-----------------------------------------------
LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.numeric_std.all;
USE work.types.all;
-----------------------------------------------

ENTITY angular_16_16_mapping IS
	PORT (
		input : IN ref_bus (0 to 146);
		block_size_control : IN std_logic_vector (3 downto 0);
		control : in std_logic_vector (1 downto 0);
		iteration_control: IN std_logic_vector (3 downto 0);
		output: OUT mapping_16_16
	);
END angular_16_16_mapping;

ARCHITECTURE comportamental OF angular_16_16_mapping IS

BEGIN
	process (input)
	begin
		if control = "000" then 
case iteration_control is
when "0000" =>
output(0, 0) <= input(0);
output(0, 1) <= input(1);
output(0, 2) <= input(2);
output(0, 3) <= input(3);
output(0, 4) <= input(4);
output(0, 5) <= input(5);
output(0, 6) <= input(6);
output(0, 7) <= input(7);
output(0, 8) <= input(8);
output(0, 9) <= input(9);
output(0, 10) <= input(10);
output(0, 11) <= input(11);
output(0, 12) <= input(12);
output(0, 13) <= input(13);
output(0, 14) <= input(14);
output(0, 15) <= input(15);
output(0, 16) <= input(1);
output(0, 17) <= input(2);
output(0, 18) <= input(3);
output(0, 19) <= input(4);
output(0, 20) <= input(5);
output(0, 21) <= input(6);
output(0, 22) <= input(7);
output(0, 23) <= input(8);
output(0, 24) <= input(9);
output(0, 25) <= input(10);
output(0, 26) <= input(11);
output(0, 27) <= input(12);
output(0, 28) <= input(13);
output(0, 29) <= input(14);
output(0, 30) <= input(15);
output(0, 31) <= input(16);
output(0, 32) <= input(2);
output(0, 33) <= input(3);
output(0, 34) <= input(4);
output(0, 35) <= input(5);
output(0, 36) <= input(6);
output(0, 37) <= input(7);
output(0, 38) <= input(8);
output(0, 39) <= input(9);
output(0, 40) <= input(10);
output(0, 41) <= input(11);
output(0, 42) <= input(12);
output(0, 43) <= input(13);
output(0, 44) <= input(14);
output(0, 45) <= input(15);
output(0, 46) <= input(16);
output(0, 47) <= input(17);
output(0, 48) <= input(3);
output(0, 49) <= input(4);
output(0, 50) <= input(5);
output(0, 51) <= input(6);
output(0, 52) <= input(7);
output(0, 53) <= input(8);
output(0, 54) <= input(9);
output(0, 55) <= input(10);
output(0, 56) <= input(11);
output(0, 57) <= input(12);
output(0, 58) <= input(13);
output(0, 59) <= input(14);
output(0, 60) <= input(15);
output(0, 61) <= input(16);
output(0, 62) <= input(17);
output(0, 63) <= input(18);
output(0, 64) <= input(4);
output(0, 65) <= input(5);
output(0, 66) <= input(6);
output(0, 67) <= input(7);
output(0, 68) <= input(8);
output(0, 69) <= input(9);
output(0, 70) <= input(10);
output(0, 71) <= input(11);
output(0, 72) <= input(12);
output(0, 73) <= input(13);
output(0, 74) <= input(14);
output(0, 75) <= input(15);
output(0, 76) <= input(16);
output(0, 77) <= input(17);
output(0, 78) <= input(18);
output(0, 79) <= input(19);
output(0, 80) <= input(5);
output(0, 81) <= input(6);
output(0, 82) <= input(7);
output(0, 83) <= input(8);
output(0, 84) <= input(9);
output(0, 85) <= input(10);
output(0, 86) <= input(11);
output(0, 87) <= input(12);
output(0, 88) <= input(13);
output(0, 89) <= input(14);
output(0, 90) <= input(15);
output(0, 91) <= input(16);
output(0, 92) <= input(17);
output(0, 93) <= input(18);
output(0, 94) <= input(19);
output(0, 95) <= input(20);
output(0, 96) <= input(6);
output(0, 97) <= input(7);
output(0, 98) <= input(8);
output(0, 99) <= input(9);
output(0, 100) <= input(10);
output(0, 101) <= input(11);
output(0, 102) <= input(12);
output(0, 103) <= input(13);
output(0, 104) <= input(14);
output(0, 105) <= input(15);
output(0, 106) <= input(16);
output(0, 107) <= input(17);
output(0, 108) <= input(18);
output(0, 109) <= input(19);
output(0, 110) <= input(20);
output(0, 111) <= input(21);
output(0, 112) <= input(7);
output(0, 113) <= input(8);
output(0, 114) <= input(9);
output(0, 115) <= input(10);
output(0, 116) <= input(11);
output(0, 117) <= input(12);
output(0, 118) <= input(13);
output(0, 119) <= input(14);
output(0, 120) <= input(15);
output(0, 121) <= input(16);
output(0, 122) <= input(17);
output(0, 123) <= input(18);
output(0, 124) <= input(19);
output(0, 125) <= input(20);
output(0, 126) <= input(21);
output(0, 127) <= input(22);
output(0, 128) <= input(8);
output(0, 129) <= input(9);
output(0, 130) <= input(10);
output(0, 131) <= input(11);
output(0, 132) <= input(12);
output(0, 133) <= input(13);
output(0, 134) <= input(14);
output(0, 135) <= input(15);
output(0, 136) <= input(16);
output(0, 137) <= input(17);
output(0, 138) <= input(18);
output(0, 139) <= input(19);
output(0, 140) <= input(20);
output(0, 141) <= input(21);
output(0, 142) <= input(22);
output(0, 143) <= input(23);
output(0, 144) <= input(9);
output(0, 145) <= input(10);
output(0, 146) <= input(11);
output(0, 147) <= input(12);
output(0, 148) <= input(13);
output(0, 149) <= input(14);
output(0, 150) <= input(15);
output(0, 151) <= input(16);
output(0, 152) <= input(17);
output(0, 153) <= input(18);
output(0, 154) <= input(19);
output(0, 155) <= input(20);
output(0, 156) <= input(21);
output(0, 157) <= input(22);
output(0, 158) <= input(23);
output(0, 159) <= input(24);
output(0, 160) <= input(10);
output(0, 161) <= input(11);
output(0, 162) <= input(12);
output(0, 163) <= input(13);
output(0, 164) <= input(14);
output(0, 165) <= input(15);
output(0, 166) <= input(16);
output(0, 167) <= input(17);
output(0, 168) <= input(18);
output(0, 169) <= input(19);
output(0, 170) <= input(20);
output(0, 171) <= input(21);
output(0, 172) <= input(22);
output(0, 173) <= input(23);
output(0, 174) <= input(24);
output(0, 175) <= input(25);
output(0, 176) <= input(11);
output(0, 177) <= input(12);
output(0, 178) <= input(13);
output(0, 179) <= input(14);
output(0, 180) <= input(15);
output(0, 181) <= input(16);
output(0, 182) <= input(17);
output(0, 183) <= input(18);
output(0, 184) <= input(19);
output(0, 185) <= input(20);
output(0, 186) <= input(21);
output(0, 187) <= input(22);
output(0, 188) <= input(23);
output(0, 189) <= input(24);
output(0, 190) <= input(25);
output(0, 191) <= input(26);
output(0, 192) <= input(12);
output(0, 193) <= input(13);
output(0, 194) <= input(14);
output(0, 195) <= input(15);
output(0, 196) <= input(16);
output(0, 197) <= input(17);
output(0, 198) <= input(18);
output(0, 199) <= input(19);
output(0, 200) <= input(20);
output(0, 201) <= input(21);
output(0, 202) <= input(22);
output(0, 203) <= input(23);
output(0, 204) <= input(24);
output(0, 205) <= input(25);
output(0, 206) <= input(26);
output(0, 207) <= input(27);
output(0, 208) <= input(13);
output(0, 209) <= input(14);
output(0, 210) <= input(15);
output(0, 211) <= input(16);
output(0, 212) <= input(17);
output(0, 213) <= input(18);
output(0, 214) <= input(19);
output(0, 215) <= input(20);
output(0, 216) <= input(21);
output(0, 217) <= input(22);
output(0, 218) <= input(23);
output(0, 219) <= input(24);
output(0, 220) <= input(25);
output(0, 221) <= input(26);
output(0, 222) <= input(27);
output(0, 223) <= input(28);
output(0, 224) <= input(14);
output(0, 225) <= input(15);
output(0, 226) <= input(16);
output(0, 227) <= input(17);
output(0, 228) <= input(18);
output(0, 229) <= input(19);
output(0, 230) <= input(20);
output(0, 231) <= input(21);
output(0, 232) <= input(22);
output(0, 233) <= input(23);
output(0, 234) <= input(24);
output(0, 235) <= input(25);
output(0, 236) <= input(26);
output(0, 237) <= input(27);
output(0, 238) <= input(28);
output(0, 239) <= input(29);
output(0, 240) <= input(15);
output(0, 241) <= input(16);
output(0, 242) <= input(17);
output(0, 243) <= input(18);
output(0, 244) <= input(19);
output(0, 245) <= input(20);
output(0, 246) <= input(21);
output(0, 247) <= input(22);
output(0, 248) <= input(23);
output(0, 249) <= input(24);
output(0, 250) <= input(25);
output(0, 251) <= input(26);
output(0, 252) <= input(27);
output(0, 253) <= input(28);
output(0, 254) <= input(29);
output(0, 255) <= input(30);
output(1, 0) <= input(31);
output(1, 1) <= input(32);
output(1, 2) <= input(33);
output(1, 3) <= input(34);
output(1, 4) <= input(35);
output(1, 5) <= input(36);
output(1, 6) <= input(37);
output(1, 7) <= input(38);
output(1, 8) <= input(39);
output(1, 9) <= input(40);
output(1, 10) <= input(41);
output(1, 11) <= input(42);
output(1, 12) <= input(43);
output(1, 13) <= input(44);
output(1, 14) <= input(45);
output(1, 15) <= input(46);
output(1, 16) <= input(32);
output(1, 17) <= input(33);
output(1, 18) <= input(34);
output(1, 19) <= input(35);
output(1, 20) <= input(36);
output(1, 21) <= input(37);
output(1, 22) <= input(38);
output(1, 23) <= input(39);
output(1, 24) <= input(40);
output(1, 25) <= input(41);
output(1, 26) <= input(42);
output(1, 27) <= input(43);
output(1, 28) <= input(44);
output(1, 29) <= input(45);
output(1, 30) <= input(46);
output(1, 31) <= input(47);
output(1, 32) <= input(33);
output(1, 33) <= input(34);
output(1, 34) <= input(35);
output(1, 35) <= input(36);
output(1, 36) <= input(37);
output(1, 37) <= input(38);
output(1, 38) <= input(39);
output(1, 39) <= input(40);
output(1, 40) <= input(41);
output(1, 41) <= input(42);
output(1, 42) <= input(43);
output(1, 43) <= input(44);
output(1, 44) <= input(45);
output(1, 45) <= input(46);
output(1, 46) <= input(47);
output(1, 47) <= input(48);
output(1, 48) <= input(34);
output(1, 49) <= input(35);
output(1, 50) <= input(36);
output(1, 51) <= input(37);
output(1, 52) <= input(38);
output(1, 53) <= input(39);
output(1, 54) <= input(40);
output(1, 55) <= input(41);
output(1, 56) <= input(42);
output(1, 57) <= input(43);
output(1, 58) <= input(44);
output(1, 59) <= input(45);
output(1, 60) <= input(46);
output(1, 61) <= input(47);
output(1, 62) <= input(48);
output(1, 63) <= input(49);
output(1, 64) <= input(35);
output(1, 65) <= input(36);
output(1, 66) <= input(37);
output(1, 67) <= input(38);
output(1, 68) <= input(39);
output(1, 69) <= input(40);
output(1, 70) <= input(41);
output(1, 71) <= input(42);
output(1, 72) <= input(43);
output(1, 73) <= input(44);
output(1, 74) <= input(45);
output(1, 75) <= input(46);
output(1, 76) <= input(47);
output(1, 77) <= input(48);
output(1, 78) <= input(49);
output(1, 79) <= input(50);
output(1, 80) <= input(4);
output(1, 81) <= input(5);
output(1, 82) <= input(6);
output(1, 83) <= input(7);
output(1, 84) <= input(8);
output(1, 85) <= input(9);
output(1, 86) <= input(10);
output(1, 87) <= input(11);
output(1, 88) <= input(12);
output(1, 89) <= input(13);
output(1, 90) <= input(14);
output(1, 91) <= input(15);
output(1, 92) <= input(16);
output(1, 93) <= input(17);
output(1, 94) <= input(18);
output(1, 95) <= input(19);
output(1, 96) <= input(5);
output(1, 97) <= input(6);
output(1, 98) <= input(7);
output(1, 99) <= input(8);
output(1, 100) <= input(9);
output(1, 101) <= input(10);
output(1, 102) <= input(11);
output(1, 103) <= input(12);
output(1, 104) <= input(13);
output(1, 105) <= input(14);
output(1, 106) <= input(15);
output(1, 107) <= input(16);
output(1, 108) <= input(17);
output(1, 109) <= input(18);
output(1, 110) <= input(19);
output(1, 111) <= input(20);
output(1, 112) <= input(6);
output(1, 113) <= input(7);
output(1, 114) <= input(8);
output(1, 115) <= input(9);
output(1, 116) <= input(10);
output(1, 117) <= input(11);
output(1, 118) <= input(12);
output(1, 119) <= input(13);
output(1, 120) <= input(14);
output(1, 121) <= input(15);
output(1, 122) <= input(16);
output(1, 123) <= input(17);
output(1, 124) <= input(18);
output(1, 125) <= input(19);
output(1, 126) <= input(20);
output(1, 127) <= input(21);
output(1, 128) <= input(7);
output(1, 129) <= input(8);
output(1, 130) <= input(9);
output(1, 131) <= input(10);
output(1, 132) <= input(11);
output(1, 133) <= input(12);
output(1, 134) <= input(13);
output(1, 135) <= input(14);
output(1, 136) <= input(15);
output(1, 137) <= input(16);
output(1, 138) <= input(17);
output(1, 139) <= input(18);
output(1, 140) <= input(19);
output(1, 141) <= input(20);
output(1, 142) <= input(21);
output(1, 143) <= input(22);
output(1, 144) <= input(8);
output(1, 145) <= input(9);
output(1, 146) <= input(10);
output(1, 147) <= input(11);
output(1, 148) <= input(12);
output(1, 149) <= input(13);
output(1, 150) <= input(14);
output(1, 151) <= input(15);
output(1, 152) <= input(16);
output(1, 153) <= input(17);
output(1, 154) <= input(18);
output(1, 155) <= input(19);
output(1, 156) <= input(20);
output(1, 157) <= input(21);
output(1, 158) <= input(22);
output(1, 159) <= input(23);
output(1, 160) <= input(40);
output(1, 161) <= input(41);
output(1, 162) <= input(42);
output(1, 163) <= input(43);
output(1, 164) <= input(44);
output(1, 165) <= input(45);
output(1, 166) <= input(46);
output(1, 167) <= input(47);
output(1, 168) <= input(48);
output(1, 169) <= input(49);
output(1, 170) <= input(50);
output(1, 171) <= input(51);
output(1, 172) <= input(52);
output(1, 173) <= input(53);
output(1, 174) <= input(54);
output(1, 175) <= input(55);
output(1, 176) <= input(41);
output(1, 177) <= input(42);
output(1, 178) <= input(43);
output(1, 179) <= input(44);
output(1, 180) <= input(45);
output(1, 181) <= input(46);
output(1, 182) <= input(47);
output(1, 183) <= input(48);
output(1, 184) <= input(49);
output(1, 185) <= input(50);
output(1, 186) <= input(51);
output(1, 187) <= input(52);
output(1, 188) <= input(53);
output(1, 189) <= input(54);
output(1, 190) <= input(55);
output(1, 191) <= input(56);
output(1, 192) <= input(42);
output(1, 193) <= input(43);
output(1, 194) <= input(44);
output(1, 195) <= input(45);
output(1, 196) <= input(46);
output(1, 197) <= input(47);
output(1, 198) <= input(48);
output(1, 199) <= input(49);
output(1, 200) <= input(50);
output(1, 201) <= input(51);
output(1, 202) <= input(52);
output(1, 203) <= input(53);
output(1, 204) <= input(54);
output(1, 205) <= input(55);
output(1, 206) <= input(56);
output(1, 207) <= input(57);
output(1, 208) <= input(43);
output(1, 209) <= input(44);
output(1, 210) <= input(45);
output(1, 211) <= input(46);
output(1, 212) <= input(47);
output(1, 213) <= input(48);
output(1, 214) <= input(49);
output(1, 215) <= input(50);
output(1, 216) <= input(51);
output(1, 217) <= input(52);
output(1, 218) <= input(53);
output(1, 219) <= input(54);
output(1, 220) <= input(55);
output(1, 221) <= input(56);
output(1, 222) <= input(57);
output(1, 223) <= input(58);
output(1, 224) <= input(44);
output(1, 225) <= input(45);
output(1, 226) <= input(46);
output(1, 227) <= input(47);
output(1, 228) <= input(48);
output(1, 229) <= input(49);
output(1, 230) <= input(50);
output(1, 231) <= input(51);
output(1, 232) <= input(52);
output(1, 233) <= input(53);
output(1, 234) <= input(54);
output(1, 235) <= input(55);
output(1, 236) <= input(56);
output(1, 237) <= input(57);
output(1, 238) <= input(58);
output(1, 239) <= input(59);
output(1, 240) <= input(45);
output(1, 241) <= input(46);
output(1, 242) <= input(47);
output(1, 243) <= input(48);
output(1, 244) <= input(49);
output(1, 245) <= input(50);
output(1, 246) <= input(51);
output(1, 247) <= input(52);
output(1, 248) <= input(53);
output(1, 249) <= input(54);
output(1, 250) <= input(55);
output(1, 251) <= input(56);
output(1, 252) <= input(57);
output(1, 253) <= input(58);
output(1, 254) <= input(59);
output(1, 255) <= input(60);
output(2, 0) <= input(31);
output(2, 1) <= input(32);
output(2, 2) <= input(33);
output(2, 3) <= input(34);
output(2, 4) <= input(35);
output(2, 5) <= input(36);
output(2, 6) <= input(37);
output(2, 7) <= input(38);
output(2, 8) <= input(39);
output(2, 9) <= input(40);
output(2, 10) <= input(41);
output(2, 11) <= input(42);
output(2, 12) <= input(43);
output(2, 13) <= input(44);
output(2, 14) <= input(45);
output(2, 15) <= input(46);
output(2, 16) <= input(32);
output(2, 17) <= input(33);
output(2, 18) <= input(34);
output(2, 19) <= input(35);
output(2, 20) <= input(36);
output(2, 21) <= input(37);
output(2, 22) <= input(38);
output(2, 23) <= input(39);
output(2, 24) <= input(40);
output(2, 25) <= input(41);
output(2, 26) <= input(42);
output(2, 27) <= input(43);
output(2, 28) <= input(44);
output(2, 29) <= input(45);
output(2, 30) <= input(46);
output(2, 31) <= input(47);
output(2, 32) <= input(1);
output(2, 33) <= input(2);
output(2, 34) <= input(3);
output(2, 35) <= input(4);
output(2, 36) <= input(5);
output(2, 37) <= input(6);
output(2, 38) <= input(7);
output(2, 39) <= input(8);
output(2, 40) <= input(9);
output(2, 41) <= input(10);
output(2, 42) <= input(11);
output(2, 43) <= input(12);
output(2, 44) <= input(13);
output(2, 45) <= input(14);
output(2, 46) <= input(15);
output(2, 47) <= input(16);
output(2, 48) <= input(2);
output(2, 49) <= input(3);
output(2, 50) <= input(4);
output(2, 51) <= input(5);
output(2, 52) <= input(6);
output(2, 53) <= input(7);
output(2, 54) <= input(8);
output(2, 55) <= input(9);
output(2, 56) <= input(10);
output(2, 57) <= input(11);
output(2, 58) <= input(12);
output(2, 59) <= input(13);
output(2, 60) <= input(14);
output(2, 61) <= input(15);
output(2, 62) <= input(16);
output(2, 63) <= input(17);
output(2, 64) <= input(3);
output(2, 65) <= input(4);
output(2, 66) <= input(5);
output(2, 67) <= input(6);
output(2, 68) <= input(7);
output(2, 69) <= input(8);
output(2, 70) <= input(9);
output(2, 71) <= input(10);
output(2, 72) <= input(11);
output(2, 73) <= input(12);
output(2, 74) <= input(13);
output(2, 75) <= input(14);
output(2, 76) <= input(15);
output(2, 77) <= input(16);
output(2, 78) <= input(17);
output(2, 79) <= input(18);
output(2, 80) <= input(35);
output(2, 81) <= input(36);
output(2, 82) <= input(37);
output(2, 83) <= input(38);
output(2, 84) <= input(39);
output(2, 85) <= input(40);
output(2, 86) <= input(41);
output(2, 87) <= input(42);
output(2, 88) <= input(43);
output(2, 89) <= input(44);
output(2, 90) <= input(45);
output(2, 91) <= input(46);
output(2, 92) <= input(47);
output(2, 93) <= input(48);
output(2, 94) <= input(49);
output(2, 95) <= input(50);
output(2, 96) <= input(36);
output(2, 97) <= input(37);
output(2, 98) <= input(38);
output(2, 99) <= input(39);
output(2, 100) <= input(40);
output(2, 101) <= input(41);
output(2, 102) <= input(42);
output(2, 103) <= input(43);
output(2, 104) <= input(44);
output(2, 105) <= input(45);
output(2, 106) <= input(46);
output(2, 107) <= input(47);
output(2, 108) <= input(48);
output(2, 109) <= input(49);
output(2, 110) <= input(50);
output(2, 111) <= input(51);
output(2, 112) <= input(37);
output(2, 113) <= input(38);
output(2, 114) <= input(39);
output(2, 115) <= input(40);
output(2, 116) <= input(41);
output(2, 117) <= input(42);
output(2, 118) <= input(43);
output(2, 119) <= input(44);
output(2, 120) <= input(45);
output(2, 121) <= input(46);
output(2, 122) <= input(47);
output(2, 123) <= input(48);
output(2, 124) <= input(49);
output(2, 125) <= input(50);
output(2, 126) <= input(51);
output(2, 127) <= input(52);
output(2, 128) <= input(6);
output(2, 129) <= input(7);
output(2, 130) <= input(8);
output(2, 131) <= input(9);
output(2, 132) <= input(10);
output(2, 133) <= input(11);
output(2, 134) <= input(12);
output(2, 135) <= input(13);
output(2, 136) <= input(14);
output(2, 137) <= input(15);
output(2, 138) <= input(16);
output(2, 139) <= input(17);
output(2, 140) <= input(18);
output(2, 141) <= input(19);
output(2, 142) <= input(20);
output(2, 143) <= input(21);
output(2, 144) <= input(7);
output(2, 145) <= input(8);
output(2, 146) <= input(9);
output(2, 147) <= input(10);
output(2, 148) <= input(11);
output(2, 149) <= input(12);
output(2, 150) <= input(13);
output(2, 151) <= input(14);
output(2, 152) <= input(15);
output(2, 153) <= input(16);
output(2, 154) <= input(17);
output(2, 155) <= input(18);
output(2, 156) <= input(19);
output(2, 157) <= input(20);
output(2, 158) <= input(21);
output(2, 159) <= input(22);
output(2, 160) <= input(39);
output(2, 161) <= input(40);
output(2, 162) <= input(41);
output(2, 163) <= input(42);
output(2, 164) <= input(43);
output(2, 165) <= input(44);
output(2, 166) <= input(45);
output(2, 167) <= input(46);
output(2, 168) <= input(47);
output(2, 169) <= input(48);
output(2, 170) <= input(49);
output(2, 171) <= input(50);
output(2, 172) <= input(51);
output(2, 173) <= input(52);
output(2, 174) <= input(53);
output(2, 175) <= input(54);
output(2, 176) <= input(40);
output(2, 177) <= input(41);
output(2, 178) <= input(42);
output(2, 179) <= input(43);
output(2, 180) <= input(44);
output(2, 181) <= input(45);
output(2, 182) <= input(46);
output(2, 183) <= input(47);
output(2, 184) <= input(48);
output(2, 185) <= input(49);
output(2, 186) <= input(50);
output(2, 187) <= input(51);
output(2, 188) <= input(52);
output(2, 189) <= input(53);
output(2, 190) <= input(54);
output(2, 191) <= input(55);
output(2, 192) <= input(41);
output(2, 193) <= input(42);
output(2, 194) <= input(43);
output(2, 195) <= input(44);
output(2, 196) <= input(45);
output(2, 197) <= input(46);
output(2, 198) <= input(47);
output(2, 199) <= input(48);
output(2, 200) <= input(49);
output(2, 201) <= input(50);
output(2, 202) <= input(51);
output(2, 203) <= input(52);
output(2, 204) <= input(53);
output(2, 205) <= input(54);
output(2, 206) <= input(55);
output(2, 207) <= input(56);
output(2, 208) <= input(10);
output(2, 209) <= input(11);
output(2, 210) <= input(12);
output(2, 211) <= input(13);
output(2, 212) <= input(14);
output(2, 213) <= input(15);
output(2, 214) <= input(16);
output(2, 215) <= input(17);
output(2, 216) <= input(18);
output(2, 217) <= input(19);
output(2, 218) <= input(20);
output(2, 219) <= input(21);
output(2, 220) <= input(22);
output(2, 221) <= input(23);
output(2, 222) <= input(24);
output(2, 223) <= input(25);
output(2, 224) <= input(11);
output(2, 225) <= input(12);
output(2, 226) <= input(13);
output(2, 227) <= input(14);
output(2, 228) <= input(15);
output(2, 229) <= input(16);
output(2, 230) <= input(17);
output(2, 231) <= input(18);
output(2, 232) <= input(19);
output(2, 233) <= input(20);
output(2, 234) <= input(21);
output(2, 235) <= input(22);
output(2, 236) <= input(23);
output(2, 237) <= input(24);
output(2, 238) <= input(25);
output(2, 239) <= input(26);
output(2, 240) <= input(12);
output(2, 241) <= input(13);
output(2, 242) <= input(14);
output(2, 243) <= input(15);
output(2, 244) <= input(16);
output(2, 245) <= input(17);
output(2, 246) <= input(18);
output(2, 247) <= input(19);
output(2, 248) <= input(20);
output(2, 249) <= input(21);
output(2, 250) <= input(22);
output(2, 251) <= input(23);
output(2, 252) <= input(24);
output(2, 253) <= input(25);
output(2, 254) <= input(26);
output(2, 255) <= input(27);
output(3, 0) <= input(31);
output(3, 1) <= input(32);
output(3, 2) <= input(33);
output(3, 3) <= input(34);
output(3, 4) <= input(35);
output(3, 5) <= input(36);
output(3, 6) <= input(37);
output(3, 7) <= input(38);
output(3, 8) <= input(39);
output(3, 9) <= input(40);
output(3, 10) <= input(41);
output(3, 11) <= input(42);
output(3, 12) <= input(43);
output(3, 13) <= input(44);
output(3, 14) <= input(45);
output(3, 15) <= input(46);
output(3, 16) <= input(0);
output(3, 17) <= input(1);
output(3, 18) <= input(2);
output(3, 19) <= input(3);
output(3, 20) <= input(4);
output(3, 21) <= input(5);
output(3, 22) <= input(6);
output(3, 23) <= input(7);
output(3, 24) <= input(8);
output(3, 25) <= input(9);
output(3, 26) <= input(10);
output(3, 27) <= input(11);
output(3, 28) <= input(12);
output(3, 29) <= input(13);
output(3, 30) <= input(14);
output(3, 31) <= input(15);
output(3, 32) <= input(1);
output(3, 33) <= input(2);
output(3, 34) <= input(3);
output(3, 35) <= input(4);
output(3, 36) <= input(5);
output(3, 37) <= input(6);
output(3, 38) <= input(7);
output(3, 39) <= input(8);
output(3, 40) <= input(9);
output(3, 41) <= input(10);
output(3, 42) <= input(11);
output(3, 43) <= input(12);
output(3, 44) <= input(13);
output(3, 45) <= input(14);
output(3, 46) <= input(15);
output(3, 47) <= input(16);
output(3, 48) <= input(33);
output(3, 49) <= input(34);
output(3, 50) <= input(35);
output(3, 51) <= input(36);
output(3, 52) <= input(37);
output(3, 53) <= input(38);
output(3, 54) <= input(39);
output(3, 55) <= input(40);
output(3, 56) <= input(41);
output(3, 57) <= input(42);
output(3, 58) <= input(43);
output(3, 59) <= input(44);
output(3, 60) <= input(45);
output(3, 61) <= input(46);
output(3, 62) <= input(47);
output(3, 63) <= input(48);
output(3, 64) <= input(34);
output(3, 65) <= input(35);
output(3, 66) <= input(36);
output(3, 67) <= input(37);
output(3, 68) <= input(38);
output(3, 69) <= input(39);
output(3, 70) <= input(40);
output(3, 71) <= input(41);
output(3, 72) <= input(42);
output(3, 73) <= input(43);
output(3, 74) <= input(44);
output(3, 75) <= input(45);
output(3, 76) <= input(46);
output(3, 77) <= input(47);
output(3, 78) <= input(48);
output(3, 79) <= input(49);
output(3, 80) <= input(3);
output(3, 81) <= input(4);
output(3, 82) <= input(5);
output(3, 83) <= input(6);
output(3, 84) <= input(7);
output(3, 85) <= input(8);
output(3, 86) <= input(9);
output(3, 87) <= input(10);
output(3, 88) <= input(11);
output(3, 89) <= input(12);
output(3, 90) <= input(13);
output(3, 91) <= input(14);
output(3, 92) <= input(15);
output(3, 93) <= input(16);
output(3, 94) <= input(17);
output(3, 95) <= input(18);
output(3, 96) <= input(4);
output(3, 97) <= input(5);
output(3, 98) <= input(6);
output(3, 99) <= input(7);
output(3, 100) <= input(8);
output(3, 101) <= input(9);
output(3, 102) <= input(10);
output(3, 103) <= input(11);
output(3, 104) <= input(12);
output(3, 105) <= input(13);
output(3, 106) <= input(14);
output(3, 107) <= input(15);
output(3, 108) <= input(16);
output(3, 109) <= input(17);
output(3, 110) <= input(18);
output(3, 111) <= input(19);
output(3, 112) <= input(36);
output(3, 113) <= input(37);
output(3, 114) <= input(38);
output(3, 115) <= input(39);
output(3, 116) <= input(40);
output(3, 117) <= input(41);
output(3, 118) <= input(42);
output(3, 119) <= input(43);
output(3, 120) <= input(44);
output(3, 121) <= input(45);
output(3, 122) <= input(46);
output(3, 123) <= input(47);
output(3, 124) <= input(48);
output(3, 125) <= input(49);
output(3, 126) <= input(50);
output(3, 127) <= input(51);
output(3, 128) <= input(5);
output(3, 129) <= input(6);
output(3, 130) <= input(7);
output(3, 131) <= input(8);
output(3, 132) <= input(9);
output(3, 133) <= input(10);
output(3, 134) <= input(11);
output(3, 135) <= input(12);
output(3, 136) <= input(13);
output(3, 137) <= input(14);
output(3, 138) <= input(15);
output(3, 139) <= input(16);
output(3, 140) <= input(17);
output(3, 141) <= input(18);
output(3, 142) <= input(19);
output(3, 143) <= input(20);
output(3, 144) <= input(6);
output(3, 145) <= input(7);
output(3, 146) <= input(8);
output(3, 147) <= input(9);
output(3, 148) <= input(10);
output(3, 149) <= input(11);
output(3, 150) <= input(12);
output(3, 151) <= input(13);
output(3, 152) <= input(14);
output(3, 153) <= input(15);
output(3, 154) <= input(16);
output(3, 155) <= input(17);
output(3, 156) <= input(18);
output(3, 157) <= input(19);
output(3, 158) <= input(20);
output(3, 159) <= input(21);
output(3, 160) <= input(38);
output(3, 161) <= input(39);
output(3, 162) <= input(40);
output(3, 163) <= input(41);
output(3, 164) <= input(42);
output(3, 165) <= input(43);
output(3, 166) <= input(44);
output(3, 167) <= input(45);
output(3, 168) <= input(46);
output(3, 169) <= input(47);
output(3, 170) <= input(48);
output(3, 171) <= input(49);
output(3, 172) <= input(50);
output(3, 173) <= input(51);
output(3, 174) <= input(52);
output(3, 175) <= input(53);
output(3, 176) <= input(39);
output(3, 177) <= input(40);
output(3, 178) <= input(41);
output(3, 179) <= input(42);
output(3, 180) <= input(43);
output(3, 181) <= input(44);
output(3, 182) <= input(45);
output(3, 183) <= input(46);
output(3, 184) <= input(47);
output(3, 185) <= input(48);
output(3, 186) <= input(49);
output(3, 187) <= input(50);
output(3, 188) <= input(51);
output(3, 189) <= input(52);
output(3, 190) <= input(53);
output(3, 191) <= input(54);
output(3, 192) <= input(8);
output(3, 193) <= input(9);
output(3, 194) <= input(10);
output(3, 195) <= input(11);
output(3, 196) <= input(12);
output(3, 197) <= input(13);
output(3, 198) <= input(14);
output(3, 199) <= input(15);
output(3, 200) <= input(16);
output(3, 201) <= input(17);
output(3, 202) <= input(18);
output(3, 203) <= input(19);
output(3, 204) <= input(20);
output(3, 205) <= input(21);
output(3, 206) <= input(22);
output(3, 207) <= input(23);
output(3, 208) <= input(9);
output(3, 209) <= input(10);
output(3, 210) <= input(11);
output(3, 211) <= input(12);
output(3, 212) <= input(13);
output(3, 213) <= input(14);
output(3, 214) <= input(15);
output(3, 215) <= input(16);
output(3, 216) <= input(17);
output(3, 217) <= input(18);
output(3, 218) <= input(19);
output(3, 219) <= input(20);
output(3, 220) <= input(21);
output(3, 221) <= input(22);
output(3, 222) <= input(23);
output(3, 223) <= input(24);
output(3, 224) <= input(41);
output(3, 225) <= input(42);
output(3, 226) <= input(43);
output(3, 227) <= input(44);
output(3, 228) <= input(45);
output(3, 229) <= input(46);
output(3, 230) <= input(47);
output(3, 231) <= input(48);
output(3, 232) <= input(49);
output(3, 233) <= input(50);
output(3, 234) <= input(51);
output(3, 235) <= input(52);
output(3, 236) <= input(53);
output(3, 237) <= input(54);
output(3, 238) <= input(55);
output(3, 239) <= input(56);
output(3, 240) <= input(42);
output(3, 241) <= input(43);
output(3, 242) <= input(44);
output(3, 243) <= input(45);
output(3, 244) <= input(46);
output(3, 245) <= input(47);
output(3, 246) <= input(48);
output(3, 247) <= input(49);
output(3, 248) <= input(50);
output(3, 249) <= input(51);
output(3, 250) <= input(52);
output(3, 251) <= input(53);
output(3, 252) <= input(54);
output(3, 253) <= input(55);
output(3, 254) <= input(56);
output(3, 255) <= input(57);
output(4, 0) <= input(31);
output(4, 1) <= input(32);
output(4, 2) <= input(33);
output(4, 3) <= input(34);
output(4, 4) <= input(35);
output(4, 5) <= input(36);
output(4, 6) <= input(37);
output(4, 7) <= input(38);
output(4, 8) <= input(39);
output(4, 9) <= input(40);
output(4, 10) <= input(41);
output(4, 11) <= input(42);
output(4, 12) <= input(43);
output(4, 13) <= input(44);
output(4, 14) <= input(45);
output(4, 15) <= input(46);
output(4, 16) <= input(0);
output(4, 17) <= input(1);
output(4, 18) <= input(2);
output(4, 19) <= input(3);
output(4, 20) <= input(4);
output(4, 21) <= input(5);
output(4, 22) <= input(6);
output(4, 23) <= input(7);
output(4, 24) <= input(8);
output(4, 25) <= input(9);
output(4, 26) <= input(10);
output(4, 27) <= input(11);
output(4, 28) <= input(12);
output(4, 29) <= input(13);
output(4, 30) <= input(14);
output(4, 31) <= input(15);
output(4, 32) <= input(32);
output(4, 33) <= input(33);
output(4, 34) <= input(34);
output(4, 35) <= input(35);
output(4, 36) <= input(36);
output(4, 37) <= input(37);
output(4, 38) <= input(38);
output(4, 39) <= input(39);
output(4, 40) <= input(40);
output(4, 41) <= input(41);
output(4, 42) <= input(42);
output(4, 43) <= input(43);
output(4, 44) <= input(44);
output(4, 45) <= input(45);
output(4, 46) <= input(46);
output(4, 47) <= input(47);
output(4, 48) <= input(33);
output(4, 49) <= input(34);
output(4, 50) <= input(35);
output(4, 51) <= input(36);
output(4, 52) <= input(37);
output(4, 53) <= input(38);
output(4, 54) <= input(39);
output(4, 55) <= input(40);
output(4, 56) <= input(41);
output(4, 57) <= input(42);
output(4, 58) <= input(43);
output(4, 59) <= input(44);
output(4, 60) <= input(45);
output(4, 61) <= input(46);
output(4, 62) <= input(47);
output(4, 63) <= input(48);
output(4, 64) <= input(2);
output(4, 65) <= input(3);
output(4, 66) <= input(4);
output(4, 67) <= input(5);
output(4, 68) <= input(6);
output(4, 69) <= input(7);
output(4, 70) <= input(8);
output(4, 71) <= input(9);
output(4, 72) <= input(10);
output(4, 73) <= input(11);
output(4, 74) <= input(12);
output(4, 75) <= input(13);
output(4, 76) <= input(14);
output(4, 77) <= input(15);
output(4, 78) <= input(16);
output(4, 79) <= input(17);
output(4, 80) <= input(34);
output(4, 81) <= input(35);
output(4, 82) <= input(36);
output(4, 83) <= input(37);
output(4, 84) <= input(38);
output(4, 85) <= input(39);
output(4, 86) <= input(40);
output(4, 87) <= input(41);
output(4, 88) <= input(42);
output(4, 89) <= input(43);
output(4, 90) <= input(44);
output(4, 91) <= input(45);
output(4, 92) <= input(46);
output(4, 93) <= input(47);
output(4, 94) <= input(48);
output(4, 95) <= input(49);
output(4, 96) <= input(3);
output(4, 97) <= input(4);
output(4, 98) <= input(5);
output(4, 99) <= input(6);
output(4, 100) <= input(7);
output(4, 101) <= input(8);
output(4, 102) <= input(9);
output(4, 103) <= input(10);
output(4, 104) <= input(11);
output(4, 105) <= input(12);
output(4, 106) <= input(13);
output(4, 107) <= input(14);
output(4, 108) <= input(15);
output(4, 109) <= input(16);
output(4, 110) <= input(17);
output(4, 111) <= input(18);
output(4, 112) <= input(4);
output(4, 113) <= input(5);
output(4, 114) <= input(6);
output(4, 115) <= input(7);
output(4, 116) <= input(8);
output(4, 117) <= input(9);
output(4, 118) <= input(10);
output(4, 119) <= input(11);
output(4, 120) <= input(12);
output(4, 121) <= input(13);
output(4, 122) <= input(14);
output(4, 123) <= input(15);
output(4, 124) <= input(16);
output(4, 125) <= input(17);
output(4, 126) <= input(18);
output(4, 127) <= input(19);
output(4, 128) <= input(36);
output(4, 129) <= input(37);
output(4, 130) <= input(38);
output(4, 131) <= input(39);
output(4, 132) <= input(40);
output(4, 133) <= input(41);
output(4, 134) <= input(42);
output(4, 135) <= input(43);
output(4, 136) <= input(44);
output(4, 137) <= input(45);
output(4, 138) <= input(46);
output(4, 139) <= input(47);
output(4, 140) <= input(48);
output(4, 141) <= input(49);
output(4, 142) <= input(50);
output(4, 143) <= input(51);
output(4, 144) <= input(5);
output(4, 145) <= input(6);
output(4, 146) <= input(7);
output(4, 147) <= input(8);
output(4, 148) <= input(9);
output(4, 149) <= input(10);
output(4, 150) <= input(11);
output(4, 151) <= input(12);
output(4, 152) <= input(13);
output(4, 153) <= input(14);
output(4, 154) <= input(15);
output(4, 155) <= input(16);
output(4, 156) <= input(17);
output(4, 157) <= input(18);
output(4, 158) <= input(19);
output(4, 159) <= input(20);
output(4, 160) <= input(37);
output(4, 161) <= input(38);
output(4, 162) <= input(39);
output(4, 163) <= input(40);
output(4, 164) <= input(41);
output(4, 165) <= input(42);
output(4, 166) <= input(43);
output(4, 167) <= input(44);
output(4, 168) <= input(45);
output(4, 169) <= input(46);
output(4, 170) <= input(47);
output(4, 171) <= input(48);
output(4, 172) <= input(49);
output(4, 173) <= input(50);
output(4, 174) <= input(51);
output(4, 175) <= input(52);
output(4, 176) <= input(38);
output(4, 177) <= input(39);
output(4, 178) <= input(40);
output(4, 179) <= input(41);
output(4, 180) <= input(42);
output(4, 181) <= input(43);
output(4, 182) <= input(44);
output(4, 183) <= input(45);
output(4, 184) <= input(46);
output(4, 185) <= input(47);
output(4, 186) <= input(48);
output(4, 187) <= input(49);
output(4, 188) <= input(50);
output(4, 189) <= input(51);
output(4, 190) <= input(52);
output(4, 191) <= input(53);
output(4, 192) <= input(7);
output(4, 193) <= input(8);
output(4, 194) <= input(9);
output(4, 195) <= input(10);
output(4, 196) <= input(11);
output(4, 197) <= input(12);
output(4, 198) <= input(13);
output(4, 199) <= input(14);
output(4, 200) <= input(15);
output(4, 201) <= input(16);
output(4, 202) <= input(17);
output(4, 203) <= input(18);
output(4, 204) <= input(19);
output(4, 205) <= input(20);
output(4, 206) <= input(21);
output(4, 207) <= input(22);
output(4, 208) <= input(39);
output(4, 209) <= input(40);
output(4, 210) <= input(41);
output(4, 211) <= input(42);
output(4, 212) <= input(43);
output(4, 213) <= input(44);
output(4, 214) <= input(45);
output(4, 215) <= input(46);
output(4, 216) <= input(47);
output(4, 217) <= input(48);
output(4, 218) <= input(49);
output(4, 219) <= input(50);
output(4, 220) <= input(51);
output(4, 221) <= input(52);
output(4, 222) <= input(53);
output(4, 223) <= input(54);
output(4, 224) <= input(8);
output(4, 225) <= input(9);
output(4, 226) <= input(10);
output(4, 227) <= input(11);
output(4, 228) <= input(12);
output(4, 229) <= input(13);
output(4, 230) <= input(14);
output(4, 231) <= input(15);
output(4, 232) <= input(16);
output(4, 233) <= input(17);
output(4, 234) <= input(18);
output(4, 235) <= input(19);
output(4, 236) <= input(20);
output(4, 237) <= input(21);
output(4, 238) <= input(22);
output(4, 239) <= input(23);
output(4, 240) <= input(9);
output(4, 241) <= input(10);
output(4, 242) <= input(11);
output(4, 243) <= input(12);
output(4, 244) <= input(13);
output(4, 245) <= input(14);
output(4, 246) <= input(15);
output(4, 247) <= input(16);
output(4, 248) <= input(17);
output(4, 249) <= input(18);
output(4, 250) <= input(19);
output(4, 251) <= input(20);
output(4, 252) <= input(21);
output(4, 253) <= input(22);
output(4, 254) <= input(23);
output(4, 255) <= input(24);
output(5, 0) <= input(31);
output(5, 1) <= input(32);
output(5, 2) <= input(33);
output(5, 3) <= input(34);
output(5, 4) <= input(35);
output(5, 5) <= input(36);
output(5, 6) <= input(37);
output(5, 7) <= input(38);
output(5, 8) <= input(39);
output(5, 9) <= input(40);
output(5, 10) <= input(41);
output(5, 11) <= input(42);
output(5, 12) <= input(43);
output(5, 13) <= input(44);
output(5, 14) <= input(45);
output(5, 15) <= input(46);
output(5, 16) <= input(0);
output(5, 17) <= input(1);
output(5, 18) <= input(2);
output(5, 19) <= input(3);
output(5, 20) <= input(4);
output(5, 21) <= input(5);
output(5, 22) <= input(6);
output(5, 23) <= input(7);
output(5, 24) <= input(8);
output(5, 25) <= input(9);
output(5, 26) <= input(10);
output(5, 27) <= input(11);
output(5, 28) <= input(12);
output(5, 29) <= input(13);
output(5, 30) <= input(14);
output(5, 31) <= input(15);
output(5, 32) <= input(32);
output(5, 33) <= input(33);
output(5, 34) <= input(34);
output(5, 35) <= input(35);
output(5, 36) <= input(36);
output(5, 37) <= input(37);
output(5, 38) <= input(38);
output(5, 39) <= input(39);
output(5, 40) <= input(40);
output(5, 41) <= input(41);
output(5, 42) <= input(42);
output(5, 43) <= input(43);
output(5, 44) <= input(44);
output(5, 45) <= input(45);
output(5, 46) <= input(46);
output(5, 47) <= input(47);
output(5, 48) <= input(1);
output(5, 49) <= input(2);
output(5, 50) <= input(3);
output(5, 51) <= input(4);
output(5, 52) <= input(5);
output(5, 53) <= input(6);
output(5, 54) <= input(7);
output(5, 55) <= input(8);
output(5, 56) <= input(9);
output(5, 57) <= input(10);
output(5, 58) <= input(11);
output(5, 59) <= input(12);
output(5, 60) <= input(13);
output(5, 61) <= input(14);
output(5, 62) <= input(15);
output(5, 63) <= input(16);
output(5, 64) <= input(33);
output(5, 65) <= input(34);
output(5, 66) <= input(35);
output(5, 67) <= input(36);
output(5, 68) <= input(37);
output(5, 69) <= input(38);
output(5, 70) <= input(39);
output(5, 71) <= input(40);
output(5, 72) <= input(41);
output(5, 73) <= input(42);
output(5, 74) <= input(43);
output(5, 75) <= input(44);
output(5, 76) <= input(45);
output(5, 77) <= input(46);
output(5, 78) <= input(47);
output(5, 79) <= input(48);
output(5, 80) <= input(2);
output(5, 81) <= input(3);
output(5, 82) <= input(4);
output(5, 83) <= input(5);
output(5, 84) <= input(6);
output(5, 85) <= input(7);
output(5, 86) <= input(8);
output(5, 87) <= input(9);
output(5, 88) <= input(10);
output(5, 89) <= input(11);
output(5, 90) <= input(12);
output(5, 91) <= input(13);
output(5, 92) <= input(14);
output(5, 93) <= input(15);
output(5, 94) <= input(16);
output(5, 95) <= input(17);
output(5, 96) <= input(34);
output(5, 97) <= input(35);
output(5, 98) <= input(36);
output(5, 99) <= input(37);
output(5, 100) <= input(38);
output(5, 101) <= input(39);
output(5, 102) <= input(40);
output(5, 103) <= input(41);
output(5, 104) <= input(42);
output(5, 105) <= input(43);
output(5, 106) <= input(44);
output(5, 107) <= input(45);
output(5, 108) <= input(46);
output(5, 109) <= input(47);
output(5, 110) <= input(48);
output(5, 111) <= input(49);
output(5, 112) <= input(35);
output(5, 113) <= input(36);
output(5, 114) <= input(37);
output(5, 115) <= input(38);
output(5, 116) <= input(39);
output(5, 117) <= input(40);
output(5, 118) <= input(41);
output(5, 119) <= input(42);
output(5, 120) <= input(43);
output(5, 121) <= input(44);
output(5, 122) <= input(45);
output(5, 123) <= input(46);
output(5, 124) <= input(47);
output(5, 125) <= input(48);
output(5, 126) <= input(49);
output(5, 127) <= input(50);
output(5, 128) <= input(4);
output(5, 129) <= input(5);
output(5, 130) <= input(6);
output(5, 131) <= input(7);
output(5, 132) <= input(8);
output(5, 133) <= input(9);
output(5, 134) <= input(10);
output(5, 135) <= input(11);
output(5, 136) <= input(12);
output(5, 137) <= input(13);
output(5, 138) <= input(14);
output(5, 139) <= input(15);
output(5, 140) <= input(16);
output(5, 141) <= input(17);
output(5, 142) <= input(18);
output(5, 143) <= input(19);
output(5, 144) <= input(36);
output(5, 145) <= input(37);
output(5, 146) <= input(38);
output(5, 147) <= input(39);
output(5, 148) <= input(40);
output(5, 149) <= input(41);
output(5, 150) <= input(42);
output(5, 151) <= input(43);
output(5, 152) <= input(44);
output(5, 153) <= input(45);
output(5, 154) <= input(46);
output(5, 155) <= input(47);
output(5, 156) <= input(48);
output(5, 157) <= input(49);
output(5, 158) <= input(50);
output(5, 159) <= input(51);
output(5, 160) <= input(5);
output(5, 161) <= input(6);
output(5, 162) <= input(7);
output(5, 163) <= input(8);
output(5, 164) <= input(9);
output(5, 165) <= input(10);
output(5, 166) <= input(11);
output(5, 167) <= input(12);
output(5, 168) <= input(13);
output(5, 169) <= input(14);
output(5, 170) <= input(15);
output(5, 171) <= input(16);
output(5, 172) <= input(17);
output(5, 173) <= input(18);
output(5, 174) <= input(19);
output(5, 175) <= input(20);
output(5, 176) <= input(37);
output(5, 177) <= input(38);
output(5, 178) <= input(39);
output(5, 179) <= input(40);
output(5, 180) <= input(41);
output(5, 181) <= input(42);
output(5, 182) <= input(43);
output(5, 183) <= input(44);
output(5, 184) <= input(45);
output(5, 185) <= input(46);
output(5, 186) <= input(47);
output(5, 187) <= input(48);
output(5, 188) <= input(49);
output(5, 189) <= input(50);
output(5, 190) <= input(51);
output(5, 191) <= input(52);
output(5, 192) <= input(6);
output(5, 193) <= input(7);
output(5, 194) <= input(8);
output(5, 195) <= input(9);
output(5, 196) <= input(10);
output(5, 197) <= input(11);
output(5, 198) <= input(12);
output(5, 199) <= input(13);
output(5, 200) <= input(14);
output(5, 201) <= input(15);
output(5, 202) <= input(16);
output(5, 203) <= input(17);
output(5, 204) <= input(18);
output(5, 205) <= input(19);
output(5, 206) <= input(20);
output(5, 207) <= input(21);
output(5, 208) <= input(38);
output(5, 209) <= input(39);
output(5, 210) <= input(40);
output(5, 211) <= input(41);
output(5, 212) <= input(42);
output(5, 213) <= input(43);
output(5, 214) <= input(44);
output(5, 215) <= input(45);
output(5, 216) <= input(46);
output(5, 217) <= input(47);
output(5, 218) <= input(48);
output(5, 219) <= input(49);
output(5, 220) <= input(50);
output(5, 221) <= input(51);
output(5, 222) <= input(52);
output(5, 223) <= input(53);
output(5, 224) <= input(7);
output(5, 225) <= input(8);
output(5, 226) <= input(9);
output(5, 227) <= input(10);
output(5, 228) <= input(11);
output(5, 229) <= input(12);
output(5, 230) <= input(13);
output(5, 231) <= input(14);
output(5, 232) <= input(15);
output(5, 233) <= input(16);
output(5, 234) <= input(17);
output(5, 235) <= input(18);
output(5, 236) <= input(19);
output(5, 237) <= input(20);
output(5, 238) <= input(21);
output(5, 239) <= input(22);
output(5, 240) <= input(8);
output(5, 241) <= input(9);
output(5, 242) <= input(10);
output(5, 243) <= input(11);
output(5, 244) <= input(12);
output(5, 245) <= input(13);
output(5, 246) <= input(14);
output(5, 247) <= input(15);
output(5, 248) <= input(16);
output(5, 249) <= input(17);
output(5, 250) <= input(18);
output(5, 251) <= input(19);
output(5, 252) <= input(20);
output(5, 253) <= input(21);
output(5, 254) <= input(22);
output(5, 255) <= input(23);
when "0001" =>
output(0, 0) <= input(0);
output(0, 1) <= input(1);
output(0, 2) <= input(2);
output(0, 3) <= input(3);
output(0, 4) <= input(4);
output(0, 5) <= input(5);
output(0, 6) <= input(6);
output(0, 7) <= input(7);
output(0, 8) <= input(8);
output(0, 9) <= input(9);
output(0, 10) <= input(10);
output(0, 11) <= input(11);
output(0, 12) <= input(12);
output(0, 13) <= input(13);
output(0, 14) <= input(14);
output(0, 15) <= input(15);
output(0, 16) <= input(16);
output(0, 17) <= input(17);
output(0, 18) <= input(18);
output(0, 19) <= input(19);
output(0, 20) <= input(20);
output(0, 21) <= input(21);
output(0, 22) <= input(22);
output(0, 23) <= input(23);
output(0, 24) <= input(24);
output(0, 25) <= input(25);
output(0, 26) <= input(26);
output(0, 27) <= input(27);
output(0, 28) <= input(28);
output(0, 29) <= input(29);
output(0, 30) <= input(30);
output(0, 31) <= input(31);
output(0, 32) <= input(1);
output(0, 33) <= input(2);
output(0, 34) <= input(3);
output(0, 35) <= input(4);
output(0, 36) <= input(5);
output(0, 37) <= input(6);
output(0, 38) <= input(7);
output(0, 39) <= input(8);
output(0, 40) <= input(9);
output(0, 41) <= input(10);
output(0, 42) <= input(11);
output(0, 43) <= input(12);
output(0, 44) <= input(13);
output(0, 45) <= input(14);
output(0, 46) <= input(15);
output(0, 47) <= input(32);
output(0, 48) <= input(17);
output(0, 49) <= input(18);
output(0, 50) <= input(19);
output(0, 51) <= input(20);
output(0, 52) <= input(21);
output(0, 53) <= input(22);
output(0, 54) <= input(23);
output(0, 55) <= input(24);
output(0, 56) <= input(25);
output(0, 57) <= input(26);
output(0, 58) <= input(27);
output(0, 59) <= input(28);
output(0, 60) <= input(29);
output(0, 61) <= input(30);
output(0, 62) <= input(31);
output(0, 63) <= input(33);
output(0, 64) <= input(2);
output(0, 65) <= input(3);
output(0, 66) <= input(4);
output(0, 67) <= input(5);
output(0, 68) <= input(6);
output(0, 69) <= input(7);
output(0, 70) <= input(8);
output(0, 71) <= input(9);
output(0, 72) <= input(10);
output(0, 73) <= input(11);
output(0, 74) <= input(12);
output(0, 75) <= input(13);
output(0, 76) <= input(14);
output(0, 77) <= input(15);
output(0, 78) <= input(32);
output(0, 79) <= input(34);
output(0, 80) <= input(18);
output(0, 81) <= input(19);
output(0, 82) <= input(20);
output(0, 83) <= input(21);
output(0, 84) <= input(22);
output(0, 85) <= input(23);
output(0, 86) <= input(24);
output(0, 87) <= input(25);
output(0, 88) <= input(26);
output(0, 89) <= input(27);
output(0, 90) <= input(28);
output(0, 91) <= input(29);
output(0, 92) <= input(30);
output(0, 93) <= input(31);
output(0, 94) <= input(33);
output(0, 95) <= input(35);
output(0, 96) <= input(3);
output(0, 97) <= input(4);
output(0, 98) <= input(5);
output(0, 99) <= input(6);
output(0, 100) <= input(7);
output(0, 101) <= input(8);
output(0, 102) <= input(9);
output(0, 103) <= input(10);
output(0, 104) <= input(11);
output(0, 105) <= input(12);
output(0, 106) <= input(13);
output(0, 107) <= input(14);
output(0, 108) <= input(15);
output(0, 109) <= input(32);
output(0, 110) <= input(34);
output(0, 111) <= input(36);
output(0, 112) <= input(19);
output(0, 113) <= input(20);
output(0, 114) <= input(21);
output(0, 115) <= input(22);
output(0, 116) <= input(23);
output(0, 117) <= input(24);
output(0, 118) <= input(25);
output(0, 119) <= input(26);
output(0, 120) <= input(27);
output(0, 121) <= input(28);
output(0, 122) <= input(29);
output(0, 123) <= input(30);
output(0, 124) <= input(31);
output(0, 125) <= input(33);
output(0, 126) <= input(35);
output(0, 127) <= input(37);
output(0, 128) <= input(4);
output(0, 129) <= input(5);
output(0, 130) <= input(6);
output(0, 131) <= input(7);
output(0, 132) <= input(8);
output(0, 133) <= input(9);
output(0, 134) <= input(10);
output(0, 135) <= input(11);
output(0, 136) <= input(12);
output(0, 137) <= input(13);
output(0, 138) <= input(14);
output(0, 139) <= input(15);
output(0, 140) <= input(32);
output(0, 141) <= input(34);
output(0, 142) <= input(36);
output(0, 143) <= input(38);
output(0, 144) <= input(20);
output(0, 145) <= input(21);
output(0, 146) <= input(22);
output(0, 147) <= input(23);
output(0, 148) <= input(24);
output(0, 149) <= input(25);
output(0, 150) <= input(26);
output(0, 151) <= input(27);
output(0, 152) <= input(28);
output(0, 153) <= input(29);
output(0, 154) <= input(30);
output(0, 155) <= input(31);
output(0, 156) <= input(33);
output(0, 157) <= input(35);
output(0, 158) <= input(37);
output(0, 159) <= input(39);
output(0, 160) <= input(5);
output(0, 161) <= input(6);
output(0, 162) <= input(7);
output(0, 163) <= input(8);
output(0, 164) <= input(9);
output(0, 165) <= input(10);
output(0, 166) <= input(11);
output(0, 167) <= input(12);
output(0, 168) <= input(13);
output(0, 169) <= input(14);
output(0, 170) <= input(15);
output(0, 171) <= input(32);
output(0, 172) <= input(34);
output(0, 173) <= input(36);
output(0, 174) <= input(38);
output(0, 175) <= input(40);
output(0, 176) <= input(21);
output(0, 177) <= input(22);
output(0, 178) <= input(23);
output(0, 179) <= input(24);
output(0, 180) <= input(25);
output(0, 181) <= input(26);
output(0, 182) <= input(27);
output(0, 183) <= input(28);
output(0, 184) <= input(29);
output(0, 185) <= input(30);
output(0, 186) <= input(31);
output(0, 187) <= input(33);
output(0, 188) <= input(35);
output(0, 189) <= input(37);
output(0, 190) <= input(39);
output(0, 191) <= input(41);
output(0, 192) <= input(6);
output(0, 193) <= input(7);
output(0, 194) <= input(8);
output(0, 195) <= input(9);
output(0, 196) <= input(10);
output(0, 197) <= input(11);
output(0, 198) <= input(12);
output(0, 199) <= input(13);
output(0, 200) <= input(14);
output(0, 201) <= input(15);
output(0, 202) <= input(32);
output(0, 203) <= input(34);
output(0, 204) <= input(36);
output(0, 205) <= input(38);
output(0, 206) <= input(40);
output(0, 207) <= input(42);
output(0, 208) <= input(22);
output(0, 209) <= input(23);
output(0, 210) <= input(24);
output(0, 211) <= input(25);
output(0, 212) <= input(26);
output(0, 213) <= input(27);
output(0, 214) <= input(28);
output(0, 215) <= input(29);
output(0, 216) <= input(30);
output(0, 217) <= input(31);
output(0, 218) <= input(33);
output(0, 219) <= input(35);
output(0, 220) <= input(37);
output(0, 221) <= input(39);
output(0, 222) <= input(41);
output(0, 223) <= input(43);
output(0, 224) <= input(7);
output(0, 225) <= input(8);
output(0, 226) <= input(9);
output(0, 227) <= input(10);
output(0, 228) <= input(11);
output(0, 229) <= input(12);
output(0, 230) <= input(13);
output(0, 231) <= input(14);
output(0, 232) <= input(15);
output(0, 233) <= input(32);
output(0, 234) <= input(34);
output(0, 235) <= input(36);
output(0, 236) <= input(38);
output(0, 237) <= input(40);
output(0, 238) <= input(42);
output(0, 239) <= input(44);
output(0, 240) <= input(23);
output(0, 241) <= input(24);
output(0, 242) <= input(25);
output(0, 243) <= input(26);
output(0, 244) <= input(27);
output(0, 245) <= input(28);
output(0, 246) <= input(29);
output(0, 247) <= input(30);
output(0, 248) <= input(31);
output(0, 249) <= input(33);
output(0, 250) <= input(35);
output(0, 251) <= input(37);
output(0, 252) <= input(39);
output(0, 253) <= input(41);
output(0, 254) <= input(43);
output(0, 255) <= input(45);
output(1, 0) <= input(46);
output(1, 1) <= input(16);
output(1, 2) <= input(17);
output(1, 3) <= input(18);
output(1, 4) <= input(19);
output(1, 5) <= input(20);
output(1, 6) <= input(21);
output(1, 7) <= input(22);
output(1, 8) <= input(23);
output(1, 9) <= input(24);
output(1, 10) <= input(25);
output(1, 11) <= input(26);
output(1, 12) <= input(27);
output(1, 13) <= input(28);
output(1, 14) <= input(29);
output(1, 15) <= input(30);
output(1, 16) <= input(0);
output(1, 17) <= input(1);
output(1, 18) <= input(2);
output(1, 19) <= input(3);
output(1, 20) <= input(4);
output(1, 21) <= input(5);
output(1, 22) <= input(6);
output(1, 23) <= input(7);
output(1, 24) <= input(8);
output(1, 25) <= input(9);
output(1, 26) <= input(10);
output(1, 27) <= input(11);
output(1, 28) <= input(12);
output(1, 29) <= input(13);
output(1, 30) <= input(14);
output(1, 31) <= input(15);
output(1, 32) <= input(16);
output(1, 33) <= input(17);
output(1, 34) <= input(18);
output(1, 35) <= input(19);
output(1, 36) <= input(20);
output(1, 37) <= input(21);
output(1, 38) <= input(22);
output(1, 39) <= input(23);
output(1, 40) <= input(24);
output(1, 41) <= input(25);
output(1, 42) <= input(26);
output(1, 43) <= input(27);
output(1, 44) <= input(28);
output(1, 45) <= input(29);
output(1, 46) <= input(30);
output(1, 47) <= input(31);
output(1, 48) <= input(1);
output(1, 49) <= input(2);
output(1, 50) <= input(3);
output(1, 51) <= input(4);
output(1, 52) <= input(5);
output(1, 53) <= input(6);
output(1, 54) <= input(7);
output(1, 55) <= input(8);
output(1, 56) <= input(9);
output(1, 57) <= input(10);
output(1, 58) <= input(11);
output(1, 59) <= input(12);
output(1, 60) <= input(13);
output(1, 61) <= input(14);
output(1, 62) <= input(15);
output(1, 63) <= input(32);
output(1, 64) <= input(17);
output(1, 65) <= input(18);
output(1, 66) <= input(19);
output(1, 67) <= input(20);
output(1, 68) <= input(21);
output(1, 69) <= input(22);
output(1, 70) <= input(23);
output(1, 71) <= input(24);
output(1, 72) <= input(25);
output(1, 73) <= input(26);
output(1, 74) <= input(27);
output(1, 75) <= input(28);
output(1, 76) <= input(29);
output(1, 77) <= input(30);
output(1, 78) <= input(31);
output(1, 79) <= input(33);
output(1, 80) <= input(2);
output(1, 81) <= input(3);
output(1, 82) <= input(4);
output(1, 83) <= input(5);
output(1, 84) <= input(6);
output(1, 85) <= input(7);
output(1, 86) <= input(8);
output(1, 87) <= input(9);
output(1, 88) <= input(10);
output(1, 89) <= input(11);
output(1, 90) <= input(12);
output(1, 91) <= input(13);
output(1, 92) <= input(14);
output(1, 93) <= input(15);
output(1, 94) <= input(32);
output(1, 95) <= input(34);
output(1, 96) <= input(18);
output(1, 97) <= input(19);
output(1, 98) <= input(20);
output(1, 99) <= input(21);
output(1, 100) <= input(22);
output(1, 101) <= input(23);
output(1, 102) <= input(24);
output(1, 103) <= input(25);
output(1, 104) <= input(26);
output(1, 105) <= input(27);
output(1, 106) <= input(28);
output(1, 107) <= input(29);
output(1, 108) <= input(30);
output(1, 109) <= input(31);
output(1, 110) <= input(33);
output(1, 111) <= input(35);
output(1, 112) <= input(3);
output(1, 113) <= input(4);
output(1, 114) <= input(5);
output(1, 115) <= input(6);
output(1, 116) <= input(7);
output(1, 117) <= input(8);
output(1, 118) <= input(9);
output(1, 119) <= input(10);
output(1, 120) <= input(11);
output(1, 121) <= input(12);
output(1, 122) <= input(13);
output(1, 123) <= input(14);
output(1, 124) <= input(15);
output(1, 125) <= input(32);
output(1, 126) <= input(34);
output(1, 127) <= input(36);
output(1, 128) <= input(3);
output(1, 129) <= input(4);
output(1, 130) <= input(5);
output(1, 131) <= input(6);
output(1, 132) <= input(7);
output(1, 133) <= input(8);
output(1, 134) <= input(9);
output(1, 135) <= input(10);
output(1, 136) <= input(11);
output(1, 137) <= input(12);
output(1, 138) <= input(13);
output(1, 139) <= input(14);
output(1, 140) <= input(15);
output(1, 141) <= input(32);
output(1, 142) <= input(34);
output(1, 143) <= input(36);
output(1, 144) <= input(19);
output(1, 145) <= input(20);
output(1, 146) <= input(21);
output(1, 147) <= input(22);
output(1, 148) <= input(23);
output(1, 149) <= input(24);
output(1, 150) <= input(25);
output(1, 151) <= input(26);
output(1, 152) <= input(27);
output(1, 153) <= input(28);
output(1, 154) <= input(29);
output(1, 155) <= input(30);
output(1, 156) <= input(31);
output(1, 157) <= input(33);
output(1, 158) <= input(35);
output(1, 159) <= input(37);
output(1, 160) <= input(4);
output(1, 161) <= input(5);
output(1, 162) <= input(6);
output(1, 163) <= input(7);
output(1, 164) <= input(8);
output(1, 165) <= input(9);
output(1, 166) <= input(10);
output(1, 167) <= input(11);
output(1, 168) <= input(12);
output(1, 169) <= input(13);
output(1, 170) <= input(14);
output(1, 171) <= input(15);
output(1, 172) <= input(32);
output(1, 173) <= input(34);
output(1, 174) <= input(36);
output(1, 175) <= input(38);
output(1, 176) <= input(20);
output(1, 177) <= input(21);
output(1, 178) <= input(22);
output(1, 179) <= input(23);
output(1, 180) <= input(24);
output(1, 181) <= input(25);
output(1, 182) <= input(26);
output(1, 183) <= input(27);
output(1, 184) <= input(28);
output(1, 185) <= input(29);
output(1, 186) <= input(30);
output(1, 187) <= input(31);
output(1, 188) <= input(33);
output(1, 189) <= input(35);
output(1, 190) <= input(37);
output(1, 191) <= input(39);
output(1, 192) <= input(5);
output(1, 193) <= input(6);
output(1, 194) <= input(7);
output(1, 195) <= input(8);
output(1, 196) <= input(9);
output(1, 197) <= input(10);
output(1, 198) <= input(11);
output(1, 199) <= input(12);
output(1, 200) <= input(13);
output(1, 201) <= input(14);
output(1, 202) <= input(15);
output(1, 203) <= input(32);
output(1, 204) <= input(34);
output(1, 205) <= input(36);
output(1, 206) <= input(38);
output(1, 207) <= input(40);
output(1, 208) <= input(21);
output(1, 209) <= input(22);
output(1, 210) <= input(23);
output(1, 211) <= input(24);
output(1, 212) <= input(25);
output(1, 213) <= input(26);
output(1, 214) <= input(27);
output(1, 215) <= input(28);
output(1, 216) <= input(29);
output(1, 217) <= input(30);
output(1, 218) <= input(31);
output(1, 219) <= input(33);
output(1, 220) <= input(35);
output(1, 221) <= input(37);
output(1, 222) <= input(39);
output(1, 223) <= input(41);
output(1, 224) <= input(6);
output(1, 225) <= input(7);
output(1, 226) <= input(8);
output(1, 227) <= input(9);
output(1, 228) <= input(10);
output(1, 229) <= input(11);
output(1, 230) <= input(12);
output(1, 231) <= input(13);
output(1, 232) <= input(14);
output(1, 233) <= input(15);
output(1, 234) <= input(32);
output(1, 235) <= input(34);
output(1, 236) <= input(36);
output(1, 237) <= input(38);
output(1, 238) <= input(40);
output(1, 239) <= input(42);
output(1, 240) <= input(22);
output(1, 241) <= input(23);
output(1, 242) <= input(24);
output(1, 243) <= input(25);
output(1, 244) <= input(26);
output(1, 245) <= input(27);
output(1, 246) <= input(28);
output(1, 247) <= input(29);
output(1, 248) <= input(30);
output(1, 249) <= input(31);
output(1, 250) <= input(33);
output(1, 251) <= input(35);
output(1, 252) <= input(37);
output(1, 253) <= input(39);
output(1, 254) <= input(41);
output(1, 255) <= input(43);
output(2, 0) <= input(46);
output(2, 1) <= input(16);
output(2, 2) <= input(17);
output(2, 3) <= input(18);
output(2, 4) <= input(19);
output(2, 5) <= input(20);
output(2, 6) <= input(21);
output(2, 7) <= input(22);
output(2, 8) <= input(23);
output(2, 9) <= input(24);
output(2, 10) <= input(25);
output(2, 11) <= input(26);
output(2, 12) <= input(27);
output(2, 13) <= input(28);
output(2, 14) <= input(29);
output(2, 15) <= input(30);
output(2, 16) <= input(0);
output(2, 17) <= input(1);
output(2, 18) <= input(2);
output(2, 19) <= input(3);
output(2, 20) <= input(4);
output(2, 21) <= input(5);
output(2, 22) <= input(6);
output(2, 23) <= input(7);
output(2, 24) <= input(8);
output(2, 25) <= input(9);
output(2, 26) <= input(10);
output(2, 27) <= input(11);
output(2, 28) <= input(12);
output(2, 29) <= input(13);
output(2, 30) <= input(14);
output(2, 31) <= input(15);
output(2, 32) <= input(16);
output(2, 33) <= input(17);
output(2, 34) <= input(18);
output(2, 35) <= input(19);
output(2, 36) <= input(20);
output(2, 37) <= input(21);
output(2, 38) <= input(22);
output(2, 39) <= input(23);
output(2, 40) <= input(24);
output(2, 41) <= input(25);
output(2, 42) <= input(26);
output(2, 43) <= input(27);
output(2, 44) <= input(28);
output(2, 45) <= input(29);
output(2, 46) <= input(30);
output(2, 47) <= input(31);
output(2, 48) <= input(1);
output(2, 49) <= input(2);
output(2, 50) <= input(3);
output(2, 51) <= input(4);
output(2, 52) <= input(5);
output(2, 53) <= input(6);
output(2, 54) <= input(7);
output(2, 55) <= input(8);
output(2, 56) <= input(9);
output(2, 57) <= input(10);
output(2, 58) <= input(11);
output(2, 59) <= input(12);
output(2, 60) <= input(13);
output(2, 61) <= input(14);
output(2, 62) <= input(15);
output(2, 63) <= input(32);
output(2, 64) <= input(1);
output(2, 65) <= input(2);
output(2, 66) <= input(3);
output(2, 67) <= input(4);
output(2, 68) <= input(5);
output(2, 69) <= input(6);
output(2, 70) <= input(7);
output(2, 71) <= input(8);
output(2, 72) <= input(9);
output(2, 73) <= input(10);
output(2, 74) <= input(11);
output(2, 75) <= input(12);
output(2, 76) <= input(13);
output(2, 77) <= input(14);
output(2, 78) <= input(15);
output(2, 79) <= input(32);
output(2, 80) <= input(17);
output(2, 81) <= input(18);
output(2, 82) <= input(19);
output(2, 83) <= input(20);
output(2, 84) <= input(21);
output(2, 85) <= input(22);
output(2, 86) <= input(23);
output(2, 87) <= input(24);
output(2, 88) <= input(25);
output(2, 89) <= input(26);
output(2, 90) <= input(27);
output(2, 91) <= input(28);
output(2, 92) <= input(29);
output(2, 93) <= input(30);
output(2, 94) <= input(31);
output(2, 95) <= input(33);
output(2, 96) <= input(2);
output(2, 97) <= input(3);
output(2, 98) <= input(4);
output(2, 99) <= input(5);
output(2, 100) <= input(6);
output(2, 101) <= input(7);
output(2, 102) <= input(8);
output(2, 103) <= input(9);
output(2, 104) <= input(10);
output(2, 105) <= input(11);
output(2, 106) <= input(12);
output(2, 107) <= input(13);
output(2, 108) <= input(14);
output(2, 109) <= input(15);
output(2, 110) <= input(32);
output(2, 111) <= input(34);
output(2, 112) <= input(18);
output(2, 113) <= input(19);
output(2, 114) <= input(20);
output(2, 115) <= input(21);
output(2, 116) <= input(22);
output(2, 117) <= input(23);
output(2, 118) <= input(24);
output(2, 119) <= input(25);
output(2, 120) <= input(26);
output(2, 121) <= input(27);
output(2, 122) <= input(28);
output(2, 123) <= input(29);
output(2, 124) <= input(30);
output(2, 125) <= input(31);
output(2, 126) <= input(33);
output(2, 127) <= input(35);
output(2, 128) <= input(18);
output(2, 129) <= input(19);
output(2, 130) <= input(20);
output(2, 131) <= input(21);
output(2, 132) <= input(22);
output(2, 133) <= input(23);
output(2, 134) <= input(24);
output(2, 135) <= input(25);
output(2, 136) <= input(26);
output(2, 137) <= input(27);
output(2, 138) <= input(28);
output(2, 139) <= input(29);
output(2, 140) <= input(30);
output(2, 141) <= input(31);
output(2, 142) <= input(33);
output(2, 143) <= input(35);
output(2, 144) <= input(3);
output(2, 145) <= input(4);
output(2, 146) <= input(5);
output(2, 147) <= input(6);
output(2, 148) <= input(7);
output(2, 149) <= input(8);
output(2, 150) <= input(9);
output(2, 151) <= input(10);
output(2, 152) <= input(11);
output(2, 153) <= input(12);
output(2, 154) <= input(13);
output(2, 155) <= input(14);
output(2, 156) <= input(15);
output(2, 157) <= input(32);
output(2, 158) <= input(34);
output(2, 159) <= input(36);
output(2, 160) <= input(19);
output(2, 161) <= input(20);
output(2, 162) <= input(21);
output(2, 163) <= input(22);
output(2, 164) <= input(23);
output(2, 165) <= input(24);
output(2, 166) <= input(25);
output(2, 167) <= input(26);
output(2, 168) <= input(27);
output(2, 169) <= input(28);
output(2, 170) <= input(29);
output(2, 171) <= input(30);
output(2, 172) <= input(31);
output(2, 173) <= input(33);
output(2, 174) <= input(35);
output(2, 175) <= input(37);
output(2, 176) <= input(4);
output(2, 177) <= input(5);
output(2, 178) <= input(6);
output(2, 179) <= input(7);
output(2, 180) <= input(8);
output(2, 181) <= input(9);
output(2, 182) <= input(10);
output(2, 183) <= input(11);
output(2, 184) <= input(12);
output(2, 185) <= input(13);
output(2, 186) <= input(14);
output(2, 187) <= input(15);
output(2, 188) <= input(32);
output(2, 189) <= input(34);
output(2, 190) <= input(36);
output(2, 191) <= input(38);
output(2, 192) <= input(4);
output(2, 193) <= input(5);
output(2, 194) <= input(6);
output(2, 195) <= input(7);
output(2, 196) <= input(8);
output(2, 197) <= input(9);
output(2, 198) <= input(10);
output(2, 199) <= input(11);
output(2, 200) <= input(12);
output(2, 201) <= input(13);
output(2, 202) <= input(14);
output(2, 203) <= input(15);
output(2, 204) <= input(32);
output(2, 205) <= input(34);
output(2, 206) <= input(36);
output(2, 207) <= input(38);
output(2, 208) <= input(20);
output(2, 209) <= input(21);
output(2, 210) <= input(22);
output(2, 211) <= input(23);
output(2, 212) <= input(24);
output(2, 213) <= input(25);
output(2, 214) <= input(26);
output(2, 215) <= input(27);
output(2, 216) <= input(28);
output(2, 217) <= input(29);
output(2, 218) <= input(30);
output(2, 219) <= input(31);
output(2, 220) <= input(33);
output(2, 221) <= input(35);
output(2, 222) <= input(37);
output(2, 223) <= input(39);
output(2, 224) <= input(5);
output(2, 225) <= input(6);
output(2, 226) <= input(7);
output(2, 227) <= input(8);
output(2, 228) <= input(9);
output(2, 229) <= input(10);
output(2, 230) <= input(11);
output(2, 231) <= input(12);
output(2, 232) <= input(13);
output(2, 233) <= input(14);
output(2, 234) <= input(15);
output(2, 235) <= input(32);
output(2, 236) <= input(34);
output(2, 237) <= input(36);
output(2, 238) <= input(38);
output(2, 239) <= input(40);
output(2, 240) <= input(21);
output(2, 241) <= input(22);
output(2, 242) <= input(23);
output(2, 243) <= input(24);
output(2, 244) <= input(25);
output(2, 245) <= input(26);
output(2, 246) <= input(27);
output(2, 247) <= input(28);
output(2, 248) <= input(29);
output(2, 249) <= input(30);
output(2, 250) <= input(31);
output(2, 251) <= input(33);
output(2, 252) <= input(35);
output(2, 253) <= input(37);
output(2, 254) <= input(39);
output(2, 255) <= input(41);
output(3, 0) <= input(46);
output(3, 1) <= input(16);
output(3, 2) <= input(17);
output(3, 3) <= input(18);
output(3, 4) <= input(19);
output(3, 5) <= input(20);
output(3, 6) <= input(21);
output(3, 7) <= input(22);
output(3, 8) <= input(23);
output(3, 9) <= input(24);
output(3, 10) <= input(25);
output(3, 11) <= input(26);
output(3, 12) <= input(27);
output(3, 13) <= input(28);
output(3, 14) <= input(29);
output(3, 15) <= input(30);
output(3, 16) <= input(0);
output(3, 17) <= input(1);
output(3, 18) <= input(2);
output(3, 19) <= input(3);
output(3, 20) <= input(4);
output(3, 21) <= input(5);
output(3, 22) <= input(6);
output(3, 23) <= input(7);
output(3, 24) <= input(8);
output(3, 25) <= input(9);
output(3, 26) <= input(10);
output(3, 27) <= input(11);
output(3, 28) <= input(12);
output(3, 29) <= input(13);
output(3, 30) <= input(14);
output(3, 31) <= input(15);
output(3, 32) <= input(0);
output(3, 33) <= input(1);
output(3, 34) <= input(2);
output(3, 35) <= input(3);
output(3, 36) <= input(4);
output(3, 37) <= input(5);
output(3, 38) <= input(6);
output(3, 39) <= input(7);
output(3, 40) <= input(8);
output(3, 41) <= input(9);
output(3, 42) <= input(10);
output(3, 43) <= input(11);
output(3, 44) <= input(12);
output(3, 45) <= input(13);
output(3, 46) <= input(14);
output(3, 47) <= input(15);
output(3, 48) <= input(16);
output(3, 49) <= input(17);
output(3, 50) <= input(18);
output(3, 51) <= input(19);
output(3, 52) <= input(20);
output(3, 53) <= input(21);
output(3, 54) <= input(22);
output(3, 55) <= input(23);
output(3, 56) <= input(24);
output(3, 57) <= input(25);
output(3, 58) <= input(26);
output(3, 59) <= input(27);
output(3, 60) <= input(28);
output(3, 61) <= input(29);
output(3, 62) <= input(30);
output(3, 63) <= input(31);
output(3, 64) <= input(1);
output(3, 65) <= input(2);
output(3, 66) <= input(3);
output(3, 67) <= input(4);
output(3, 68) <= input(5);
output(3, 69) <= input(6);
output(3, 70) <= input(7);
output(3, 71) <= input(8);
output(3, 72) <= input(9);
output(3, 73) <= input(10);
output(3, 74) <= input(11);
output(3, 75) <= input(12);
output(3, 76) <= input(13);
output(3, 77) <= input(14);
output(3, 78) <= input(15);
output(3, 79) <= input(32);
output(3, 80) <= input(1);
output(3, 81) <= input(2);
output(3, 82) <= input(3);
output(3, 83) <= input(4);
output(3, 84) <= input(5);
output(3, 85) <= input(6);
output(3, 86) <= input(7);
output(3, 87) <= input(8);
output(3, 88) <= input(9);
output(3, 89) <= input(10);
output(3, 90) <= input(11);
output(3, 91) <= input(12);
output(3, 92) <= input(13);
output(3, 93) <= input(14);
output(3, 94) <= input(15);
output(3, 95) <= input(32);
output(3, 96) <= input(17);
output(3, 97) <= input(18);
output(3, 98) <= input(19);
output(3, 99) <= input(20);
output(3, 100) <= input(21);
output(3, 101) <= input(22);
output(3, 102) <= input(23);
output(3, 103) <= input(24);
output(3, 104) <= input(25);
output(3, 105) <= input(26);
output(3, 106) <= input(27);
output(3, 107) <= input(28);
output(3, 108) <= input(29);
output(3, 109) <= input(30);
output(3, 110) <= input(31);
output(3, 111) <= input(33);
output(3, 112) <= input(2);
output(3, 113) <= input(3);
output(3, 114) <= input(4);
output(3, 115) <= input(5);
output(3, 116) <= input(6);
output(3, 117) <= input(7);
output(3, 118) <= input(8);
output(3, 119) <= input(9);
output(3, 120) <= input(10);
output(3, 121) <= input(11);
output(3, 122) <= input(12);
output(3, 123) <= input(13);
output(3, 124) <= input(14);
output(3, 125) <= input(15);
output(3, 126) <= input(32);
output(3, 127) <= input(34);
output(3, 128) <= input(2);
output(3, 129) <= input(3);
output(3, 130) <= input(4);
output(3, 131) <= input(5);
output(3, 132) <= input(6);
output(3, 133) <= input(7);
output(3, 134) <= input(8);
output(3, 135) <= input(9);
output(3, 136) <= input(10);
output(3, 137) <= input(11);
output(3, 138) <= input(12);
output(3, 139) <= input(13);
output(3, 140) <= input(14);
output(3, 141) <= input(15);
output(3, 142) <= input(32);
output(3, 143) <= input(34);
output(3, 144) <= input(18);
output(3, 145) <= input(19);
output(3, 146) <= input(20);
output(3, 147) <= input(21);
output(3, 148) <= input(22);
output(3, 149) <= input(23);
output(3, 150) <= input(24);
output(3, 151) <= input(25);
output(3, 152) <= input(26);
output(3, 153) <= input(27);
output(3, 154) <= input(28);
output(3, 155) <= input(29);
output(3, 156) <= input(30);
output(3, 157) <= input(31);
output(3, 158) <= input(33);
output(3, 159) <= input(35);
output(3, 160) <= input(18);
output(3, 161) <= input(19);
output(3, 162) <= input(20);
output(3, 163) <= input(21);
output(3, 164) <= input(22);
output(3, 165) <= input(23);
output(3, 166) <= input(24);
output(3, 167) <= input(25);
output(3, 168) <= input(26);
output(3, 169) <= input(27);
output(3, 170) <= input(28);
output(3, 171) <= input(29);
output(3, 172) <= input(30);
output(3, 173) <= input(31);
output(3, 174) <= input(33);
output(3, 175) <= input(35);
output(3, 176) <= input(3);
output(3, 177) <= input(4);
output(3, 178) <= input(5);
output(3, 179) <= input(6);
output(3, 180) <= input(7);
output(3, 181) <= input(8);
output(3, 182) <= input(9);
output(3, 183) <= input(10);
output(3, 184) <= input(11);
output(3, 185) <= input(12);
output(3, 186) <= input(13);
output(3, 187) <= input(14);
output(3, 188) <= input(15);
output(3, 189) <= input(32);
output(3, 190) <= input(34);
output(3, 191) <= input(36);
output(3, 192) <= input(19);
output(3, 193) <= input(20);
output(3, 194) <= input(21);
output(3, 195) <= input(22);
output(3, 196) <= input(23);
output(3, 197) <= input(24);
output(3, 198) <= input(25);
output(3, 199) <= input(26);
output(3, 200) <= input(27);
output(3, 201) <= input(28);
output(3, 202) <= input(29);
output(3, 203) <= input(30);
output(3, 204) <= input(31);
output(3, 205) <= input(33);
output(3, 206) <= input(35);
output(3, 207) <= input(37);
output(3, 208) <= input(19);
output(3, 209) <= input(20);
output(3, 210) <= input(21);
output(3, 211) <= input(22);
output(3, 212) <= input(23);
output(3, 213) <= input(24);
output(3, 214) <= input(25);
output(3, 215) <= input(26);
output(3, 216) <= input(27);
output(3, 217) <= input(28);
output(3, 218) <= input(29);
output(3, 219) <= input(30);
output(3, 220) <= input(31);
output(3, 221) <= input(33);
output(3, 222) <= input(35);
output(3, 223) <= input(37);
output(3, 224) <= input(4);
output(3, 225) <= input(5);
output(3, 226) <= input(6);
output(3, 227) <= input(7);
output(3, 228) <= input(8);
output(3, 229) <= input(9);
output(3, 230) <= input(10);
output(3, 231) <= input(11);
output(3, 232) <= input(12);
output(3, 233) <= input(13);
output(3, 234) <= input(14);
output(3, 235) <= input(15);
output(3, 236) <= input(32);
output(3, 237) <= input(34);
output(3, 238) <= input(36);
output(3, 239) <= input(38);
output(3, 240) <= input(20);
output(3, 241) <= input(21);
output(3, 242) <= input(22);
output(3, 243) <= input(23);
output(3, 244) <= input(24);
output(3, 245) <= input(25);
output(3, 246) <= input(26);
output(3, 247) <= input(27);
output(3, 248) <= input(28);
output(3, 249) <= input(29);
output(3, 250) <= input(30);
output(3, 251) <= input(31);
output(3, 252) <= input(33);
output(3, 253) <= input(35);
output(3, 254) <= input(37);
output(3, 255) <= input(39);
output(4, 0) <= input(46);
output(4, 1) <= input(16);
output(4, 2) <= input(17);
output(4, 3) <= input(18);
output(4, 4) <= input(19);
output(4, 5) <= input(20);
output(4, 6) <= input(21);
output(4, 7) <= input(22);
output(4, 8) <= input(23);
output(4, 9) <= input(24);
output(4, 10) <= input(25);
output(4, 11) <= input(26);
output(4, 12) <= input(27);
output(4, 13) <= input(28);
output(4, 14) <= input(29);
output(4, 15) <= input(30);
output(4, 16) <= input(0);
output(4, 17) <= input(1);
output(4, 18) <= input(2);
output(4, 19) <= input(3);
output(4, 20) <= input(4);
output(4, 21) <= input(5);
output(4, 22) <= input(6);
output(4, 23) <= input(7);
output(4, 24) <= input(8);
output(4, 25) <= input(9);
output(4, 26) <= input(10);
output(4, 27) <= input(11);
output(4, 28) <= input(12);
output(4, 29) <= input(13);
output(4, 30) <= input(14);
output(4, 31) <= input(15);
output(4, 32) <= input(0);
output(4, 33) <= input(1);
output(4, 34) <= input(2);
output(4, 35) <= input(3);
output(4, 36) <= input(4);
output(4, 37) <= input(5);
output(4, 38) <= input(6);
output(4, 39) <= input(7);
output(4, 40) <= input(8);
output(4, 41) <= input(9);
output(4, 42) <= input(10);
output(4, 43) <= input(11);
output(4, 44) <= input(12);
output(4, 45) <= input(13);
output(4, 46) <= input(14);
output(4, 47) <= input(15);
output(4, 48) <= input(16);
output(4, 49) <= input(17);
output(4, 50) <= input(18);
output(4, 51) <= input(19);
output(4, 52) <= input(20);
output(4, 53) <= input(21);
output(4, 54) <= input(22);
output(4, 55) <= input(23);
output(4, 56) <= input(24);
output(4, 57) <= input(25);
output(4, 58) <= input(26);
output(4, 59) <= input(27);
output(4, 60) <= input(28);
output(4, 61) <= input(29);
output(4, 62) <= input(30);
output(4, 63) <= input(31);
output(4, 64) <= input(16);
output(4, 65) <= input(17);
output(4, 66) <= input(18);
output(4, 67) <= input(19);
output(4, 68) <= input(20);
output(4, 69) <= input(21);
output(4, 70) <= input(22);
output(4, 71) <= input(23);
output(4, 72) <= input(24);
output(4, 73) <= input(25);
output(4, 74) <= input(26);
output(4, 75) <= input(27);
output(4, 76) <= input(28);
output(4, 77) <= input(29);
output(4, 78) <= input(30);
output(4, 79) <= input(31);
output(4, 80) <= input(1);
output(4, 81) <= input(2);
output(4, 82) <= input(3);
output(4, 83) <= input(4);
output(4, 84) <= input(5);
output(4, 85) <= input(6);
output(4, 86) <= input(7);
output(4, 87) <= input(8);
output(4, 88) <= input(9);
output(4, 89) <= input(10);
output(4, 90) <= input(11);
output(4, 91) <= input(12);
output(4, 92) <= input(13);
output(4, 93) <= input(14);
output(4, 94) <= input(15);
output(4, 95) <= input(32);
output(4, 96) <= input(1);
output(4, 97) <= input(2);
output(4, 98) <= input(3);
output(4, 99) <= input(4);
output(4, 100) <= input(5);
output(4, 101) <= input(6);
output(4, 102) <= input(7);
output(4, 103) <= input(8);
output(4, 104) <= input(9);
output(4, 105) <= input(10);
output(4, 106) <= input(11);
output(4, 107) <= input(12);
output(4, 108) <= input(13);
output(4, 109) <= input(14);
output(4, 110) <= input(15);
output(4, 111) <= input(32);
output(4, 112) <= input(17);
output(4, 113) <= input(18);
output(4, 114) <= input(19);
output(4, 115) <= input(20);
output(4, 116) <= input(21);
output(4, 117) <= input(22);
output(4, 118) <= input(23);
output(4, 119) <= input(24);
output(4, 120) <= input(25);
output(4, 121) <= input(26);
output(4, 122) <= input(27);
output(4, 123) <= input(28);
output(4, 124) <= input(29);
output(4, 125) <= input(30);
output(4, 126) <= input(31);
output(4, 127) <= input(33);
output(4, 128) <= input(17);
output(4, 129) <= input(18);
output(4, 130) <= input(19);
output(4, 131) <= input(20);
output(4, 132) <= input(21);
output(4, 133) <= input(22);
output(4, 134) <= input(23);
output(4, 135) <= input(24);
output(4, 136) <= input(25);
output(4, 137) <= input(26);
output(4, 138) <= input(27);
output(4, 139) <= input(28);
output(4, 140) <= input(29);
output(4, 141) <= input(30);
output(4, 142) <= input(31);
output(4, 143) <= input(33);
output(4, 144) <= input(2);
output(4, 145) <= input(3);
output(4, 146) <= input(4);
output(4, 147) <= input(5);
output(4, 148) <= input(6);
output(4, 149) <= input(7);
output(4, 150) <= input(8);
output(4, 151) <= input(9);
output(4, 152) <= input(10);
output(4, 153) <= input(11);
output(4, 154) <= input(12);
output(4, 155) <= input(13);
output(4, 156) <= input(14);
output(4, 157) <= input(15);
output(4, 158) <= input(32);
output(4, 159) <= input(34);
output(4, 160) <= input(2);
output(4, 161) <= input(3);
output(4, 162) <= input(4);
output(4, 163) <= input(5);
output(4, 164) <= input(6);
output(4, 165) <= input(7);
output(4, 166) <= input(8);
output(4, 167) <= input(9);
output(4, 168) <= input(10);
output(4, 169) <= input(11);
output(4, 170) <= input(12);
output(4, 171) <= input(13);
output(4, 172) <= input(14);
output(4, 173) <= input(15);
output(4, 174) <= input(32);
output(4, 175) <= input(34);
output(4, 176) <= input(18);
output(4, 177) <= input(19);
output(4, 178) <= input(20);
output(4, 179) <= input(21);
output(4, 180) <= input(22);
output(4, 181) <= input(23);
output(4, 182) <= input(24);
output(4, 183) <= input(25);
output(4, 184) <= input(26);
output(4, 185) <= input(27);
output(4, 186) <= input(28);
output(4, 187) <= input(29);
output(4, 188) <= input(30);
output(4, 189) <= input(31);
output(4, 190) <= input(33);
output(4, 191) <= input(35);
output(4, 192) <= input(18);
output(4, 193) <= input(19);
output(4, 194) <= input(20);
output(4, 195) <= input(21);
output(4, 196) <= input(22);
output(4, 197) <= input(23);
output(4, 198) <= input(24);
output(4, 199) <= input(25);
output(4, 200) <= input(26);
output(4, 201) <= input(27);
output(4, 202) <= input(28);
output(4, 203) <= input(29);
output(4, 204) <= input(30);
output(4, 205) <= input(31);
output(4, 206) <= input(33);
output(4, 207) <= input(35);
output(4, 208) <= input(3);
output(4, 209) <= input(4);
output(4, 210) <= input(5);
output(4, 211) <= input(6);
output(4, 212) <= input(7);
output(4, 213) <= input(8);
output(4, 214) <= input(9);
output(4, 215) <= input(10);
output(4, 216) <= input(11);
output(4, 217) <= input(12);
output(4, 218) <= input(13);
output(4, 219) <= input(14);
output(4, 220) <= input(15);
output(4, 221) <= input(32);
output(4, 222) <= input(34);
output(4, 223) <= input(36);
output(4, 224) <= input(3);
output(4, 225) <= input(4);
output(4, 226) <= input(5);
output(4, 227) <= input(6);
output(4, 228) <= input(7);
output(4, 229) <= input(8);
output(4, 230) <= input(9);
output(4, 231) <= input(10);
output(4, 232) <= input(11);
output(4, 233) <= input(12);
output(4, 234) <= input(13);
output(4, 235) <= input(14);
output(4, 236) <= input(15);
output(4, 237) <= input(32);
output(4, 238) <= input(34);
output(4, 239) <= input(36);
output(4, 240) <= input(19);
output(4, 241) <= input(20);
output(4, 242) <= input(21);
output(4, 243) <= input(22);
output(4, 244) <= input(23);
output(4, 245) <= input(24);
output(4, 246) <= input(25);
output(4, 247) <= input(26);
output(4, 248) <= input(27);
output(4, 249) <= input(28);
output(4, 250) <= input(29);
output(4, 251) <= input(30);
output(4, 252) <= input(31);
output(4, 253) <= input(33);
output(4, 254) <= input(35);
output(4, 255) <= input(37);
output(5, 0) <= input(46);
output(5, 1) <= input(16);
output(5, 2) <= input(17);
output(5, 3) <= input(18);
output(5, 4) <= input(19);
output(5, 5) <= input(20);
output(5, 6) <= input(21);
output(5, 7) <= input(22);
output(5, 8) <= input(23);
output(5, 9) <= input(24);
output(5, 10) <= input(25);
output(5, 11) <= input(26);
output(5, 12) <= input(27);
output(5, 13) <= input(28);
output(5, 14) <= input(29);
output(5, 15) <= input(30);
output(5, 16) <= input(46);
output(5, 17) <= input(16);
output(5, 18) <= input(17);
output(5, 19) <= input(18);
output(5, 20) <= input(19);
output(5, 21) <= input(20);
output(5, 22) <= input(21);
output(5, 23) <= input(22);
output(5, 24) <= input(23);
output(5, 25) <= input(24);
output(5, 26) <= input(25);
output(5, 27) <= input(26);
output(5, 28) <= input(27);
output(5, 29) <= input(28);
output(5, 30) <= input(29);
output(5, 31) <= input(30);
output(5, 32) <= input(0);
output(5, 33) <= input(1);
output(5, 34) <= input(2);
output(5, 35) <= input(3);
output(5, 36) <= input(4);
output(5, 37) <= input(5);
output(5, 38) <= input(6);
output(5, 39) <= input(7);
output(5, 40) <= input(8);
output(5, 41) <= input(9);
output(5, 42) <= input(10);
output(5, 43) <= input(11);
output(5, 44) <= input(12);
output(5, 45) <= input(13);
output(5, 46) <= input(14);
output(5, 47) <= input(15);
output(5, 48) <= input(0);
output(5, 49) <= input(1);
output(5, 50) <= input(2);
output(5, 51) <= input(3);
output(5, 52) <= input(4);
output(5, 53) <= input(5);
output(5, 54) <= input(6);
output(5, 55) <= input(7);
output(5, 56) <= input(8);
output(5, 57) <= input(9);
output(5, 58) <= input(10);
output(5, 59) <= input(11);
output(5, 60) <= input(12);
output(5, 61) <= input(13);
output(5, 62) <= input(14);
output(5, 63) <= input(15);
output(5, 64) <= input(0);
output(5, 65) <= input(1);
output(5, 66) <= input(2);
output(5, 67) <= input(3);
output(5, 68) <= input(4);
output(5, 69) <= input(5);
output(5, 70) <= input(6);
output(5, 71) <= input(7);
output(5, 72) <= input(8);
output(5, 73) <= input(9);
output(5, 74) <= input(10);
output(5, 75) <= input(11);
output(5, 76) <= input(12);
output(5, 77) <= input(13);
output(5, 78) <= input(14);
output(5, 79) <= input(15);
output(5, 80) <= input(16);
output(5, 81) <= input(17);
output(5, 82) <= input(18);
output(5, 83) <= input(19);
output(5, 84) <= input(20);
output(5, 85) <= input(21);
output(5, 86) <= input(22);
output(5, 87) <= input(23);
output(5, 88) <= input(24);
output(5, 89) <= input(25);
output(5, 90) <= input(26);
output(5, 91) <= input(27);
output(5, 92) <= input(28);
output(5, 93) <= input(29);
output(5, 94) <= input(30);
output(5, 95) <= input(31);
output(5, 96) <= input(16);
output(5, 97) <= input(17);
output(5, 98) <= input(18);
output(5, 99) <= input(19);
output(5, 100) <= input(20);
output(5, 101) <= input(21);
output(5, 102) <= input(22);
output(5, 103) <= input(23);
output(5, 104) <= input(24);
output(5, 105) <= input(25);
output(5, 106) <= input(26);
output(5, 107) <= input(27);
output(5, 108) <= input(28);
output(5, 109) <= input(29);
output(5, 110) <= input(30);
output(5, 111) <= input(31);
output(5, 112) <= input(1);
output(5, 113) <= input(2);
output(5, 114) <= input(3);
output(5, 115) <= input(4);
output(5, 116) <= input(5);
output(5, 117) <= input(6);
output(5, 118) <= input(7);
output(5, 119) <= input(8);
output(5, 120) <= input(9);
output(5, 121) <= input(10);
output(5, 122) <= input(11);
output(5, 123) <= input(12);
output(5, 124) <= input(13);
output(5, 125) <= input(14);
output(5, 126) <= input(15);
output(5, 127) <= input(32);
output(5, 128) <= input(1);
output(5, 129) <= input(2);
output(5, 130) <= input(3);
output(5, 131) <= input(4);
output(5, 132) <= input(5);
output(5, 133) <= input(6);
output(5, 134) <= input(7);
output(5, 135) <= input(8);
output(5, 136) <= input(9);
output(5, 137) <= input(10);
output(5, 138) <= input(11);
output(5, 139) <= input(12);
output(5, 140) <= input(13);
output(5, 141) <= input(14);
output(5, 142) <= input(15);
output(5, 143) <= input(32);
output(5, 144) <= input(1);
output(5, 145) <= input(2);
output(5, 146) <= input(3);
output(5, 147) <= input(4);
output(5, 148) <= input(5);
output(5, 149) <= input(6);
output(5, 150) <= input(7);
output(5, 151) <= input(8);
output(5, 152) <= input(9);
output(5, 153) <= input(10);
output(5, 154) <= input(11);
output(5, 155) <= input(12);
output(5, 156) <= input(13);
output(5, 157) <= input(14);
output(5, 158) <= input(15);
output(5, 159) <= input(32);
output(5, 160) <= input(17);
output(5, 161) <= input(18);
output(5, 162) <= input(19);
output(5, 163) <= input(20);
output(5, 164) <= input(21);
output(5, 165) <= input(22);
output(5, 166) <= input(23);
output(5, 167) <= input(24);
output(5, 168) <= input(25);
output(5, 169) <= input(26);
output(5, 170) <= input(27);
output(5, 171) <= input(28);
output(5, 172) <= input(29);
output(5, 173) <= input(30);
output(5, 174) <= input(31);
output(5, 175) <= input(33);
output(5, 176) <= input(17);
output(5, 177) <= input(18);
output(5, 178) <= input(19);
output(5, 179) <= input(20);
output(5, 180) <= input(21);
output(5, 181) <= input(22);
output(5, 182) <= input(23);
output(5, 183) <= input(24);
output(5, 184) <= input(25);
output(5, 185) <= input(26);
output(5, 186) <= input(27);
output(5, 187) <= input(28);
output(5, 188) <= input(29);
output(5, 189) <= input(30);
output(5, 190) <= input(31);
output(5, 191) <= input(33);
output(5, 192) <= input(17);
output(5, 193) <= input(18);
output(5, 194) <= input(19);
output(5, 195) <= input(20);
output(5, 196) <= input(21);
output(5, 197) <= input(22);
output(5, 198) <= input(23);
output(5, 199) <= input(24);
output(5, 200) <= input(25);
output(5, 201) <= input(26);
output(5, 202) <= input(27);
output(5, 203) <= input(28);
output(5, 204) <= input(29);
output(5, 205) <= input(30);
output(5, 206) <= input(31);
output(5, 207) <= input(33);
output(5, 208) <= input(2);
output(5, 209) <= input(3);
output(5, 210) <= input(4);
output(5, 211) <= input(5);
output(5, 212) <= input(6);
output(5, 213) <= input(7);
output(5, 214) <= input(8);
output(5, 215) <= input(9);
output(5, 216) <= input(10);
output(5, 217) <= input(11);
output(5, 218) <= input(12);
output(5, 219) <= input(13);
output(5, 220) <= input(14);
output(5, 221) <= input(15);
output(5, 222) <= input(32);
output(5, 223) <= input(34);
output(5, 224) <= input(2);
output(5, 225) <= input(3);
output(5, 226) <= input(4);
output(5, 227) <= input(5);
output(5, 228) <= input(6);
output(5, 229) <= input(7);
output(5, 230) <= input(8);
output(5, 231) <= input(9);
output(5, 232) <= input(10);
output(5, 233) <= input(11);
output(5, 234) <= input(12);
output(5, 235) <= input(13);
output(5, 236) <= input(14);
output(5, 237) <= input(15);
output(5, 238) <= input(32);
output(5, 239) <= input(34);
output(5, 240) <= input(18);
output(5, 241) <= input(19);
output(5, 242) <= input(20);
output(5, 243) <= input(21);
output(5, 244) <= input(22);
output(5, 245) <= input(23);
output(5, 246) <= input(24);
output(5, 247) <= input(25);
output(5, 248) <= input(26);
output(5, 249) <= input(27);
output(5, 250) <= input(28);
output(5, 251) <= input(29);
output(5, 252) <= input(30);
output(5, 253) <= input(31);
output(5, 254) <= input(33);
output(5, 255) <= input(35);
when "0010" =>
output(0, 0) <= input(0);
output(0, 1) <= input(1);
output(0, 2) <= input(2);
output(0, 3) <= input(3);
output(0, 4) <= input(4);
output(0, 5) <= input(5);
output(0, 6) <= input(6);
output(0, 7) <= input(7);
output(0, 8) <= input(8);
output(0, 9) <= input(9);
output(0, 10) <= input(10);
output(0, 11) <= input(11);
output(0, 12) <= input(12);
output(0, 13) <= input(13);
output(0, 14) <= input(14);
output(0, 15) <= input(15);
output(0, 16) <= input(0);
output(0, 17) <= input(1);
output(0, 18) <= input(2);
output(0, 19) <= input(3);
output(0, 20) <= input(4);
output(0, 21) <= input(5);
output(0, 22) <= input(6);
output(0, 23) <= input(7);
output(0, 24) <= input(8);
output(0, 25) <= input(9);
output(0, 26) <= input(10);
output(0, 27) <= input(11);
output(0, 28) <= input(12);
output(0, 29) <= input(13);
output(0, 30) <= input(14);
output(0, 31) <= input(15);
output(0, 32) <= input(0);
output(0, 33) <= input(1);
output(0, 34) <= input(2);
output(0, 35) <= input(3);
output(0, 36) <= input(4);
output(0, 37) <= input(5);
output(0, 38) <= input(6);
output(0, 39) <= input(7);
output(0, 40) <= input(8);
output(0, 41) <= input(9);
output(0, 42) <= input(10);
output(0, 43) <= input(11);
output(0, 44) <= input(12);
output(0, 45) <= input(13);
output(0, 46) <= input(14);
output(0, 47) <= input(15);
output(0, 48) <= input(16);
output(0, 49) <= input(17);
output(0, 50) <= input(18);
output(0, 51) <= input(19);
output(0, 52) <= input(20);
output(0, 53) <= input(21);
output(0, 54) <= input(22);
output(0, 55) <= input(23);
output(0, 56) <= input(24);
output(0, 57) <= input(25);
output(0, 58) <= input(26);
output(0, 59) <= input(27);
output(0, 60) <= input(28);
output(0, 61) <= input(29);
output(0, 62) <= input(30);
output(0, 63) <= input(31);
output(0, 64) <= input(16);
output(0, 65) <= input(17);
output(0, 66) <= input(18);
output(0, 67) <= input(19);
output(0, 68) <= input(20);
output(0, 69) <= input(21);
output(0, 70) <= input(22);
output(0, 71) <= input(23);
output(0, 72) <= input(24);
output(0, 73) <= input(25);
output(0, 74) <= input(26);
output(0, 75) <= input(27);
output(0, 76) <= input(28);
output(0, 77) <= input(29);
output(0, 78) <= input(30);
output(0, 79) <= input(31);
output(0, 80) <= input(16);
output(0, 81) <= input(17);
output(0, 82) <= input(18);
output(0, 83) <= input(19);
output(0, 84) <= input(20);
output(0, 85) <= input(21);
output(0, 86) <= input(22);
output(0, 87) <= input(23);
output(0, 88) <= input(24);
output(0, 89) <= input(25);
output(0, 90) <= input(26);
output(0, 91) <= input(27);
output(0, 92) <= input(28);
output(0, 93) <= input(29);
output(0, 94) <= input(30);
output(0, 95) <= input(31);
output(0, 96) <= input(16);
output(0, 97) <= input(17);
output(0, 98) <= input(18);
output(0, 99) <= input(19);
output(0, 100) <= input(20);
output(0, 101) <= input(21);
output(0, 102) <= input(22);
output(0, 103) <= input(23);
output(0, 104) <= input(24);
output(0, 105) <= input(25);
output(0, 106) <= input(26);
output(0, 107) <= input(27);
output(0, 108) <= input(28);
output(0, 109) <= input(29);
output(0, 110) <= input(30);
output(0, 111) <= input(31);
output(0, 112) <= input(1);
output(0, 113) <= input(2);
output(0, 114) <= input(3);
output(0, 115) <= input(4);
output(0, 116) <= input(5);
output(0, 117) <= input(6);
output(0, 118) <= input(7);
output(0, 119) <= input(8);
output(0, 120) <= input(9);
output(0, 121) <= input(10);
output(0, 122) <= input(11);
output(0, 123) <= input(12);
output(0, 124) <= input(13);
output(0, 125) <= input(14);
output(0, 126) <= input(15);
output(0, 127) <= input(32);
output(0, 128) <= input(1);
output(0, 129) <= input(2);
output(0, 130) <= input(3);
output(0, 131) <= input(4);
output(0, 132) <= input(5);
output(0, 133) <= input(6);
output(0, 134) <= input(7);
output(0, 135) <= input(8);
output(0, 136) <= input(9);
output(0, 137) <= input(10);
output(0, 138) <= input(11);
output(0, 139) <= input(12);
output(0, 140) <= input(13);
output(0, 141) <= input(14);
output(0, 142) <= input(15);
output(0, 143) <= input(32);
output(0, 144) <= input(1);
output(0, 145) <= input(2);
output(0, 146) <= input(3);
output(0, 147) <= input(4);
output(0, 148) <= input(5);
output(0, 149) <= input(6);
output(0, 150) <= input(7);
output(0, 151) <= input(8);
output(0, 152) <= input(9);
output(0, 153) <= input(10);
output(0, 154) <= input(11);
output(0, 155) <= input(12);
output(0, 156) <= input(13);
output(0, 157) <= input(14);
output(0, 158) <= input(15);
output(0, 159) <= input(32);
output(0, 160) <= input(1);
output(0, 161) <= input(2);
output(0, 162) <= input(3);
output(0, 163) <= input(4);
output(0, 164) <= input(5);
output(0, 165) <= input(6);
output(0, 166) <= input(7);
output(0, 167) <= input(8);
output(0, 168) <= input(9);
output(0, 169) <= input(10);
output(0, 170) <= input(11);
output(0, 171) <= input(12);
output(0, 172) <= input(13);
output(0, 173) <= input(14);
output(0, 174) <= input(15);
output(0, 175) <= input(32);
output(0, 176) <= input(17);
output(0, 177) <= input(18);
output(0, 178) <= input(19);
output(0, 179) <= input(20);
output(0, 180) <= input(21);
output(0, 181) <= input(22);
output(0, 182) <= input(23);
output(0, 183) <= input(24);
output(0, 184) <= input(25);
output(0, 185) <= input(26);
output(0, 186) <= input(27);
output(0, 187) <= input(28);
output(0, 188) <= input(29);
output(0, 189) <= input(30);
output(0, 190) <= input(31);
output(0, 191) <= input(33);
output(0, 192) <= input(17);
output(0, 193) <= input(18);
output(0, 194) <= input(19);
output(0, 195) <= input(20);
output(0, 196) <= input(21);
output(0, 197) <= input(22);
output(0, 198) <= input(23);
output(0, 199) <= input(24);
output(0, 200) <= input(25);
output(0, 201) <= input(26);
output(0, 202) <= input(27);
output(0, 203) <= input(28);
output(0, 204) <= input(29);
output(0, 205) <= input(30);
output(0, 206) <= input(31);
output(0, 207) <= input(33);
output(0, 208) <= input(17);
output(0, 209) <= input(18);
output(0, 210) <= input(19);
output(0, 211) <= input(20);
output(0, 212) <= input(21);
output(0, 213) <= input(22);
output(0, 214) <= input(23);
output(0, 215) <= input(24);
output(0, 216) <= input(25);
output(0, 217) <= input(26);
output(0, 218) <= input(27);
output(0, 219) <= input(28);
output(0, 220) <= input(29);
output(0, 221) <= input(30);
output(0, 222) <= input(31);
output(0, 223) <= input(33);
output(0, 224) <= input(17);
output(0, 225) <= input(18);
output(0, 226) <= input(19);
output(0, 227) <= input(20);
output(0, 228) <= input(21);
output(0, 229) <= input(22);
output(0, 230) <= input(23);
output(0, 231) <= input(24);
output(0, 232) <= input(25);
output(0, 233) <= input(26);
output(0, 234) <= input(27);
output(0, 235) <= input(28);
output(0, 236) <= input(29);
output(0, 237) <= input(30);
output(0, 238) <= input(31);
output(0, 239) <= input(33);
output(0, 240) <= input(2);
output(0, 241) <= input(3);
output(0, 242) <= input(4);
output(0, 243) <= input(5);
output(0, 244) <= input(6);
output(0, 245) <= input(7);
output(0, 246) <= input(8);
output(0, 247) <= input(9);
output(0, 248) <= input(10);
output(0, 249) <= input(11);
output(0, 250) <= input(12);
output(0, 251) <= input(13);
output(0, 252) <= input(14);
output(0, 253) <= input(15);
output(0, 254) <= input(32);
output(0, 255) <= input(34);
output(1, 0) <= input(0);
output(1, 1) <= input(1);
output(1, 2) <= input(2);
output(1, 3) <= input(3);
output(1, 4) <= input(4);
output(1, 5) <= input(5);
output(1, 6) <= input(6);
output(1, 7) <= input(7);
output(1, 8) <= input(8);
output(1, 9) <= input(9);
output(1, 10) <= input(10);
output(1, 11) <= input(11);
output(1, 12) <= input(12);
output(1, 13) <= input(13);
output(1, 14) <= input(14);
output(1, 15) <= input(15);
output(1, 16) <= input(0);
output(1, 17) <= input(1);
output(1, 18) <= input(2);
output(1, 19) <= input(3);
output(1, 20) <= input(4);
output(1, 21) <= input(5);
output(1, 22) <= input(6);
output(1, 23) <= input(7);
output(1, 24) <= input(8);
output(1, 25) <= input(9);
output(1, 26) <= input(10);
output(1, 27) <= input(11);
output(1, 28) <= input(12);
output(1, 29) <= input(13);
output(1, 30) <= input(14);
output(1, 31) <= input(15);
output(1, 32) <= input(0);
output(1, 33) <= input(1);
output(1, 34) <= input(2);
output(1, 35) <= input(3);
output(1, 36) <= input(4);
output(1, 37) <= input(5);
output(1, 38) <= input(6);
output(1, 39) <= input(7);
output(1, 40) <= input(8);
output(1, 41) <= input(9);
output(1, 42) <= input(10);
output(1, 43) <= input(11);
output(1, 44) <= input(12);
output(1, 45) <= input(13);
output(1, 46) <= input(14);
output(1, 47) <= input(15);
output(1, 48) <= input(0);
output(1, 49) <= input(1);
output(1, 50) <= input(2);
output(1, 51) <= input(3);
output(1, 52) <= input(4);
output(1, 53) <= input(5);
output(1, 54) <= input(6);
output(1, 55) <= input(7);
output(1, 56) <= input(8);
output(1, 57) <= input(9);
output(1, 58) <= input(10);
output(1, 59) <= input(11);
output(1, 60) <= input(12);
output(1, 61) <= input(13);
output(1, 62) <= input(14);
output(1, 63) <= input(15);
output(1, 64) <= input(0);
output(1, 65) <= input(1);
output(1, 66) <= input(2);
output(1, 67) <= input(3);
output(1, 68) <= input(4);
output(1, 69) <= input(5);
output(1, 70) <= input(6);
output(1, 71) <= input(7);
output(1, 72) <= input(8);
output(1, 73) <= input(9);
output(1, 74) <= input(10);
output(1, 75) <= input(11);
output(1, 76) <= input(12);
output(1, 77) <= input(13);
output(1, 78) <= input(14);
output(1, 79) <= input(15);
output(1, 80) <= input(16);
output(1, 81) <= input(17);
output(1, 82) <= input(18);
output(1, 83) <= input(19);
output(1, 84) <= input(20);
output(1, 85) <= input(21);
output(1, 86) <= input(22);
output(1, 87) <= input(23);
output(1, 88) <= input(24);
output(1, 89) <= input(25);
output(1, 90) <= input(26);
output(1, 91) <= input(27);
output(1, 92) <= input(28);
output(1, 93) <= input(29);
output(1, 94) <= input(30);
output(1, 95) <= input(31);
output(1, 96) <= input(16);
output(1, 97) <= input(17);
output(1, 98) <= input(18);
output(1, 99) <= input(19);
output(1, 100) <= input(20);
output(1, 101) <= input(21);
output(1, 102) <= input(22);
output(1, 103) <= input(23);
output(1, 104) <= input(24);
output(1, 105) <= input(25);
output(1, 106) <= input(26);
output(1, 107) <= input(27);
output(1, 108) <= input(28);
output(1, 109) <= input(29);
output(1, 110) <= input(30);
output(1, 111) <= input(31);
output(1, 112) <= input(16);
output(1, 113) <= input(17);
output(1, 114) <= input(18);
output(1, 115) <= input(19);
output(1, 116) <= input(20);
output(1, 117) <= input(21);
output(1, 118) <= input(22);
output(1, 119) <= input(23);
output(1, 120) <= input(24);
output(1, 121) <= input(25);
output(1, 122) <= input(26);
output(1, 123) <= input(27);
output(1, 124) <= input(28);
output(1, 125) <= input(29);
output(1, 126) <= input(30);
output(1, 127) <= input(31);
output(1, 128) <= input(16);
output(1, 129) <= input(17);
output(1, 130) <= input(18);
output(1, 131) <= input(19);
output(1, 132) <= input(20);
output(1, 133) <= input(21);
output(1, 134) <= input(22);
output(1, 135) <= input(23);
output(1, 136) <= input(24);
output(1, 137) <= input(25);
output(1, 138) <= input(26);
output(1, 139) <= input(27);
output(1, 140) <= input(28);
output(1, 141) <= input(29);
output(1, 142) <= input(30);
output(1, 143) <= input(31);
output(1, 144) <= input(16);
output(1, 145) <= input(17);
output(1, 146) <= input(18);
output(1, 147) <= input(19);
output(1, 148) <= input(20);
output(1, 149) <= input(21);
output(1, 150) <= input(22);
output(1, 151) <= input(23);
output(1, 152) <= input(24);
output(1, 153) <= input(25);
output(1, 154) <= input(26);
output(1, 155) <= input(27);
output(1, 156) <= input(28);
output(1, 157) <= input(29);
output(1, 158) <= input(30);
output(1, 159) <= input(31);
output(1, 160) <= input(1);
output(1, 161) <= input(2);
output(1, 162) <= input(3);
output(1, 163) <= input(4);
output(1, 164) <= input(5);
output(1, 165) <= input(6);
output(1, 166) <= input(7);
output(1, 167) <= input(8);
output(1, 168) <= input(9);
output(1, 169) <= input(10);
output(1, 170) <= input(11);
output(1, 171) <= input(12);
output(1, 172) <= input(13);
output(1, 173) <= input(14);
output(1, 174) <= input(15);
output(1, 175) <= input(32);
output(1, 176) <= input(1);
output(1, 177) <= input(2);
output(1, 178) <= input(3);
output(1, 179) <= input(4);
output(1, 180) <= input(5);
output(1, 181) <= input(6);
output(1, 182) <= input(7);
output(1, 183) <= input(8);
output(1, 184) <= input(9);
output(1, 185) <= input(10);
output(1, 186) <= input(11);
output(1, 187) <= input(12);
output(1, 188) <= input(13);
output(1, 189) <= input(14);
output(1, 190) <= input(15);
output(1, 191) <= input(32);
output(1, 192) <= input(1);
output(1, 193) <= input(2);
output(1, 194) <= input(3);
output(1, 195) <= input(4);
output(1, 196) <= input(5);
output(1, 197) <= input(6);
output(1, 198) <= input(7);
output(1, 199) <= input(8);
output(1, 200) <= input(9);
output(1, 201) <= input(10);
output(1, 202) <= input(11);
output(1, 203) <= input(12);
output(1, 204) <= input(13);
output(1, 205) <= input(14);
output(1, 206) <= input(15);
output(1, 207) <= input(32);
output(1, 208) <= input(1);
output(1, 209) <= input(2);
output(1, 210) <= input(3);
output(1, 211) <= input(4);
output(1, 212) <= input(5);
output(1, 213) <= input(6);
output(1, 214) <= input(7);
output(1, 215) <= input(8);
output(1, 216) <= input(9);
output(1, 217) <= input(10);
output(1, 218) <= input(11);
output(1, 219) <= input(12);
output(1, 220) <= input(13);
output(1, 221) <= input(14);
output(1, 222) <= input(15);
output(1, 223) <= input(32);
output(1, 224) <= input(1);
output(1, 225) <= input(2);
output(1, 226) <= input(3);
output(1, 227) <= input(4);
output(1, 228) <= input(5);
output(1, 229) <= input(6);
output(1, 230) <= input(7);
output(1, 231) <= input(8);
output(1, 232) <= input(9);
output(1, 233) <= input(10);
output(1, 234) <= input(11);
output(1, 235) <= input(12);
output(1, 236) <= input(13);
output(1, 237) <= input(14);
output(1, 238) <= input(15);
output(1, 239) <= input(32);
output(1, 240) <= input(17);
output(1, 241) <= input(18);
output(1, 242) <= input(19);
output(1, 243) <= input(20);
output(1, 244) <= input(21);
output(1, 245) <= input(22);
output(1, 246) <= input(23);
output(1, 247) <= input(24);
output(1, 248) <= input(25);
output(1, 249) <= input(26);
output(1, 250) <= input(27);
output(1, 251) <= input(28);
output(1, 252) <= input(29);
output(1, 253) <= input(30);
output(1, 254) <= input(31);
output(1, 255) <= input(33);
output(2, 0) <= input(0);
output(2, 1) <= input(1);
output(2, 2) <= input(2);
output(2, 3) <= input(3);
output(2, 4) <= input(4);
output(2, 5) <= input(5);
output(2, 6) <= input(6);
output(2, 7) <= input(7);
output(2, 8) <= input(8);
output(2, 9) <= input(9);
output(2, 10) <= input(10);
output(2, 11) <= input(11);
output(2, 12) <= input(12);
output(2, 13) <= input(13);
output(2, 14) <= input(14);
output(2, 15) <= input(15);
output(2, 16) <= input(0);
output(2, 17) <= input(1);
output(2, 18) <= input(2);
output(2, 19) <= input(3);
output(2, 20) <= input(4);
output(2, 21) <= input(5);
output(2, 22) <= input(6);
output(2, 23) <= input(7);
output(2, 24) <= input(8);
output(2, 25) <= input(9);
output(2, 26) <= input(10);
output(2, 27) <= input(11);
output(2, 28) <= input(12);
output(2, 29) <= input(13);
output(2, 30) <= input(14);
output(2, 31) <= input(15);
output(2, 32) <= input(0);
output(2, 33) <= input(1);
output(2, 34) <= input(2);
output(2, 35) <= input(3);
output(2, 36) <= input(4);
output(2, 37) <= input(5);
output(2, 38) <= input(6);
output(2, 39) <= input(7);
output(2, 40) <= input(8);
output(2, 41) <= input(9);
output(2, 42) <= input(10);
output(2, 43) <= input(11);
output(2, 44) <= input(12);
output(2, 45) <= input(13);
output(2, 46) <= input(14);
output(2, 47) <= input(15);
output(2, 48) <= input(0);
output(2, 49) <= input(1);
output(2, 50) <= input(2);
output(2, 51) <= input(3);
output(2, 52) <= input(4);
output(2, 53) <= input(5);
output(2, 54) <= input(6);
output(2, 55) <= input(7);
output(2, 56) <= input(8);
output(2, 57) <= input(9);
output(2, 58) <= input(10);
output(2, 59) <= input(11);
output(2, 60) <= input(12);
output(2, 61) <= input(13);
output(2, 62) <= input(14);
output(2, 63) <= input(15);
output(2, 64) <= input(0);
output(2, 65) <= input(1);
output(2, 66) <= input(2);
output(2, 67) <= input(3);
output(2, 68) <= input(4);
output(2, 69) <= input(5);
output(2, 70) <= input(6);
output(2, 71) <= input(7);
output(2, 72) <= input(8);
output(2, 73) <= input(9);
output(2, 74) <= input(10);
output(2, 75) <= input(11);
output(2, 76) <= input(12);
output(2, 77) <= input(13);
output(2, 78) <= input(14);
output(2, 79) <= input(15);
output(2, 80) <= input(0);
output(2, 81) <= input(1);
output(2, 82) <= input(2);
output(2, 83) <= input(3);
output(2, 84) <= input(4);
output(2, 85) <= input(5);
output(2, 86) <= input(6);
output(2, 87) <= input(7);
output(2, 88) <= input(8);
output(2, 89) <= input(9);
output(2, 90) <= input(10);
output(2, 91) <= input(11);
output(2, 92) <= input(12);
output(2, 93) <= input(13);
output(2, 94) <= input(14);
output(2, 95) <= input(15);
output(2, 96) <= input(0);
output(2, 97) <= input(1);
output(2, 98) <= input(2);
output(2, 99) <= input(3);
output(2, 100) <= input(4);
output(2, 101) <= input(5);
output(2, 102) <= input(6);
output(2, 103) <= input(7);
output(2, 104) <= input(8);
output(2, 105) <= input(9);
output(2, 106) <= input(10);
output(2, 107) <= input(11);
output(2, 108) <= input(12);
output(2, 109) <= input(13);
output(2, 110) <= input(14);
output(2, 111) <= input(15);
output(2, 112) <= input(16);
output(2, 113) <= input(17);
output(2, 114) <= input(18);
output(2, 115) <= input(19);
output(2, 116) <= input(20);
output(2, 117) <= input(21);
output(2, 118) <= input(22);
output(2, 119) <= input(23);
output(2, 120) <= input(24);
output(2, 121) <= input(25);
output(2, 122) <= input(26);
output(2, 123) <= input(27);
output(2, 124) <= input(28);
output(2, 125) <= input(29);
output(2, 126) <= input(30);
output(2, 127) <= input(31);
output(2, 128) <= input(16);
output(2, 129) <= input(17);
output(2, 130) <= input(18);
output(2, 131) <= input(19);
output(2, 132) <= input(20);
output(2, 133) <= input(21);
output(2, 134) <= input(22);
output(2, 135) <= input(23);
output(2, 136) <= input(24);
output(2, 137) <= input(25);
output(2, 138) <= input(26);
output(2, 139) <= input(27);
output(2, 140) <= input(28);
output(2, 141) <= input(29);
output(2, 142) <= input(30);
output(2, 143) <= input(31);
output(2, 144) <= input(16);
output(2, 145) <= input(17);
output(2, 146) <= input(18);
output(2, 147) <= input(19);
output(2, 148) <= input(20);
output(2, 149) <= input(21);
output(2, 150) <= input(22);
output(2, 151) <= input(23);
output(2, 152) <= input(24);
output(2, 153) <= input(25);
output(2, 154) <= input(26);
output(2, 155) <= input(27);
output(2, 156) <= input(28);
output(2, 157) <= input(29);
output(2, 158) <= input(30);
output(2, 159) <= input(31);
output(2, 160) <= input(16);
output(2, 161) <= input(17);
output(2, 162) <= input(18);
output(2, 163) <= input(19);
output(2, 164) <= input(20);
output(2, 165) <= input(21);
output(2, 166) <= input(22);
output(2, 167) <= input(23);
output(2, 168) <= input(24);
output(2, 169) <= input(25);
output(2, 170) <= input(26);
output(2, 171) <= input(27);
output(2, 172) <= input(28);
output(2, 173) <= input(29);
output(2, 174) <= input(30);
output(2, 175) <= input(31);
output(2, 176) <= input(16);
output(2, 177) <= input(17);
output(2, 178) <= input(18);
output(2, 179) <= input(19);
output(2, 180) <= input(20);
output(2, 181) <= input(21);
output(2, 182) <= input(22);
output(2, 183) <= input(23);
output(2, 184) <= input(24);
output(2, 185) <= input(25);
output(2, 186) <= input(26);
output(2, 187) <= input(27);
output(2, 188) <= input(28);
output(2, 189) <= input(29);
output(2, 190) <= input(30);
output(2, 191) <= input(31);
output(2, 192) <= input(16);
output(2, 193) <= input(17);
output(2, 194) <= input(18);
output(2, 195) <= input(19);
output(2, 196) <= input(20);
output(2, 197) <= input(21);
output(2, 198) <= input(22);
output(2, 199) <= input(23);
output(2, 200) <= input(24);
output(2, 201) <= input(25);
output(2, 202) <= input(26);
output(2, 203) <= input(27);
output(2, 204) <= input(28);
output(2, 205) <= input(29);
output(2, 206) <= input(30);
output(2, 207) <= input(31);
output(2, 208) <= input(16);
output(2, 209) <= input(17);
output(2, 210) <= input(18);
output(2, 211) <= input(19);
output(2, 212) <= input(20);
output(2, 213) <= input(21);
output(2, 214) <= input(22);
output(2, 215) <= input(23);
output(2, 216) <= input(24);
output(2, 217) <= input(25);
output(2, 218) <= input(26);
output(2, 219) <= input(27);
output(2, 220) <= input(28);
output(2, 221) <= input(29);
output(2, 222) <= input(30);
output(2, 223) <= input(31);
output(2, 224) <= input(16);
output(2, 225) <= input(17);
output(2, 226) <= input(18);
output(2, 227) <= input(19);
output(2, 228) <= input(20);
output(2, 229) <= input(21);
output(2, 230) <= input(22);
output(2, 231) <= input(23);
output(2, 232) <= input(24);
output(2, 233) <= input(25);
output(2, 234) <= input(26);
output(2, 235) <= input(27);
output(2, 236) <= input(28);
output(2, 237) <= input(29);
output(2, 238) <= input(30);
output(2, 239) <= input(31);
output(2, 240) <= input(1);
output(2, 241) <= input(2);
output(2, 242) <= input(3);
output(2, 243) <= input(4);
output(2, 244) <= input(5);
output(2, 245) <= input(6);
output(2, 246) <= input(7);
output(2, 247) <= input(8);
output(2, 248) <= input(9);
output(2, 249) <= input(10);
output(2, 250) <= input(11);
output(2, 251) <= input(12);
output(2, 252) <= input(13);
output(2, 253) <= input(14);
output(2, 254) <= input(15);
output(2, 255) <= input(32);
output(3, 0) <= input(0);
output(3, 1) <= input(1);
output(3, 2) <= input(2);
output(3, 3) <= input(3);
output(3, 4) <= input(4);
output(3, 5) <= input(5);
output(3, 6) <= input(6);
output(3, 7) <= input(7);
output(3, 8) <= input(8);
output(3, 9) <= input(9);
output(3, 10) <= input(10);
output(3, 11) <= input(11);
output(3, 12) <= input(12);
output(3, 13) <= input(13);
output(3, 14) <= input(14);
output(3, 15) <= input(15);
output(3, 16) <= input(0);
output(3, 17) <= input(1);
output(3, 18) <= input(2);
output(3, 19) <= input(3);
output(3, 20) <= input(4);
output(3, 21) <= input(5);
output(3, 22) <= input(6);
output(3, 23) <= input(7);
output(3, 24) <= input(8);
output(3, 25) <= input(9);
output(3, 26) <= input(10);
output(3, 27) <= input(11);
output(3, 28) <= input(12);
output(3, 29) <= input(13);
output(3, 30) <= input(14);
output(3, 31) <= input(15);
output(3, 32) <= input(0);
output(3, 33) <= input(1);
output(3, 34) <= input(2);
output(3, 35) <= input(3);
output(3, 36) <= input(4);
output(3, 37) <= input(5);
output(3, 38) <= input(6);
output(3, 39) <= input(7);
output(3, 40) <= input(8);
output(3, 41) <= input(9);
output(3, 42) <= input(10);
output(3, 43) <= input(11);
output(3, 44) <= input(12);
output(3, 45) <= input(13);
output(3, 46) <= input(14);
output(3, 47) <= input(15);
output(3, 48) <= input(0);
output(3, 49) <= input(1);
output(3, 50) <= input(2);
output(3, 51) <= input(3);
output(3, 52) <= input(4);
output(3, 53) <= input(5);
output(3, 54) <= input(6);
output(3, 55) <= input(7);
output(3, 56) <= input(8);
output(3, 57) <= input(9);
output(3, 58) <= input(10);
output(3, 59) <= input(11);
output(3, 60) <= input(12);
output(3, 61) <= input(13);
output(3, 62) <= input(14);
output(3, 63) <= input(15);
output(3, 64) <= input(0);
output(3, 65) <= input(1);
output(3, 66) <= input(2);
output(3, 67) <= input(3);
output(3, 68) <= input(4);
output(3, 69) <= input(5);
output(3, 70) <= input(6);
output(3, 71) <= input(7);
output(3, 72) <= input(8);
output(3, 73) <= input(9);
output(3, 74) <= input(10);
output(3, 75) <= input(11);
output(3, 76) <= input(12);
output(3, 77) <= input(13);
output(3, 78) <= input(14);
output(3, 79) <= input(15);
output(3, 80) <= input(0);
output(3, 81) <= input(1);
output(3, 82) <= input(2);
output(3, 83) <= input(3);
output(3, 84) <= input(4);
output(3, 85) <= input(5);
output(3, 86) <= input(6);
output(3, 87) <= input(7);
output(3, 88) <= input(8);
output(3, 89) <= input(9);
output(3, 90) <= input(10);
output(3, 91) <= input(11);
output(3, 92) <= input(12);
output(3, 93) <= input(13);
output(3, 94) <= input(14);
output(3, 95) <= input(15);
output(3, 96) <= input(0);
output(3, 97) <= input(1);
output(3, 98) <= input(2);
output(3, 99) <= input(3);
output(3, 100) <= input(4);
output(3, 101) <= input(5);
output(3, 102) <= input(6);
output(3, 103) <= input(7);
output(3, 104) <= input(8);
output(3, 105) <= input(9);
output(3, 106) <= input(10);
output(3, 107) <= input(11);
output(3, 108) <= input(12);
output(3, 109) <= input(13);
output(3, 110) <= input(14);
output(3, 111) <= input(15);
output(3, 112) <= input(0);
output(3, 113) <= input(1);
output(3, 114) <= input(2);
output(3, 115) <= input(3);
output(3, 116) <= input(4);
output(3, 117) <= input(5);
output(3, 118) <= input(6);
output(3, 119) <= input(7);
output(3, 120) <= input(8);
output(3, 121) <= input(9);
output(3, 122) <= input(10);
output(3, 123) <= input(11);
output(3, 124) <= input(12);
output(3, 125) <= input(13);
output(3, 126) <= input(14);
output(3, 127) <= input(15);
output(3, 128) <= input(0);
output(3, 129) <= input(1);
output(3, 130) <= input(2);
output(3, 131) <= input(3);
output(3, 132) <= input(4);
output(3, 133) <= input(5);
output(3, 134) <= input(6);
output(3, 135) <= input(7);
output(3, 136) <= input(8);
output(3, 137) <= input(9);
output(3, 138) <= input(10);
output(3, 139) <= input(11);
output(3, 140) <= input(12);
output(3, 141) <= input(13);
output(3, 142) <= input(14);
output(3, 143) <= input(15);
output(3, 144) <= input(0);
output(3, 145) <= input(1);
output(3, 146) <= input(2);
output(3, 147) <= input(3);
output(3, 148) <= input(4);
output(3, 149) <= input(5);
output(3, 150) <= input(6);
output(3, 151) <= input(7);
output(3, 152) <= input(8);
output(3, 153) <= input(9);
output(3, 154) <= input(10);
output(3, 155) <= input(11);
output(3, 156) <= input(12);
output(3, 157) <= input(13);
output(3, 158) <= input(14);
output(3, 159) <= input(15);
output(3, 160) <= input(0);
output(3, 161) <= input(1);
output(3, 162) <= input(2);
output(3, 163) <= input(3);
output(3, 164) <= input(4);
output(3, 165) <= input(5);
output(3, 166) <= input(6);
output(3, 167) <= input(7);
output(3, 168) <= input(8);
output(3, 169) <= input(9);
output(3, 170) <= input(10);
output(3, 171) <= input(11);
output(3, 172) <= input(12);
output(3, 173) <= input(13);
output(3, 174) <= input(14);
output(3, 175) <= input(15);
output(3, 176) <= input(0);
output(3, 177) <= input(1);
output(3, 178) <= input(2);
output(3, 179) <= input(3);
output(3, 180) <= input(4);
output(3, 181) <= input(5);
output(3, 182) <= input(6);
output(3, 183) <= input(7);
output(3, 184) <= input(8);
output(3, 185) <= input(9);
output(3, 186) <= input(10);
output(3, 187) <= input(11);
output(3, 188) <= input(12);
output(3, 189) <= input(13);
output(3, 190) <= input(14);
output(3, 191) <= input(15);
output(3, 192) <= input(0);
output(3, 193) <= input(1);
output(3, 194) <= input(2);
output(3, 195) <= input(3);
output(3, 196) <= input(4);
output(3, 197) <= input(5);
output(3, 198) <= input(6);
output(3, 199) <= input(7);
output(3, 200) <= input(8);
output(3, 201) <= input(9);
output(3, 202) <= input(10);
output(3, 203) <= input(11);
output(3, 204) <= input(12);
output(3, 205) <= input(13);
output(3, 206) <= input(14);
output(3, 207) <= input(15);
output(3, 208) <= input(0);
output(3, 209) <= input(1);
output(3, 210) <= input(2);
output(3, 211) <= input(3);
output(3, 212) <= input(4);
output(3, 213) <= input(5);
output(3, 214) <= input(6);
output(3, 215) <= input(7);
output(3, 216) <= input(8);
output(3, 217) <= input(9);
output(3, 218) <= input(10);
output(3, 219) <= input(11);
output(3, 220) <= input(12);
output(3, 221) <= input(13);
output(3, 222) <= input(14);
output(3, 223) <= input(15);
output(3, 224) <= input(0);
output(3, 225) <= input(1);
output(3, 226) <= input(2);
output(3, 227) <= input(3);
output(3, 228) <= input(4);
output(3, 229) <= input(5);
output(3, 230) <= input(6);
output(3, 231) <= input(7);
output(3, 232) <= input(8);
output(3, 233) <= input(9);
output(3, 234) <= input(10);
output(3, 235) <= input(11);
output(3, 236) <= input(12);
output(3, 237) <= input(13);
output(3, 238) <= input(14);
output(3, 239) <= input(15);
output(3, 240) <= input(16);
output(3, 241) <= input(17);
output(3, 242) <= input(18);
output(3, 243) <= input(19);
output(3, 244) <= input(20);
output(3, 245) <= input(21);
output(3, 246) <= input(22);
output(3, 247) <= input(23);
output(3, 248) <= input(24);
output(3, 249) <= input(25);
output(3, 250) <= input(26);
output(3, 251) <= input(27);
output(3, 252) <= input(28);
output(3, 253) <= input(29);
output(3, 254) <= input(30);
output(3, 255) <= input(31);
output(4, 0) <= input(0);
output(4, 1) <= input(1);
output(4, 2) <= input(2);
output(4, 3) <= input(3);
output(4, 4) <= input(4);
output(4, 5) <= input(5);
output(4, 6) <= input(6);
output(4, 7) <= input(7);
output(4, 8) <= input(8);
output(4, 9) <= input(9);
output(4, 10) <= input(10);
output(4, 11) <= input(11);
output(4, 12) <= input(12);
output(4, 13) <= input(13);
output(4, 14) <= input(14);
output(4, 15) <= input(15);
output(4, 16) <= input(0);
output(4, 17) <= input(1);
output(4, 18) <= input(2);
output(4, 19) <= input(3);
output(4, 20) <= input(4);
output(4, 21) <= input(5);
output(4, 22) <= input(6);
output(4, 23) <= input(7);
output(4, 24) <= input(8);
output(4, 25) <= input(9);
output(4, 26) <= input(10);
output(4, 27) <= input(11);
output(4, 28) <= input(12);
output(4, 29) <= input(13);
output(4, 30) <= input(14);
output(4, 31) <= input(15);
output(4, 32) <= input(0);
output(4, 33) <= input(1);
output(4, 34) <= input(2);
output(4, 35) <= input(3);
output(4, 36) <= input(4);
output(4, 37) <= input(5);
output(4, 38) <= input(6);
output(4, 39) <= input(7);
output(4, 40) <= input(8);
output(4, 41) <= input(9);
output(4, 42) <= input(10);
output(4, 43) <= input(11);
output(4, 44) <= input(12);
output(4, 45) <= input(13);
output(4, 46) <= input(14);
output(4, 47) <= input(15);
output(4, 48) <= input(0);
output(4, 49) <= input(1);
output(4, 50) <= input(2);
output(4, 51) <= input(3);
output(4, 52) <= input(4);
output(4, 53) <= input(5);
output(4, 54) <= input(6);
output(4, 55) <= input(7);
output(4, 56) <= input(8);
output(4, 57) <= input(9);
output(4, 58) <= input(10);
output(4, 59) <= input(11);
output(4, 60) <= input(12);
output(4, 61) <= input(13);
output(4, 62) <= input(14);
output(4, 63) <= input(15);
output(4, 64) <= input(0);
output(4, 65) <= input(1);
output(4, 66) <= input(2);
output(4, 67) <= input(3);
output(4, 68) <= input(4);
output(4, 69) <= input(5);
output(4, 70) <= input(6);
output(4, 71) <= input(7);
output(4, 72) <= input(8);
output(4, 73) <= input(9);
output(4, 74) <= input(10);
output(4, 75) <= input(11);
output(4, 76) <= input(12);
output(4, 77) <= input(13);
output(4, 78) <= input(14);
output(4, 79) <= input(15);
output(4, 80) <= input(0);
output(4, 81) <= input(1);
output(4, 82) <= input(2);
output(4, 83) <= input(3);
output(4, 84) <= input(4);
output(4, 85) <= input(5);
output(4, 86) <= input(6);
output(4, 87) <= input(7);
output(4, 88) <= input(8);
output(4, 89) <= input(9);
output(4, 90) <= input(10);
output(4, 91) <= input(11);
output(4, 92) <= input(12);
output(4, 93) <= input(13);
output(4, 94) <= input(14);
output(4, 95) <= input(15);
output(4, 96) <= input(0);
output(4, 97) <= input(1);
output(4, 98) <= input(2);
output(4, 99) <= input(3);
output(4, 100) <= input(4);
output(4, 101) <= input(5);
output(4, 102) <= input(6);
output(4, 103) <= input(7);
output(4, 104) <= input(8);
output(4, 105) <= input(9);
output(4, 106) <= input(10);
output(4, 107) <= input(11);
output(4, 108) <= input(12);
output(4, 109) <= input(13);
output(4, 110) <= input(14);
output(4, 111) <= input(15);
output(4, 112) <= input(0);
output(4, 113) <= input(1);
output(4, 114) <= input(2);
output(4, 115) <= input(3);
output(4, 116) <= input(4);
output(4, 117) <= input(5);
output(4, 118) <= input(6);
output(4, 119) <= input(7);
output(4, 120) <= input(8);
output(4, 121) <= input(9);
output(4, 122) <= input(10);
output(4, 123) <= input(11);
output(4, 124) <= input(12);
output(4, 125) <= input(13);
output(4, 126) <= input(14);
output(4, 127) <= input(15);
output(4, 128) <= input(0);
output(4, 129) <= input(1);
output(4, 130) <= input(2);
output(4, 131) <= input(3);
output(4, 132) <= input(4);
output(4, 133) <= input(5);
output(4, 134) <= input(6);
output(4, 135) <= input(7);
output(4, 136) <= input(8);
output(4, 137) <= input(9);
output(4, 138) <= input(10);
output(4, 139) <= input(11);
output(4, 140) <= input(12);
output(4, 141) <= input(13);
output(4, 142) <= input(14);
output(4, 143) <= input(15);
output(4, 144) <= input(0);
output(4, 145) <= input(1);
output(4, 146) <= input(2);
output(4, 147) <= input(3);
output(4, 148) <= input(4);
output(4, 149) <= input(5);
output(4, 150) <= input(6);
output(4, 151) <= input(7);
output(4, 152) <= input(8);
output(4, 153) <= input(9);
output(4, 154) <= input(10);
output(4, 155) <= input(11);
output(4, 156) <= input(12);
output(4, 157) <= input(13);
output(4, 158) <= input(14);
output(4, 159) <= input(15);
output(4, 160) <= input(0);
output(4, 161) <= input(1);
output(4, 162) <= input(2);
output(4, 163) <= input(3);
output(4, 164) <= input(4);
output(4, 165) <= input(5);
output(4, 166) <= input(6);
output(4, 167) <= input(7);
output(4, 168) <= input(8);
output(4, 169) <= input(9);
output(4, 170) <= input(10);
output(4, 171) <= input(11);
output(4, 172) <= input(12);
output(4, 173) <= input(13);
output(4, 174) <= input(14);
output(4, 175) <= input(15);
output(4, 176) <= input(0);
output(4, 177) <= input(1);
output(4, 178) <= input(2);
output(4, 179) <= input(3);
output(4, 180) <= input(4);
output(4, 181) <= input(5);
output(4, 182) <= input(6);
output(4, 183) <= input(7);
output(4, 184) <= input(8);
output(4, 185) <= input(9);
output(4, 186) <= input(10);
output(4, 187) <= input(11);
output(4, 188) <= input(12);
output(4, 189) <= input(13);
output(4, 190) <= input(14);
output(4, 191) <= input(15);
output(4, 192) <= input(0);
output(4, 193) <= input(1);
output(4, 194) <= input(2);
output(4, 195) <= input(3);
output(4, 196) <= input(4);
output(4, 197) <= input(5);
output(4, 198) <= input(6);
output(4, 199) <= input(7);
output(4, 200) <= input(8);
output(4, 201) <= input(9);
output(4, 202) <= input(10);
output(4, 203) <= input(11);
output(4, 204) <= input(12);
output(4, 205) <= input(13);
output(4, 206) <= input(14);
output(4, 207) <= input(15);
output(4, 208) <= input(0);
output(4, 209) <= input(1);
output(4, 210) <= input(2);
output(4, 211) <= input(3);
output(4, 212) <= input(4);
output(4, 213) <= input(5);
output(4, 214) <= input(6);
output(4, 215) <= input(7);
output(4, 216) <= input(8);
output(4, 217) <= input(9);
output(4, 218) <= input(10);
output(4, 219) <= input(11);
output(4, 220) <= input(12);
output(4, 221) <= input(13);
output(4, 222) <= input(14);
output(4, 223) <= input(15);
output(4, 224) <= input(0);
output(4, 225) <= input(1);
output(4, 226) <= input(2);
output(4, 227) <= input(3);
output(4, 228) <= input(4);
output(4, 229) <= input(5);
output(4, 230) <= input(6);
output(4, 231) <= input(7);
output(4, 232) <= input(8);
output(4, 233) <= input(9);
output(4, 234) <= input(10);
output(4, 235) <= input(11);
output(4, 236) <= input(12);
output(4, 237) <= input(13);
output(4, 238) <= input(14);
output(4, 239) <= input(15);
output(4, 240) <= input(0);
output(4, 241) <= input(1);
output(4, 242) <= input(2);
output(4, 243) <= input(3);
output(4, 244) <= input(4);
output(4, 245) <= input(5);
output(4, 246) <= input(6);
output(4, 247) <= input(7);
output(4, 248) <= input(8);
output(4, 249) <= input(9);
output(4, 250) <= input(10);
output(4, 251) <= input(11);
output(4, 252) <= input(12);
output(4, 253) <= input(13);
output(4, 254) <= input(14);
output(4, 255) <= input(15);
output(5, 0) <= input(35);
output(5, 1) <= input(16);
output(5, 2) <= input(17);
output(5, 3) <= input(18);
output(5, 4) <= input(19);
output(5, 5) <= input(20);
output(5, 6) <= input(21);
output(5, 7) <= input(22);
output(5, 8) <= input(23);
output(5, 9) <= input(24);
output(5, 10) <= input(25);
output(5, 11) <= input(26);
output(5, 12) <= input(27);
output(5, 13) <= input(28);
output(5, 14) <= input(29);
output(5, 15) <= input(30);
output(5, 16) <= input(35);
output(5, 17) <= input(16);
output(5, 18) <= input(17);
output(5, 19) <= input(18);
output(5, 20) <= input(19);
output(5, 21) <= input(20);
output(5, 22) <= input(21);
output(5, 23) <= input(22);
output(5, 24) <= input(23);
output(5, 25) <= input(24);
output(5, 26) <= input(25);
output(5, 27) <= input(26);
output(5, 28) <= input(27);
output(5, 29) <= input(28);
output(5, 30) <= input(29);
output(5, 31) <= input(30);
output(5, 32) <= input(35);
output(5, 33) <= input(16);
output(5, 34) <= input(17);
output(5, 35) <= input(18);
output(5, 36) <= input(19);
output(5, 37) <= input(20);
output(5, 38) <= input(21);
output(5, 39) <= input(22);
output(5, 40) <= input(23);
output(5, 41) <= input(24);
output(5, 42) <= input(25);
output(5, 43) <= input(26);
output(5, 44) <= input(27);
output(5, 45) <= input(28);
output(5, 46) <= input(29);
output(5, 47) <= input(30);
output(5, 48) <= input(35);
output(5, 49) <= input(16);
output(5, 50) <= input(17);
output(5, 51) <= input(18);
output(5, 52) <= input(19);
output(5, 53) <= input(20);
output(5, 54) <= input(21);
output(5, 55) <= input(22);
output(5, 56) <= input(23);
output(5, 57) <= input(24);
output(5, 58) <= input(25);
output(5, 59) <= input(26);
output(5, 60) <= input(27);
output(5, 61) <= input(28);
output(5, 62) <= input(29);
output(5, 63) <= input(30);
output(5, 64) <= input(35);
output(5, 65) <= input(16);
output(5, 66) <= input(17);
output(5, 67) <= input(18);
output(5, 68) <= input(19);
output(5, 69) <= input(20);
output(5, 70) <= input(21);
output(5, 71) <= input(22);
output(5, 72) <= input(23);
output(5, 73) <= input(24);
output(5, 74) <= input(25);
output(5, 75) <= input(26);
output(5, 76) <= input(27);
output(5, 77) <= input(28);
output(5, 78) <= input(29);
output(5, 79) <= input(30);
output(5, 80) <= input(35);
output(5, 81) <= input(16);
output(5, 82) <= input(17);
output(5, 83) <= input(18);
output(5, 84) <= input(19);
output(5, 85) <= input(20);
output(5, 86) <= input(21);
output(5, 87) <= input(22);
output(5, 88) <= input(23);
output(5, 89) <= input(24);
output(5, 90) <= input(25);
output(5, 91) <= input(26);
output(5, 92) <= input(27);
output(5, 93) <= input(28);
output(5, 94) <= input(29);
output(5, 95) <= input(30);
output(5, 96) <= input(35);
output(5, 97) <= input(16);
output(5, 98) <= input(17);
output(5, 99) <= input(18);
output(5, 100) <= input(19);
output(5, 101) <= input(20);
output(5, 102) <= input(21);
output(5, 103) <= input(22);
output(5, 104) <= input(23);
output(5, 105) <= input(24);
output(5, 106) <= input(25);
output(5, 107) <= input(26);
output(5, 108) <= input(27);
output(5, 109) <= input(28);
output(5, 110) <= input(29);
output(5, 111) <= input(30);
output(5, 112) <= input(35);
output(5, 113) <= input(16);
output(5, 114) <= input(17);
output(5, 115) <= input(18);
output(5, 116) <= input(19);
output(5, 117) <= input(20);
output(5, 118) <= input(21);
output(5, 119) <= input(22);
output(5, 120) <= input(23);
output(5, 121) <= input(24);
output(5, 122) <= input(25);
output(5, 123) <= input(26);
output(5, 124) <= input(27);
output(5, 125) <= input(28);
output(5, 126) <= input(29);
output(5, 127) <= input(30);
output(5, 128) <= input(35);
output(5, 129) <= input(16);
output(5, 130) <= input(17);
output(5, 131) <= input(18);
output(5, 132) <= input(19);
output(5, 133) <= input(20);
output(5, 134) <= input(21);
output(5, 135) <= input(22);
output(5, 136) <= input(23);
output(5, 137) <= input(24);
output(5, 138) <= input(25);
output(5, 139) <= input(26);
output(5, 140) <= input(27);
output(5, 141) <= input(28);
output(5, 142) <= input(29);
output(5, 143) <= input(30);
output(5, 144) <= input(35);
output(5, 145) <= input(16);
output(5, 146) <= input(17);
output(5, 147) <= input(18);
output(5, 148) <= input(19);
output(5, 149) <= input(20);
output(5, 150) <= input(21);
output(5, 151) <= input(22);
output(5, 152) <= input(23);
output(5, 153) <= input(24);
output(5, 154) <= input(25);
output(5, 155) <= input(26);
output(5, 156) <= input(27);
output(5, 157) <= input(28);
output(5, 158) <= input(29);
output(5, 159) <= input(30);
output(5, 160) <= input(35);
output(5, 161) <= input(16);
output(5, 162) <= input(17);
output(5, 163) <= input(18);
output(5, 164) <= input(19);
output(5, 165) <= input(20);
output(5, 166) <= input(21);
output(5, 167) <= input(22);
output(5, 168) <= input(23);
output(5, 169) <= input(24);
output(5, 170) <= input(25);
output(5, 171) <= input(26);
output(5, 172) <= input(27);
output(5, 173) <= input(28);
output(5, 174) <= input(29);
output(5, 175) <= input(30);
output(5, 176) <= input(35);
output(5, 177) <= input(16);
output(5, 178) <= input(17);
output(5, 179) <= input(18);
output(5, 180) <= input(19);
output(5, 181) <= input(20);
output(5, 182) <= input(21);
output(5, 183) <= input(22);
output(5, 184) <= input(23);
output(5, 185) <= input(24);
output(5, 186) <= input(25);
output(5, 187) <= input(26);
output(5, 188) <= input(27);
output(5, 189) <= input(28);
output(5, 190) <= input(29);
output(5, 191) <= input(30);
output(5, 192) <= input(35);
output(5, 193) <= input(16);
output(5, 194) <= input(17);
output(5, 195) <= input(18);
output(5, 196) <= input(19);
output(5, 197) <= input(20);
output(5, 198) <= input(21);
output(5, 199) <= input(22);
output(5, 200) <= input(23);
output(5, 201) <= input(24);
output(5, 202) <= input(25);
output(5, 203) <= input(26);
output(5, 204) <= input(27);
output(5, 205) <= input(28);
output(5, 206) <= input(29);
output(5, 207) <= input(30);
output(5, 208) <= input(35);
output(5, 209) <= input(16);
output(5, 210) <= input(17);
output(5, 211) <= input(18);
output(5, 212) <= input(19);
output(5, 213) <= input(20);
output(5, 214) <= input(21);
output(5, 215) <= input(22);
output(5, 216) <= input(23);
output(5, 217) <= input(24);
output(5, 218) <= input(25);
output(5, 219) <= input(26);
output(5, 220) <= input(27);
output(5, 221) <= input(28);
output(5, 222) <= input(29);
output(5, 223) <= input(30);
output(5, 224) <= input(35);
output(5, 225) <= input(16);
output(5, 226) <= input(17);
output(5, 227) <= input(18);
output(5, 228) <= input(19);
output(5, 229) <= input(20);
output(5, 230) <= input(21);
output(5, 231) <= input(22);
output(5, 232) <= input(23);
output(5, 233) <= input(24);
output(5, 234) <= input(25);
output(5, 235) <= input(26);
output(5, 236) <= input(27);
output(5, 237) <= input(28);
output(5, 238) <= input(29);
output(5, 239) <= input(30);
output(5, 240) <= input(35);
output(5, 241) <= input(16);
output(5, 242) <= input(17);
output(5, 243) <= input(18);
output(5, 244) <= input(19);
output(5, 245) <= input(20);
output(5, 246) <= input(21);
output(5, 247) <= input(22);
output(5, 248) <= input(23);
output(5, 249) <= input(24);
output(5, 250) <= input(25);
output(5, 251) <= input(26);
output(5, 252) <= input(27);
output(5, 253) <= input(28);
output(5, 254) <= input(29);
output(5, 255) <= input(30);
output(6, 0) <= input(36);
output(6, 1) <= input(16);
output(6, 2) <= input(17);
output(6, 3) <= input(18);
output(6, 4) <= input(19);
output(6, 5) <= input(20);
output(6, 6) <= input(21);
output(6, 7) <= input(22);
output(6, 8) <= input(23);
output(6, 9) <= input(24);
output(6, 10) <= input(25);
output(6, 11) <= input(26);
output(6, 12) <= input(27);
output(6, 13) <= input(28);
output(6, 14) <= input(29);
output(6, 15) <= input(30);
output(6, 16) <= input(36);
output(6, 17) <= input(16);
output(6, 18) <= input(17);
output(6, 19) <= input(18);
output(6, 20) <= input(19);
output(6, 21) <= input(20);
output(6, 22) <= input(21);
output(6, 23) <= input(22);
output(6, 24) <= input(23);
output(6, 25) <= input(24);
output(6, 26) <= input(25);
output(6, 27) <= input(26);
output(6, 28) <= input(27);
output(6, 29) <= input(28);
output(6, 30) <= input(29);
output(6, 31) <= input(30);
output(6, 32) <= input(36);
output(6, 33) <= input(16);
output(6, 34) <= input(17);
output(6, 35) <= input(18);
output(6, 36) <= input(19);
output(6, 37) <= input(20);
output(6, 38) <= input(21);
output(6, 39) <= input(22);
output(6, 40) <= input(23);
output(6, 41) <= input(24);
output(6, 42) <= input(25);
output(6, 43) <= input(26);
output(6, 44) <= input(27);
output(6, 45) <= input(28);
output(6, 46) <= input(29);
output(6, 47) <= input(30);
output(6, 48) <= input(36);
output(6, 49) <= input(16);
output(6, 50) <= input(17);
output(6, 51) <= input(18);
output(6, 52) <= input(19);
output(6, 53) <= input(20);
output(6, 54) <= input(21);
output(6, 55) <= input(22);
output(6, 56) <= input(23);
output(6, 57) <= input(24);
output(6, 58) <= input(25);
output(6, 59) <= input(26);
output(6, 60) <= input(27);
output(6, 61) <= input(28);
output(6, 62) <= input(29);
output(6, 63) <= input(30);
output(6, 64) <= input(36);
output(6, 65) <= input(16);
output(6, 66) <= input(17);
output(6, 67) <= input(18);
output(6, 68) <= input(19);
output(6, 69) <= input(20);
output(6, 70) <= input(21);
output(6, 71) <= input(22);
output(6, 72) <= input(23);
output(6, 73) <= input(24);
output(6, 74) <= input(25);
output(6, 75) <= input(26);
output(6, 76) <= input(27);
output(6, 77) <= input(28);
output(6, 78) <= input(29);
output(6, 79) <= input(30);
output(6, 80) <= input(36);
output(6, 81) <= input(16);
output(6, 82) <= input(17);
output(6, 83) <= input(18);
output(6, 84) <= input(19);
output(6, 85) <= input(20);
output(6, 86) <= input(21);
output(6, 87) <= input(22);
output(6, 88) <= input(23);
output(6, 89) <= input(24);
output(6, 90) <= input(25);
output(6, 91) <= input(26);
output(6, 92) <= input(27);
output(6, 93) <= input(28);
output(6, 94) <= input(29);
output(6, 95) <= input(30);
output(6, 96) <= input(36);
output(6, 97) <= input(16);
output(6, 98) <= input(17);
output(6, 99) <= input(18);
output(6, 100) <= input(19);
output(6, 101) <= input(20);
output(6, 102) <= input(21);
output(6, 103) <= input(22);
output(6, 104) <= input(23);
output(6, 105) <= input(24);
output(6, 106) <= input(25);
output(6, 107) <= input(26);
output(6, 108) <= input(27);
output(6, 109) <= input(28);
output(6, 110) <= input(29);
output(6, 111) <= input(30);
output(6, 112) <= input(36);
output(6, 113) <= input(16);
output(6, 114) <= input(17);
output(6, 115) <= input(18);
output(6, 116) <= input(19);
output(6, 117) <= input(20);
output(6, 118) <= input(21);
output(6, 119) <= input(22);
output(6, 120) <= input(23);
output(6, 121) <= input(24);
output(6, 122) <= input(25);
output(6, 123) <= input(26);
output(6, 124) <= input(27);
output(6, 125) <= input(28);
output(6, 126) <= input(29);
output(6, 127) <= input(30);
output(6, 128) <= input(37);
output(6, 129) <= input(0);
output(6, 130) <= input(1);
output(6, 131) <= input(2);
output(6, 132) <= input(3);
output(6, 133) <= input(4);
output(6, 134) <= input(5);
output(6, 135) <= input(6);
output(6, 136) <= input(7);
output(6, 137) <= input(8);
output(6, 138) <= input(9);
output(6, 139) <= input(10);
output(6, 140) <= input(11);
output(6, 141) <= input(12);
output(6, 142) <= input(13);
output(6, 143) <= input(14);
output(6, 144) <= input(37);
output(6, 145) <= input(0);
output(6, 146) <= input(1);
output(6, 147) <= input(2);
output(6, 148) <= input(3);
output(6, 149) <= input(4);
output(6, 150) <= input(5);
output(6, 151) <= input(6);
output(6, 152) <= input(7);
output(6, 153) <= input(8);
output(6, 154) <= input(9);
output(6, 155) <= input(10);
output(6, 156) <= input(11);
output(6, 157) <= input(12);
output(6, 158) <= input(13);
output(6, 159) <= input(14);
output(6, 160) <= input(37);
output(6, 161) <= input(0);
output(6, 162) <= input(1);
output(6, 163) <= input(2);
output(6, 164) <= input(3);
output(6, 165) <= input(4);
output(6, 166) <= input(5);
output(6, 167) <= input(6);
output(6, 168) <= input(7);
output(6, 169) <= input(8);
output(6, 170) <= input(9);
output(6, 171) <= input(10);
output(6, 172) <= input(11);
output(6, 173) <= input(12);
output(6, 174) <= input(13);
output(6, 175) <= input(14);
output(6, 176) <= input(37);
output(6, 177) <= input(0);
output(6, 178) <= input(1);
output(6, 179) <= input(2);
output(6, 180) <= input(3);
output(6, 181) <= input(4);
output(6, 182) <= input(5);
output(6, 183) <= input(6);
output(6, 184) <= input(7);
output(6, 185) <= input(8);
output(6, 186) <= input(9);
output(6, 187) <= input(10);
output(6, 188) <= input(11);
output(6, 189) <= input(12);
output(6, 190) <= input(13);
output(6, 191) <= input(14);
output(6, 192) <= input(37);
output(6, 193) <= input(0);
output(6, 194) <= input(1);
output(6, 195) <= input(2);
output(6, 196) <= input(3);
output(6, 197) <= input(4);
output(6, 198) <= input(5);
output(6, 199) <= input(6);
output(6, 200) <= input(7);
output(6, 201) <= input(8);
output(6, 202) <= input(9);
output(6, 203) <= input(10);
output(6, 204) <= input(11);
output(6, 205) <= input(12);
output(6, 206) <= input(13);
output(6, 207) <= input(14);
output(6, 208) <= input(37);
output(6, 209) <= input(0);
output(6, 210) <= input(1);
output(6, 211) <= input(2);
output(6, 212) <= input(3);
output(6, 213) <= input(4);
output(6, 214) <= input(5);
output(6, 215) <= input(6);
output(6, 216) <= input(7);
output(6, 217) <= input(8);
output(6, 218) <= input(9);
output(6, 219) <= input(10);
output(6, 220) <= input(11);
output(6, 221) <= input(12);
output(6, 222) <= input(13);
output(6, 223) <= input(14);
output(6, 224) <= input(37);
output(6, 225) <= input(0);
output(6, 226) <= input(1);
output(6, 227) <= input(2);
output(6, 228) <= input(3);
output(6, 229) <= input(4);
output(6, 230) <= input(5);
output(6, 231) <= input(6);
output(6, 232) <= input(7);
output(6, 233) <= input(8);
output(6, 234) <= input(9);
output(6, 235) <= input(10);
output(6, 236) <= input(11);
output(6, 237) <= input(12);
output(6, 238) <= input(13);
output(6, 239) <= input(14);
output(6, 240) <= input(37);
output(6, 241) <= input(0);
output(6, 242) <= input(1);
output(6, 243) <= input(2);
output(6, 244) <= input(3);
output(6, 245) <= input(4);
output(6, 246) <= input(5);
output(6, 247) <= input(6);
output(6, 248) <= input(7);
output(6, 249) <= input(8);
output(6, 250) <= input(9);
output(6, 251) <= input(10);
output(6, 252) <= input(11);
output(6, 253) <= input(12);
output(6, 254) <= input(13);
output(6, 255) <= input(14);
output(7, 0) <= input(38);
output(7, 1) <= input(16);
output(7, 2) <= input(17);
output(7, 3) <= input(18);
output(7, 4) <= input(19);
output(7, 5) <= input(20);
output(7, 6) <= input(21);
output(7, 7) <= input(22);
output(7, 8) <= input(23);
output(7, 9) <= input(24);
output(7, 10) <= input(25);
output(7, 11) <= input(26);
output(7, 12) <= input(27);
output(7, 13) <= input(28);
output(7, 14) <= input(29);
output(7, 15) <= input(30);
output(7, 16) <= input(38);
output(7, 17) <= input(16);
output(7, 18) <= input(17);
output(7, 19) <= input(18);
output(7, 20) <= input(19);
output(7, 21) <= input(20);
output(7, 22) <= input(21);
output(7, 23) <= input(22);
output(7, 24) <= input(23);
output(7, 25) <= input(24);
output(7, 26) <= input(25);
output(7, 27) <= input(26);
output(7, 28) <= input(27);
output(7, 29) <= input(28);
output(7, 30) <= input(29);
output(7, 31) <= input(30);
output(7, 32) <= input(38);
output(7, 33) <= input(16);
output(7, 34) <= input(17);
output(7, 35) <= input(18);
output(7, 36) <= input(19);
output(7, 37) <= input(20);
output(7, 38) <= input(21);
output(7, 39) <= input(22);
output(7, 40) <= input(23);
output(7, 41) <= input(24);
output(7, 42) <= input(25);
output(7, 43) <= input(26);
output(7, 44) <= input(27);
output(7, 45) <= input(28);
output(7, 46) <= input(29);
output(7, 47) <= input(30);
output(7, 48) <= input(38);
output(7, 49) <= input(16);
output(7, 50) <= input(17);
output(7, 51) <= input(18);
output(7, 52) <= input(19);
output(7, 53) <= input(20);
output(7, 54) <= input(21);
output(7, 55) <= input(22);
output(7, 56) <= input(23);
output(7, 57) <= input(24);
output(7, 58) <= input(25);
output(7, 59) <= input(26);
output(7, 60) <= input(27);
output(7, 61) <= input(28);
output(7, 62) <= input(29);
output(7, 63) <= input(30);
output(7, 64) <= input(38);
output(7, 65) <= input(16);
output(7, 66) <= input(17);
output(7, 67) <= input(18);
output(7, 68) <= input(19);
output(7, 69) <= input(20);
output(7, 70) <= input(21);
output(7, 71) <= input(22);
output(7, 72) <= input(23);
output(7, 73) <= input(24);
output(7, 74) <= input(25);
output(7, 75) <= input(26);
output(7, 76) <= input(27);
output(7, 77) <= input(28);
output(7, 78) <= input(29);
output(7, 79) <= input(30);
output(7, 80) <= input(39);
output(7, 81) <= input(0);
output(7, 82) <= input(1);
output(7, 83) <= input(2);
output(7, 84) <= input(3);
output(7, 85) <= input(4);
output(7, 86) <= input(5);
output(7, 87) <= input(6);
output(7, 88) <= input(7);
output(7, 89) <= input(8);
output(7, 90) <= input(9);
output(7, 91) <= input(10);
output(7, 92) <= input(11);
output(7, 93) <= input(12);
output(7, 94) <= input(13);
output(7, 95) <= input(14);
output(7, 96) <= input(39);
output(7, 97) <= input(0);
output(7, 98) <= input(1);
output(7, 99) <= input(2);
output(7, 100) <= input(3);
output(7, 101) <= input(4);
output(7, 102) <= input(5);
output(7, 103) <= input(6);
output(7, 104) <= input(7);
output(7, 105) <= input(8);
output(7, 106) <= input(9);
output(7, 107) <= input(10);
output(7, 108) <= input(11);
output(7, 109) <= input(12);
output(7, 110) <= input(13);
output(7, 111) <= input(14);
output(7, 112) <= input(39);
output(7, 113) <= input(0);
output(7, 114) <= input(1);
output(7, 115) <= input(2);
output(7, 116) <= input(3);
output(7, 117) <= input(4);
output(7, 118) <= input(5);
output(7, 119) <= input(6);
output(7, 120) <= input(7);
output(7, 121) <= input(8);
output(7, 122) <= input(9);
output(7, 123) <= input(10);
output(7, 124) <= input(11);
output(7, 125) <= input(12);
output(7, 126) <= input(13);
output(7, 127) <= input(14);
output(7, 128) <= input(39);
output(7, 129) <= input(0);
output(7, 130) <= input(1);
output(7, 131) <= input(2);
output(7, 132) <= input(3);
output(7, 133) <= input(4);
output(7, 134) <= input(5);
output(7, 135) <= input(6);
output(7, 136) <= input(7);
output(7, 137) <= input(8);
output(7, 138) <= input(9);
output(7, 139) <= input(10);
output(7, 140) <= input(11);
output(7, 141) <= input(12);
output(7, 142) <= input(13);
output(7, 143) <= input(14);
output(7, 144) <= input(39);
output(7, 145) <= input(0);
output(7, 146) <= input(1);
output(7, 147) <= input(2);
output(7, 148) <= input(3);
output(7, 149) <= input(4);
output(7, 150) <= input(5);
output(7, 151) <= input(6);
output(7, 152) <= input(7);
output(7, 153) <= input(8);
output(7, 154) <= input(9);
output(7, 155) <= input(10);
output(7, 156) <= input(11);
output(7, 157) <= input(12);
output(7, 158) <= input(13);
output(7, 159) <= input(14);
output(7, 160) <= input(40);
output(7, 161) <= input(38);
output(7, 162) <= input(16);
output(7, 163) <= input(17);
output(7, 164) <= input(18);
output(7, 165) <= input(19);
output(7, 166) <= input(20);
output(7, 167) <= input(21);
output(7, 168) <= input(22);
output(7, 169) <= input(23);
output(7, 170) <= input(24);
output(7, 171) <= input(25);
output(7, 172) <= input(26);
output(7, 173) <= input(27);
output(7, 174) <= input(28);
output(7, 175) <= input(29);
output(7, 176) <= input(40);
output(7, 177) <= input(38);
output(7, 178) <= input(16);
output(7, 179) <= input(17);
output(7, 180) <= input(18);
output(7, 181) <= input(19);
output(7, 182) <= input(20);
output(7, 183) <= input(21);
output(7, 184) <= input(22);
output(7, 185) <= input(23);
output(7, 186) <= input(24);
output(7, 187) <= input(25);
output(7, 188) <= input(26);
output(7, 189) <= input(27);
output(7, 190) <= input(28);
output(7, 191) <= input(29);
output(7, 192) <= input(40);
output(7, 193) <= input(38);
output(7, 194) <= input(16);
output(7, 195) <= input(17);
output(7, 196) <= input(18);
output(7, 197) <= input(19);
output(7, 198) <= input(20);
output(7, 199) <= input(21);
output(7, 200) <= input(22);
output(7, 201) <= input(23);
output(7, 202) <= input(24);
output(7, 203) <= input(25);
output(7, 204) <= input(26);
output(7, 205) <= input(27);
output(7, 206) <= input(28);
output(7, 207) <= input(29);
output(7, 208) <= input(40);
output(7, 209) <= input(38);
output(7, 210) <= input(16);
output(7, 211) <= input(17);
output(7, 212) <= input(18);
output(7, 213) <= input(19);
output(7, 214) <= input(20);
output(7, 215) <= input(21);
output(7, 216) <= input(22);
output(7, 217) <= input(23);
output(7, 218) <= input(24);
output(7, 219) <= input(25);
output(7, 220) <= input(26);
output(7, 221) <= input(27);
output(7, 222) <= input(28);
output(7, 223) <= input(29);
output(7, 224) <= input(40);
output(7, 225) <= input(38);
output(7, 226) <= input(16);
output(7, 227) <= input(17);
output(7, 228) <= input(18);
output(7, 229) <= input(19);
output(7, 230) <= input(20);
output(7, 231) <= input(21);
output(7, 232) <= input(22);
output(7, 233) <= input(23);
output(7, 234) <= input(24);
output(7, 235) <= input(25);
output(7, 236) <= input(26);
output(7, 237) <= input(27);
output(7, 238) <= input(28);
output(7, 239) <= input(29);
output(7, 240) <= input(40);
output(7, 241) <= input(38);
output(7, 242) <= input(16);
output(7, 243) <= input(17);
output(7, 244) <= input(18);
output(7, 245) <= input(19);
output(7, 246) <= input(20);
output(7, 247) <= input(21);
output(7, 248) <= input(22);
output(7, 249) <= input(23);
output(7, 250) <= input(24);
output(7, 251) <= input(25);
output(7, 252) <= input(26);
output(7, 253) <= input(27);
output(7, 254) <= input(28);
output(7, 255) <= input(29);
when "0011" =>
output(0, 0) <= input(0);
output(0, 1) <= input(1);
output(0, 2) <= input(2);
output(0, 3) <= input(3);
output(0, 4) <= input(4);
output(0, 5) <= input(5);
output(0, 6) <= input(6);
output(0, 7) <= input(7);
output(0, 8) <= input(8);
output(0, 9) <= input(9);
output(0, 10) <= input(10);
output(0, 11) <= input(11);
output(0, 12) <= input(12);
output(0, 13) <= input(13);
output(0, 14) <= input(14);
output(0, 15) <= input(15);
output(0, 16) <= input(0);
output(0, 17) <= input(1);
output(0, 18) <= input(2);
output(0, 19) <= input(3);
output(0, 20) <= input(4);
output(0, 21) <= input(5);
output(0, 22) <= input(6);
output(0, 23) <= input(7);
output(0, 24) <= input(8);
output(0, 25) <= input(9);
output(0, 26) <= input(10);
output(0, 27) <= input(11);
output(0, 28) <= input(12);
output(0, 29) <= input(13);
output(0, 30) <= input(14);
output(0, 31) <= input(15);
output(0, 32) <= input(0);
output(0, 33) <= input(1);
output(0, 34) <= input(2);
output(0, 35) <= input(3);
output(0, 36) <= input(4);
output(0, 37) <= input(5);
output(0, 38) <= input(6);
output(0, 39) <= input(7);
output(0, 40) <= input(8);
output(0, 41) <= input(9);
output(0, 42) <= input(10);
output(0, 43) <= input(11);
output(0, 44) <= input(12);
output(0, 45) <= input(13);
output(0, 46) <= input(14);
output(0, 47) <= input(15);
output(0, 48) <= input(0);
output(0, 49) <= input(1);
output(0, 50) <= input(2);
output(0, 51) <= input(3);
output(0, 52) <= input(4);
output(0, 53) <= input(5);
output(0, 54) <= input(6);
output(0, 55) <= input(7);
output(0, 56) <= input(8);
output(0, 57) <= input(9);
output(0, 58) <= input(10);
output(0, 59) <= input(11);
output(0, 60) <= input(12);
output(0, 61) <= input(13);
output(0, 62) <= input(14);
output(0, 63) <= input(15);
output(0, 64) <= input(16);
output(0, 65) <= input(17);
output(0, 66) <= input(18);
output(0, 67) <= input(19);
output(0, 68) <= input(20);
output(0, 69) <= input(21);
output(0, 70) <= input(22);
output(0, 71) <= input(23);
output(0, 72) <= input(24);
output(0, 73) <= input(25);
output(0, 74) <= input(26);
output(0, 75) <= input(27);
output(0, 76) <= input(28);
output(0, 77) <= input(29);
output(0, 78) <= input(30);
output(0, 79) <= input(31);
output(0, 80) <= input(16);
output(0, 81) <= input(17);
output(0, 82) <= input(18);
output(0, 83) <= input(19);
output(0, 84) <= input(20);
output(0, 85) <= input(21);
output(0, 86) <= input(22);
output(0, 87) <= input(23);
output(0, 88) <= input(24);
output(0, 89) <= input(25);
output(0, 90) <= input(26);
output(0, 91) <= input(27);
output(0, 92) <= input(28);
output(0, 93) <= input(29);
output(0, 94) <= input(30);
output(0, 95) <= input(31);
output(0, 96) <= input(16);
output(0, 97) <= input(17);
output(0, 98) <= input(18);
output(0, 99) <= input(19);
output(0, 100) <= input(20);
output(0, 101) <= input(21);
output(0, 102) <= input(22);
output(0, 103) <= input(23);
output(0, 104) <= input(24);
output(0, 105) <= input(25);
output(0, 106) <= input(26);
output(0, 107) <= input(27);
output(0, 108) <= input(28);
output(0, 109) <= input(29);
output(0, 110) <= input(30);
output(0, 111) <= input(31);
output(0, 112) <= input(16);
output(0, 113) <= input(17);
output(0, 114) <= input(18);
output(0, 115) <= input(19);
output(0, 116) <= input(20);
output(0, 117) <= input(21);
output(0, 118) <= input(22);
output(0, 119) <= input(23);
output(0, 120) <= input(24);
output(0, 121) <= input(25);
output(0, 122) <= input(26);
output(0, 123) <= input(27);
output(0, 124) <= input(28);
output(0, 125) <= input(29);
output(0, 126) <= input(30);
output(0, 127) <= input(31);
output(0, 128) <= input(32);
output(0, 129) <= input(0);
output(0, 130) <= input(1);
output(0, 131) <= input(2);
output(0, 132) <= input(3);
output(0, 133) <= input(4);
output(0, 134) <= input(5);
output(0, 135) <= input(6);
output(0, 136) <= input(7);
output(0, 137) <= input(8);
output(0, 138) <= input(9);
output(0, 139) <= input(10);
output(0, 140) <= input(11);
output(0, 141) <= input(12);
output(0, 142) <= input(13);
output(0, 143) <= input(14);
output(0, 144) <= input(32);
output(0, 145) <= input(0);
output(0, 146) <= input(1);
output(0, 147) <= input(2);
output(0, 148) <= input(3);
output(0, 149) <= input(4);
output(0, 150) <= input(5);
output(0, 151) <= input(6);
output(0, 152) <= input(7);
output(0, 153) <= input(8);
output(0, 154) <= input(9);
output(0, 155) <= input(10);
output(0, 156) <= input(11);
output(0, 157) <= input(12);
output(0, 158) <= input(13);
output(0, 159) <= input(14);
output(0, 160) <= input(32);
output(0, 161) <= input(0);
output(0, 162) <= input(1);
output(0, 163) <= input(2);
output(0, 164) <= input(3);
output(0, 165) <= input(4);
output(0, 166) <= input(5);
output(0, 167) <= input(6);
output(0, 168) <= input(7);
output(0, 169) <= input(8);
output(0, 170) <= input(9);
output(0, 171) <= input(10);
output(0, 172) <= input(11);
output(0, 173) <= input(12);
output(0, 174) <= input(13);
output(0, 175) <= input(14);
output(0, 176) <= input(32);
output(0, 177) <= input(0);
output(0, 178) <= input(1);
output(0, 179) <= input(2);
output(0, 180) <= input(3);
output(0, 181) <= input(4);
output(0, 182) <= input(5);
output(0, 183) <= input(6);
output(0, 184) <= input(7);
output(0, 185) <= input(8);
output(0, 186) <= input(9);
output(0, 187) <= input(10);
output(0, 188) <= input(11);
output(0, 189) <= input(12);
output(0, 190) <= input(13);
output(0, 191) <= input(14);
output(0, 192) <= input(33);
output(0, 193) <= input(16);
output(0, 194) <= input(17);
output(0, 195) <= input(18);
output(0, 196) <= input(19);
output(0, 197) <= input(20);
output(0, 198) <= input(21);
output(0, 199) <= input(22);
output(0, 200) <= input(23);
output(0, 201) <= input(24);
output(0, 202) <= input(25);
output(0, 203) <= input(26);
output(0, 204) <= input(27);
output(0, 205) <= input(28);
output(0, 206) <= input(29);
output(0, 207) <= input(30);
output(0, 208) <= input(33);
output(0, 209) <= input(16);
output(0, 210) <= input(17);
output(0, 211) <= input(18);
output(0, 212) <= input(19);
output(0, 213) <= input(20);
output(0, 214) <= input(21);
output(0, 215) <= input(22);
output(0, 216) <= input(23);
output(0, 217) <= input(24);
output(0, 218) <= input(25);
output(0, 219) <= input(26);
output(0, 220) <= input(27);
output(0, 221) <= input(28);
output(0, 222) <= input(29);
output(0, 223) <= input(30);
output(0, 224) <= input(33);
output(0, 225) <= input(16);
output(0, 226) <= input(17);
output(0, 227) <= input(18);
output(0, 228) <= input(19);
output(0, 229) <= input(20);
output(0, 230) <= input(21);
output(0, 231) <= input(22);
output(0, 232) <= input(23);
output(0, 233) <= input(24);
output(0, 234) <= input(25);
output(0, 235) <= input(26);
output(0, 236) <= input(27);
output(0, 237) <= input(28);
output(0, 238) <= input(29);
output(0, 239) <= input(30);
output(0, 240) <= input(33);
output(0, 241) <= input(16);
output(0, 242) <= input(17);
output(0, 243) <= input(18);
output(0, 244) <= input(19);
output(0, 245) <= input(20);
output(0, 246) <= input(21);
output(0, 247) <= input(22);
output(0, 248) <= input(23);
output(0, 249) <= input(24);
output(0, 250) <= input(25);
output(0, 251) <= input(26);
output(0, 252) <= input(27);
output(0, 253) <= input(28);
output(0, 254) <= input(29);
output(0, 255) <= input(30);
output(1, 0) <= input(34);
output(1, 1) <= input(1);
output(1, 2) <= input(2);
output(1, 3) <= input(3);
output(1, 4) <= input(4);
output(1, 5) <= input(5);
output(1, 6) <= input(6);
output(1, 7) <= input(7);
output(1, 8) <= input(8);
output(1, 9) <= input(9);
output(1, 10) <= input(10);
output(1, 11) <= input(11);
output(1, 12) <= input(12);
output(1, 13) <= input(13);
output(1, 14) <= input(14);
output(1, 15) <= input(15);
output(1, 16) <= input(34);
output(1, 17) <= input(1);
output(1, 18) <= input(2);
output(1, 19) <= input(3);
output(1, 20) <= input(4);
output(1, 21) <= input(5);
output(1, 22) <= input(6);
output(1, 23) <= input(7);
output(1, 24) <= input(8);
output(1, 25) <= input(9);
output(1, 26) <= input(10);
output(1, 27) <= input(11);
output(1, 28) <= input(12);
output(1, 29) <= input(13);
output(1, 30) <= input(14);
output(1, 31) <= input(15);
output(1, 32) <= input(35);
output(1, 33) <= input(17);
output(1, 34) <= input(18);
output(1, 35) <= input(19);
output(1, 36) <= input(20);
output(1, 37) <= input(21);
output(1, 38) <= input(22);
output(1, 39) <= input(23);
output(1, 40) <= input(24);
output(1, 41) <= input(25);
output(1, 42) <= input(26);
output(1, 43) <= input(27);
output(1, 44) <= input(28);
output(1, 45) <= input(29);
output(1, 46) <= input(30);
output(1, 47) <= input(31);
output(1, 48) <= input(35);
output(1, 49) <= input(17);
output(1, 50) <= input(18);
output(1, 51) <= input(19);
output(1, 52) <= input(20);
output(1, 53) <= input(21);
output(1, 54) <= input(22);
output(1, 55) <= input(23);
output(1, 56) <= input(24);
output(1, 57) <= input(25);
output(1, 58) <= input(26);
output(1, 59) <= input(27);
output(1, 60) <= input(28);
output(1, 61) <= input(29);
output(1, 62) <= input(30);
output(1, 63) <= input(31);
output(1, 64) <= input(35);
output(1, 65) <= input(17);
output(1, 66) <= input(18);
output(1, 67) <= input(19);
output(1, 68) <= input(20);
output(1, 69) <= input(21);
output(1, 70) <= input(22);
output(1, 71) <= input(23);
output(1, 72) <= input(24);
output(1, 73) <= input(25);
output(1, 74) <= input(26);
output(1, 75) <= input(27);
output(1, 76) <= input(28);
output(1, 77) <= input(29);
output(1, 78) <= input(30);
output(1, 79) <= input(31);
output(1, 80) <= input(36);
output(1, 81) <= input(34);
output(1, 82) <= input(1);
output(1, 83) <= input(2);
output(1, 84) <= input(3);
output(1, 85) <= input(4);
output(1, 86) <= input(5);
output(1, 87) <= input(6);
output(1, 88) <= input(7);
output(1, 89) <= input(8);
output(1, 90) <= input(9);
output(1, 91) <= input(10);
output(1, 92) <= input(11);
output(1, 93) <= input(12);
output(1, 94) <= input(13);
output(1, 95) <= input(14);
output(1, 96) <= input(36);
output(1, 97) <= input(34);
output(1, 98) <= input(1);
output(1, 99) <= input(2);
output(1, 100) <= input(3);
output(1, 101) <= input(4);
output(1, 102) <= input(5);
output(1, 103) <= input(6);
output(1, 104) <= input(7);
output(1, 105) <= input(8);
output(1, 106) <= input(9);
output(1, 107) <= input(10);
output(1, 108) <= input(11);
output(1, 109) <= input(12);
output(1, 110) <= input(13);
output(1, 111) <= input(14);
output(1, 112) <= input(36);
output(1, 113) <= input(34);
output(1, 114) <= input(1);
output(1, 115) <= input(2);
output(1, 116) <= input(3);
output(1, 117) <= input(4);
output(1, 118) <= input(5);
output(1, 119) <= input(6);
output(1, 120) <= input(7);
output(1, 121) <= input(8);
output(1, 122) <= input(9);
output(1, 123) <= input(10);
output(1, 124) <= input(11);
output(1, 125) <= input(12);
output(1, 126) <= input(13);
output(1, 127) <= input(14);
output(1, 128) <= input(37);
output(1, 129) <= input(35);
output(1, 130) <= input(17);
output(1, 131) <= input(18);
output(1, 132) <= input(19);
output(1, 133) <= input(20);
output(1, 134) <= input(21);
output(1, 135) <= input(22);
output(1, 136) <= input(23);
output(1, 137) <= input(24);
output(1, 138) <= input(25);
output(1, 139) <= input(26);
output(1, 140) <= input(27);
output(1, 141) <= input(28);
output(1, 142) <= input(29);
output(1, 143) <= input(30);
output(1, 144) <= input(37);
output(1, 145) <= input(35);
output(1, 146) <= input(17);
output(1, 147) <= input(18);
output(1, 148) <= input(19);
output(1, 149) <= input(20);
output(1, 150) <= input(21);
output(1, 151) <= input(22);
output(1, 152) <= input(23);
output(1, 153) <= input(24);
output(1, 154) <= input(25);
output(1, 155) <= input(26);
output(1, 156) <= input(27);
output(1, 157) <= input(28);
output(1, 158) <= input(29);
output(1, 159) <= input(30);
output(1, 160) <= input(38);
output(1, 161) <= input(36);
output(1, 162) <= input(34);
output(1, 163) <= input(1);
output(1, 164) <= input(2);
output(1, 165) <= input(3);
output(1, 166) <= input(4);
output(1, 167) <= input(5);
output(1, 168) <= input(6);
output(1, 169) <= input(7);
output(1, 170) <= input(8);
output(1, 171) <= input(9);
output(1, 172) <= input(10);
output(1, 173) <= input(11);
output(1, 174) <= input(12);
output(1, 175) <= input(13);
output(1, 176) <= input(38);
output(1, 177) <= input(36);
output(1, 178) <= input(34);
output(1, 179) <= input(1);
output(1, 180) <= input(2);
output(1, 181) <= input(3);
output(1, 182) <= input(4);
output(1, 183) <= input(5);
output(1, 184) <= input(6);
output(1, 185) <= input(7);
output(1, 186) <= input(8);
output(1, 187) <= input(9);
output(1, 188) <= input(10);
output(1, 189) <= input(11);
output(1, 190) <= input(12);
output(1, 191) <= input(13);
output(1, 192) <= input(38);
output(1, 193) <= input(36);
output(1, 194) <= input(34);
output(1, 195) <= input(1);
output(1, 196) <= input(2);
output(1, 197) <= input(3);
output(1, 198) <= input(4);
output(1, 199) <= input(5);
output(1, 200) <= input(6);
output(1, 201) <= input(7);
output(1, 202) <= input(8);
output(1, 203) <= input(9);
output(1, 204) <= input(10);
output(1, 205) <= input(11);
output(1, 206) <= input(12);
output(1, 207) <= input(13);
output(1, 208) <= input(39);
output(1, 209) <= input(37);
output(1, 210) <= input(35);
output(1, 211) <= input(17);
output(1, 212) <= input(18);
output(1, 213) <= input(19);
output(1, 214) <= input(20);
output(1, 215) <= input(21);
output(1, 216) <= input(22);
output(1, 217) <= input(23);
output(1, 218) <= input(24);
output(1, 219) <= input(25);
output(1, 220) <= input(26);
output(1, 221) <= input(27);
output(1, 222) <= input(28);
output(1, 223) <= input(29);
output(1, 224) <= input(39);
output(1, 225) <= input(37);
output(1, 226) <= input(35);
output(1, 227) <= input(17);
output(1, 228) <= input(18);
output(1, 229) <= input(19);
output(1, 230) <= input(20);
output(1, 231) <= input(21);
output(1, 232) <= input(22);
output(1, 233) <= input(23);
output(1, 234) <= input(24);
output(1, 235) <= input(25);
output(1, 236) <= input(26);
output(1, 237) <= input(27);
output(1, 238) <= input(28);
output(1, 239) <= input(29);
output(1, 240) <= input(39);
output(1, 241) <= input(37);
output(1, 242) <= input(35);
output(1, 243) <= input(17);
output(1, 244) <= input(18);
output(1, 245) <= input(19);
output(1, 246) <= input(20);
output(1, 247) <= input(21);
output(1, 248) <= input(22);
output(1, 249) <= input(23);
output(1, 250) <= input(24);
output(1, 251) <= input(25);
output(1, 252) <= input(26);
output(1, 253) <= input(27);
output(1, 254) <= input(28);
output(1, 255) <= input(29);
output(2, 0) <= input(40);
output(2, 1) <= input(1);
output(2, 2) <= input(2);
output(2, 3) <= input(3);
output(2, 4) <= input(4);
output(2, 5) <= input(5);
output(2, 6) <= input(6);
output(2, 7) <= input(7);
output(2, 8) <= input(8);
output(2, 9) <= input(9);
output(2, 10) <= input(10);
output(2, 11) <= input(11);
output(2, 12) <= input(12);
output(2, 13) <= input(13);
output(2, 14) <= input(14);
output(2, 15) <= input(15);
output(2, 16) <= input(40);
output(2, 17) <= input(1);
output(2, 18) <= input(2);
output(2, 19) <= input(3);
output(2, 20) <= input(4);
output(2, 21) <= input(5);
output(2, 22) <= input(6);
output(2, 23) <= input(7);
output(2, 24) <= input(8);
output(2, 25) <= input(9);
output(2, 26) <= input(10);
output(2, 27) <= input(11);
output(2, 28) <= input(12);
output(2, 29) <= input(13);
output(2, 30) <= input(14);
output(2, 31) <= input(15);
output(2, 32) <= input(41);
output(2, 33) <= input(17);
output(2, 34) <= input(18);
output(2, 35) <= input(19);
output(2, 36) <= input(20);
output(2, 37) <= input(21);
output(2, 38) <= input(22);
output(2, 39) <= input(23);
output(2, 40) <= input(24);
output(2, 41) <= input(25);
output(2, 42) <= input(26);
output(2, 43) <= input(27);
output(2, 44) <= input(28);
output(2, 45) <= input(29);
output(2, 46) <= input(30);
output(2, 47) <= input(31);
output(2, 48) <= input(41);
output(2, 49) <= input(17);
output(2, 50) <= input(18);
output(2, 51) <= input(19);
output(2, 52) <= input(20);
output(2, 53) <= input(21);
output(2, 54) <= input(22);
output(2, 55) <= input(23);
output(2, 56) <= input(24);
output(2, 57) <= input(25);
output(2, 58) <= input(26);
output(2, 59) <= input(27);
output(2, 60) <= input(28);
output(2, 61) <= input(29);
output(2, 62) <= input(30);
output(2, 63) <= input(31);
output(2, 64) <= input(42);
output(2, 65) <= input(40);
output(2, 66) <= input(1);
output(2, 67) <= input(2);
output(2, 68) <= input(3);
output(2, 69) <= input(4);
output(2, 70) <= input(5);
output(2, 71) <= input(6);
output(2, 72) <= input(7);
output(2, 73) <= input(8);
output(2, 74) <= input(9);
output(2, 75) <= input(10);
output(2, 76) <= input(11);
output(2, 77) <= input(12);
output(2, 78) <= input(13);
output(2, 79) <= input(14);
output(2, 80) <= input(42);
output(2, 81) <= input(40);
output(2, 82) <= input(1);
output(2, 83) <= input(2);
output(2, 84) <= input(3);
output(2, 85) <= input(4);
output(2, 86) <= input(5);
output(2, 87) <= input(6);
output(2, 88) <= input(7);
output(2, 89) <= input(8);
output(2, 90) <= input(9);
output(2, 91) <= input(10);
output(2, 92) <= input(11);
output(2, 93) <= input(12);
output(2, 94) <= input(13);
output(2, 95) <= input(14);
output(2, 96) <= input(43);
output(2, 97) <= input(41);
output(2, 98) <= input(17);
output(2, 99) <= input(18);
output(2, 100) <= input(19);
output(2, 101) <= input(20);
output(2, 102) <= input(21);
output(2, 103) <= input(22);
output(2, 104) <= input(23);
output(2, 105) <= input(24);
output(2, 106) <= input(25);
output(2, 107) <= input(26);
output(2, 108) <= input(27);
output(2, 109) <= input(28);
output(2, 110) <= input(29);
output(2, 111) <= input(30);
output(2, 112) <= input(43);
output(2, 113) <= input(41);
output(2, 114) <= input(17);
output(2, 115) <= input(18);
output(2, 116) <= input(19);
output(2, 117) <= input(20);
output(2, 118) <= input(21);
output(2, 119) <= input(22);
output(2, 120) <= input(23);
output(2, 121) <= input(24);
output(2, 122) <= input(25);
output(2, 123) <= input(26);
output(2, 124) <= input(27);
output(2, 125) <= input(28);
output(2, 126) <= input(29);
output(2, 127) <= input(30);
output(2, 128) <= input(44);
output(2, 129) <= input(42);
output(2, 130) <= input(40);
output(2, 131) <= input(1);
output(2, 132) <= input(2);
output(2, 133) <= input(3);
output(2, 134) <= input(4);
output(2, 135) <= input(5);
output(2, 136) <= input(6);
output(2, 137) <= input(7);
output(2, 138) <= input(8);
output(2, 139) <= input(9);
output(2, 140) <= input(10);
output(2, 141) <= input(11);
output(2, 142) <= input(12);
output(2, 143) <= input(13);
output(2, 144) <= input(44);
output(2, 145) <= input(42);
output(2, 146) <= input(40);
output(2, 147) <= input(1);
output(2, 148) <= input(2);
output(2, 149) <= input(3);
output(2, 150) <= input(4);
output(2, 151) <= input(5);
output(2, 152) <= input(6);
output(2, 153) <= input(7);
output(2, 154) <= input(8);
output(2, 155) <= input(9);
output(2, 156) <= input(10);
output(2, 157) <= input(11);
output(2, 158) <= input(12);
output(2, 159) <= input(13);
output(2, 160) <= input(45);
output(2, 161) <= input(43);
output(2, 162) <= input(41);
output(2, 163) <= input(17);
output(2, 164) <= input(18);
output(2, 165) <= input(19);
output(2, 166) <= input(20);
output(2, 167) <= input(21);
output(2, 168) <= input(22);
output(2, 169) <= input(23);
output(2, 170) <= input(24);
output(2, 171) <= input(25);
output(2, 172) <= input(26);
output(2, 173) <= input(27);
output(2, 174) <= input(28);
output(2, 175) <= input(29);
output(2, 176) <= input(45);
output(2, 177) <= input(43);
output(2, 178) <= input(41);
output(2, 179) <= input(17);
output(2, 180) <= input(18);
output(2, 181) <= input(19);
output(2, 182) <= input(20);
output(2, 183) <= input(21);
output(2, 184) <= input(22);
output(2, 185) <= input(23);
output(2, 186) <= input(24);
output(2, 187) <= input(25);
output(2, 188) <= input(26);
output(2, 189) <= input(27);
output(2, 190) <= input(28);
output(2, 191) <= input(29);
output(2, 192) <= input(46);
output(2, 193) <= input(44);
output(2, 194) <= input(42);
output(2, 195) <= input(40);
output(2, 196) <= input(1);
output(2, 197) <= input(2);
output(2, 198) <= input(3);
output(2, 199) <= input(4);
output(2, 200) <= input(5);
output(2, 201) <= input(6);
output(2, 202) <= input(7);
output(2, 203) <= input(8);
output(2, 204) <= input(9);
output(2, 205) <= input(10);
output(2, 206) <= input(11);
output(2, 207) <= input(12);
output(2, 208) <= input(46);
output(2, 209) <= input(44);
output(2, 210) <= input(42);
output(2, 211) <= input(40);
output(2, 212) <= input(1);
output(2, 213) <= input(2);
output(2, 214) <= input(3);
output(2, 215) <= input(4);
output(2, 216) <= input(5);
output(2, 217) <= input(6);
output(2, 218) <= input(7);
output(2, 219) <= input(8);
output(2, 220) <= input(9);
output(2, 221) <= input(10);
output(2, 222) <= input(11);
output(2, 223) <= input(12);
output(2, 224) <= input(47);
output(2, 225) <= input(45);
output(2, 226) <= input(43);
output(2, 227) <= input(41);
output(2, 228) <= input(17);
output(2, 229) <= input(18);
output(2, 230) <= input(19);
output(2, 231) <= input(20);
output(2, 232) <= input(21);
output(2, 233) <= input(22);
output(2, 234) <= input(23);
output(2, 235) <= input(24);
output(2, 236) <= input(25);
output(2, 237) <= input(26);
output(2, 238) <= input(27);
output(2, 239) <= input(28);
output(2, 240) <= input(47);
output(2, 241) <= input(45);
output(2, 242) <= input(43);
output(2, 243) <= input(41);
output(2, 244) <= input(17);
output(2, 245) <= input(18);
output(2, 246) <= input(19);
output(2, 247) <= input(20);
output(2, 248) <= input(21);
output(2, 249) <= input(22);
output(2, 250) <= input(23);
output(2, 251) <= input(24);
output(2, 252) <= input(25);
output(2, 253) <= input(26);
output(2, 254) <= input(27);
output(2, 255) <= input(28);
when "0100" =>
output(0, 0) <= input(0);
output(0, 1) <= input(1);
output(0, 2) <= input(2);
output(0, 3) <= input(3);
output(0, 4) <= input(4);
output(0, 5) <= input(5);
output(0, 6) <= input(6);
output(0, 7) <= input(7);
output(0, 8) <= input(8);
output(0, 9) <= input(9);
output(0, 10) <= input(10);
output(0, 11) <= input(11);
output(0, 12) <= input(12);
output(0, 13) <= input(13);
output(0, 14) <= input(14);
output(0, 15) <= input(15);
output(0, 16) <= input(16);
output(0, 17) <= input(17);
output(0, 18) <= input(18);
output(0, 19) <= input(19);
output(0, 20) <= input(20);
output(0, 21) <= input(21);
output(0, 22) <= input(22);
output(0, 23) <= input(23);
output(0, 24) <= input(24);
output(0, 25) <= input(25);
output(0, 26) <= input(26);
output(0, 27) <= input(27);
output(0, 28) <= input(28);
output(0, 29) <= input(29);
output(0, 30) <= input(30);
output(0, 31) <= input(31);
output(0, 32) <= input(16);
output(0, 33) <= input(17);
output(0, 34) <= input(18);
output(0, 35) <= input(19);
output(0, 36) <= input(20);
output(0, 37) <= input(21);
output(0, 38) <= input(22);
output(0, 39) <= input(23);
output(0, 40) <= input(24);
output(0, 41) <= input(25);
output(0, 42) <= input(26);
output(0, 43) <= input(27);
output(0, 44) <= input(28);
output(0, 45) <= input(29);
output(0, 46) <= input(30);
output(0, 47) <= input(31);
output(0, 48) <= input(32);
output(0, 49) <= input(0);
output(0, 50) <= input(1);
output(0, 51) <= input(2);
output(0, 52) <= input(3);
output(0, 53) <= input(4);
output(0, 54) <= input(5);
output(0, 55) <= input(6);
output(0, 56) <= input(7);
output(0, 57) <= input(8);
output(0, 58) <= input(9);
output(0, 59) <= input(10);
output(0, 60) <= input(11);
output(0, 61) <= input(12);
output(0, 62) <= input(13);
output(0, 63) <= input(14);
output(0, 64) <= input(33);
output(0, 65) <= input(16);
output(0, 66) <= input(17);
output(0, 67) <= input(18);
output(0, 68) <= input(19);
output(0, 69) <= input(20);
output(0, 70) <= input(21);
output(0, 71) <= input(22);
output(0, 72) <= input(23);
output(0, 73) <= input(24);
output(0, 74) <= input(25);
output(0, 75) <= input(26);
output(0, 76) <= input(27);
output(0, 77) <= input(28);
output(0, 78) <= input(29);
output(0, 79) <= input(30);
output(0, 80) <= input(33);
output(0, 81) <= input(16);
output(0, 82) <= input(17);
output(0, 83) <= input(18);
output(0, 84) <= input(19);
output(0, 85) <= input(20);
output(0, 86) <= input(21);
output(0, 87) <= input(22);
output(0, 88) <= input(23);
output(0, 89) <= input(24);
output(0, 90) <= input(25);
output(0, 91) <= input(26);
output(0, 92) <= input(27);
output(0, 93) <= input(28);
output(0, 94) <= input(29);
output(0, 95) <= input(30);
output(0, 96) <= input(34);
output(0, 97) <= input(32);
output(0, 98) <= input(0);
output(0, 99) <= input(1);
output(0, 100) <= input(2);
output(0, 101) <= input(3);
output(0, 102) <= input(4);
output(0, 103) <= input(5);
output(0, 104) <= input(6);
output(0, 105) <= input(7);
output(0, 106) <= input(8);
output(0, 107) <= input(9);
output(0, 108) <= input(10);
output(0, 109) <= input(11);
output(0, 110) <= input(12);
output(0, 111) <= input(13);
output(0, 112) <= input(34);
output(0, 113) <= input(32);
output(0, 114) <= input(0);
output(0, 115) <= input(1);
output(0, 116) <= input(2);
output(0, 117) <= input(3);
output(0, 118) <= input(4);
output(0, 119) <= input(5);
output(0, 120) <= input(6);
output(0, 121) <= input(7);
output(0, 122) <= input(8);
output(0, 123) <= input(9);
output(0, 124) <= input(10);
output(0, 125) <= input(11);
output(0, 126) <= input(12);
output(0, 127) <= input(13);
output(0, 128) <= input(35);
output(0, 129) <= input(33);
output(0, 130) <= input(16);
output(0, 131) <= input(17);
output(0, 132) <= input(18);
output(0, 133) <= input(19);
output(0, 134) <= input(20);
output(0, 135) <= input(21);
output(0, 136) <= input(22);
output(0, 137) <= input(23);
output(0, 138) <= input(24);
output(0, 139) <= input(25);
output(0, 140) <= input(26);
output(0, 141) <= input(27);
output(0, 142) <= input(28);
output(0, 143) <= input(29);
output(0, 144) <= input(36);
output(0, 145) <= input(34);
output(0, 146) <= input(32);
output(0, 147) <= input(0);
output(0, 148) <= input(1);
output(0, 149) <= input(2);
output(0, 150) <= input(3);
output(0, 151) <= input(4);
output(0, 152) <= input(5);
output(0, 153) <= input(6);
output(0, 154) <= input(7);
output(0, 155) <= input(8);
output(0, 156) <= input(9);
output(0, 157) <= input(10);
output(0, 158) <= input(11);
output(0, 159) <= input(12);
output(0, 160) <= input(36);
output(0, 161) <= input(34);
output(0, 162) <= input(32);
output(0, 163) <= input(0);
output(0, 164) <= input(1);
output(0, 165) <= input(2);
output(0, 166) <= input(3);
output(0, 167) <= input(4);
output(0, 168) <= input(5);
output(0, 169) <= input(6);
output(0, 170) <= input(7);
output(0, 171) <= input(8);
output(0, 172) <= input(9);
output(0, 173) <= input(10);
output(0, 174) <= input(11);
output(0, 175) <= input(12);
output(0, 176) <= input(37);
output(0, 177) <= input(35);
output(0, 178) <= input(33);
output(0, 179) <= input(16);
output(0, 180) <= input(17);
output(0, 181) <= input(18);
output(0, 182) <= input(19);
output(0, 183) <= input(20);
output(0, 184) <= input(21);
output(0, 185) <= input(22);
output(0, 186) <= input(23);
output(0, 187) <= input(24);
output(0, 188) <= input(25);
output(0, 189) <= input(26);
output(0, 190) <= input(27);
output(0, 191) <= input(28);
output(0, 192) <= input(38);
output(0, 193) <= input(36);
output(0, 194) <= input(34);
output(0, 195) <= input(32);
output(0, 196) <= input(0);
output(0, 197) <= input(1);
output(0, 198) <= input(2);
output(0, 199) <= input(3);
output(0, 200) <= input(4);
output(0, 201) <= input(5);
output(0, 202) <= input(6);
output(0, 203) <= input(7);
output(0, 204) <= input(8);
output(0, 205) <= input(9);
output(0, 206) <= input(10);
output(0, 207) <= input(11);
output(0, 208) <= input(38);
output(0, 209) <= input(36);
output(0, 210) <= input(34);
output(0, 211) <= input(32);
output(0, 212) <= input(0);
output(0, 213) <= input(1);
output(0, 214) <= input(2);
output(0, 215) <= input(3);
output(0, 216) <= input(4);
output(0, 217) <= input(5);
output(0, 218) <= input(6);
output(0, 219) <= input(7);
output(0, 220) <= input(8);
output(0, 221) <= input(9);
output(0, 222) <= input(10);
output(0, 223) <= input(11);
output(0, 224) <= input(39);
output(0, 225) <= input(37);
output(0, 226) <= input(35);
output(0, 227) <= input(33);
output(0, 228) <= input(16);
output(0, 229) <= input(17);
output(0, 230) <= input(18);
output(0, 231) <= input(19);
output(0, 232) <= input(20);
output(0, 233) <= input(21);
output(0, 234) <= input(22);
output(0, 235) <= input(23);
output(0, 236) <= input(24);
output(0, 237) <= input(25);
output(0, 238) <= input(26);
output(0, 239) <= input(27);
output(0, 240) <= input(39);
output(0, 241) <= input(37);
output(0, 242) <= input(35);
output(0, 243) <= input(33);
output(0, 244) <= input(16);
output(0, 245) <= input(17);
output(0, 246) <= input(18);
output(0, 247) <= input(19);
output(0, 248) <= input(20);
output(0, 249) <= input(21);
output(0, 250) <= input(22);
output(0, 251) <= input(23);
output(0, 252) <= input(24);
output(0, 253) <= input(25);
output(0, 254) <= input(26);
output(0, 255) <= input(27);
output(1, 0) <= input(0);
output(1, 1) <= input(1);
output(1, 2) <= input(2);
output(1, 3) <= input(3);
output(1, 4) <= input(4);
output(1, 5) <= input(5);
output(1, 6) <= input(6);
output(1, 7) <= input(7);
output(1, 8) <= input(8);
output(1, 9) <= input(9);
output(1, 10) <= input(10);
output(1, 11) <= input(11);
output(1, 12) <= input(12);
output(1, 13) <= input(13);
output(1, 14) <= input(14);
output(1, 15) <= input(15);
output(1, 16) <= input(16);
output(1, 17) <= input(17);
output(1, 18) <= input(18);
output(1, 19) <= input(19);
output(1, 20) <= input(20);
output(1, 21) <= input(21);
output(1, 22) <= input(22);
output(1, 23) <= input(23);
output(1, 24) <= input(24);
output(1, 25) <= input(25);
output(1, 26) <= input(26);
output(1, 27) <= input(27);
output(1, 28) <= input(28);
output(1, 29) <= input(29);
output(1, 30) <= input(30);
output(1, 31) <= input(31);
output(1, 32) <= input(40);
output(1, 33) <= input(0);
output(1, 34) <= input(1);
output(1, 35) <= input(2);
output(1, 36) <= input(3);
output(1, 37) <= input(4);
output(1, 38) <= input(5);
output(1, 39) <= input(6);
output(1, 40) <= input(7);
output(1, 41) <= input(8);
output(1, 42) <= input(9);
output(1, 43) <= input(10);
output(1, 44) <= input(11);
output(1, 45) <= input(12);
output(1, 46) <= input(13);
output(1, 47) <= input(14);
output(1, 48) <= input(40);
output(1, 49) <= input(0);
output(1, 50) <= input(1);
output(1, 51) <= input(2);
output(1, 52) <= input(3);
output(1, 53) <= input(4);
output(1, 54) <= input(5);
output(1, 55) <= input(6);
output(1, 56) <= input(7);
output(1, 57) <= input(8);
output(1, 58) <= input(9);
output(1, 59) <= input(10);
output(1, 60) <= input(11);
output(1, 61) <= input(12);
output(1, 62) <= input(13);
output(1, 63) <= input(14);
output(1, 64) <= input(41);
output(1, 65) <= input(16);
output(1, 66) <= input(17);
output(1, 67) <= input(18);
output(1, 68) <= input(19);
output(1, 69) <= input(20);
output(1, 70) <= input(21);
output(1, 71) <= input(22);
output(1, 72) <= input(23);
output(1, 73) <= input(24);
output(1, 74) <= input(25);
output(1, 75) <= input(26);
output(1, 76) <= input(27);
output(1, 77) <= input(28);
output(1, 78) <= input(29);
output(1, 79) <= input(30);
output(1, 80) <= input(42);
output(1, 81) <= input(40);
output(1, 82) <= input(0);
output(1, 83) <= input(1);
output(1, 84) <= input(2);
output(1, 85) <= input(3);
output(1, 86) <= input(4);
output(1, 87) <= input(5);
output(1, 88) <= input(6);
output(1, 89) <= input(7);
output(1, 90) <= input(8);
output(1, 91) <= input(9);
output(1, 92) <= input(10);
output(1, 93) <= input(11);
output(1, 94) <= input(12);
output(1, 95) <= input(13);
output(1, 96) <= input(43);
output(1, 97) <= input(41);
output(1, 98) <= input(16);
output(1, 99) <= input(17);
output(1, 100) <= input(18);
output(1, 101) <= input(19);
output(1, 102) <= input(20);
output(1, 103) <= input(21);
output(1, 104) <= input(22);
output(1, 105) <= input(23);
output(1, 106) <= input(24);
output(1, 107) <= input(25);
output(1, 108) <= input(26);
output(1, 109) <= input(27);
output(1, 110) <= input(28);
output(1, 111) <= input(29);
output(1, 112) <= input(43);
output(1, 113) <= input(41);
output(1, 114) <= input(16);
output(1, 115) <= input(17);
output(1, 116) <= input(18);
output(1, 117) <= input(19);
output(1, 118) <= input(20);
output(1, 119) <= input(21);
output(1, 120) <= input(22);
output(1, 121) <= input(23);
output(1, 122) <= input(24);
output(1, 123) <= input(25);
output(1, 124) <= input(26);
output(1, 125) <= input(27);
output(1, 126) <= input(28);
output(1, 127) <= input(29);
output(1, 128) <= input(44);
output(1, 129) <= input(42);
output(1, 130) <= input(40);
output(1, 131) <= input(0);
output(1, 132) <= input(1);
output(1, 133) <= input(2);
output(1, 134) <= input(3);
output(1, 135) <= input(4);
output(1, 136) <= input(5);
output(1, 137) <= input(6);
output(1, 138) <= input(7);
output(1, 139) <= input(8);
output(1, 140) <= input(9);
output(1, 141) <= input(10);
output(1, 142) <= input(11);
output(1, 143) <= input(12);
output(1, 144) <= input(45);
output(1, 145) <= input(43);
output(1, 146) <= input(41);
output(1, 147) <= input(16);
output(1, 148) <= input(17);
output(1, 149) <= input(18);
output(1, 150) <= input(19);
output(1, 151) <= input(20);
output(1, 152) <= input(21);
output(1, 153) <= input(22);
output(1, 154) <= input(23);
output(1, 155) <= input(24);
output(1, 156) <= input(25);
output(1, 157) <= input(26);
output(1, 158) <= input(27);
output(1, 159) <= input(28);
output(1, 160) <= input(46);
output(1, 161) <= input(44);
output(1, 162) <= input(42);
output(1, 163) <= input(40);
output(1, 164) <= input(0);
output(1, 165) <= input(1);
output(1, 166) <= input(2);
output(1, 167) <= input(3);
output(1, 168) <= input(4);
output(1, 169) <= input(5);
output(1, 170) <= input(6);
output(1, 171) <= input(7);
output(1, 172) <= input(8);
output(1, 173) <= input(9);
output(1, 174) <= input(10);
output(1, 175) <= input(11);
output(1, 176) <= input(46);
output(1, 177) <= input(44);
output(1, 178) <= input(42);
output(1, 179) <= input(40);
output(1, 180) <= input(0);
output(1, 181) <= input(1);
output(1, 182) <= input(2);
output(1, 183) <= input(3);
output(1, 184) <= input(4);
output(1, 185) <= input(5);
output(1, 186) <= input(6);
output(1, 187) <= input(7);
output(1, 188) <= input(8);
output(1, 189) <= input(9);
output(1, 190) <= input(10);
output(1, 191) <= input(11);
output(1, 192) <= input(47);
output(1, 193) <= input(45);
output(1, 194) <= input(43);
output(1, 195) <= input(41);
output(1, 196) <= input(16);
output(1, 197) <= input(17);
output(1, 198) <= input(18);
output(1, 199) <= input(19);
output(1, 200) <= input(20);
output(1, 201) <= input(21);
output(1, 202) <= input(22);
output(1, 203) <= input(23);
output(1, 204) <= input(24);
output(1, 205) <= input(25);
output(1, 206) <= input(26);
output(1, 207) <= input(27);
output(1, 208) <= input(48);
output(1, 209) <= input(46);
output(1, 210) <= input(44);
output(1, 211) <= input(42);
output(1, 212) <= input(40);
output(1, 213) <= input(0);
output(1, 214) <= input(1);
output(1, 215) <= input(2);
output(1, 216) <= input(3);
output(1, 217) <= input(4);
output(1, 218) <= input(5);
output(1, 219) <= input(6);
output(1, 220) <= input(7);
output(1, 221) <= input(8);
output(1, 222) <= input(9);
output(1, 223) <= input(10);
output(1, 224) <= input(49);
output(1, 225) <= input(47);
output(1, 226) <= input(45);
output(1, 227) <= input(43);
output(1, 228) <= input(41);
output(1, 229) <= input(16);
output(1, 230) <= input(17);
output(1, 231) <= input(18);
output(1, 232) <= input(19);
output(1, 233) <= input(20);
output(1, 234) <= input(21);
output(1, 235) <= input(22);
output(1, 236) <= input(23);
output(1, 237) <= input(24);
output(1, 238) <= input(25);
output(1, 239) <= input(26);
output(1, 240) <= input(49);
output(1, 241) <= input(47);
output(1, 242) <= input(45);
output(1, 243) <= input(43);
output(1, 244) <= input(41);
output(1, 245) <= input(16);
output(1, 246) <= input(17);
output(1, 247) <= input(18);
output(1, 248) <= input(19);
output(1, 249) <= input(20);
output(1, 250) <= input(21);
output(1, 251) <= input(22);
output(1, 252) <= input(23);
output(1, 253) <= input(24);
output(1, 254) <= input(25);
output(1, 255) <= input(26);
output(2, 0) <= input(50);
output(2, 1) <= input(1);
output(2, 2) <= input(2);
output(2, 3) <= input(3);
output(2, 4) <= input(4);
output(2, 5) <= input(5);
output(2, 6) <= input(6);
output(2, 7) <= input(7);
output(2, 8) <= input(8);
output(2, 9) <= input(9);
output(2, 10) <= input(10);
output(2, 11) <= input(11);
output(2, 12) <= input(12);
output(2, 13) <= input(13);
output(2, 14) <= input(14);
output(2, 15) <= input(15);
output(2, 16) <= input(51);
output(2, 17) <= input(17);
output(2, 18) <= input(18);
output(2, 19) <= input(19);
output(2, 20) <= input(20);
output(2, 21) <= input(21);
output(2, 22) <= input(22);
output(2, 23) <= input(23);
output(2, 24) <= input(24);
output(2, 25) <= input(25);
output(2, 26) <= input(26);
output(2, 27) <= input(27);
output(2, 28) <= input(28);
output(2, 29) <= input(29);
output(2, 30) <= input(30);
output(2, 31) <= input(31);
output(2, 32) <= input(52);
output(2, 33) <= input(50);
output(2, 34) <= input(1);
output(2, 35) <= input(2);
output(2, 36) <= input(3);
output(2, 37) <= input(4);
output(2, 38) <= input(5);
output(2, 39) <= input(6);
output(2, 40) <= input(7);
output(2, 41) <= input(8);
output(2, 42) <= input(9);
output(2, 43) <= input(10);
output(2, 44) <= input(11);
output(2, 45) <= input(12);
output(2, 46) <= input(13);
output(2, 47) <= input(14);
output(2, 48) <= input(53);
output(2, 49) <= input(51);
output(2, 50) <= input(17);
output(2, 51) <= input(18);
output(2, 52) <= input(19);
output(2, 53) <= input(20);
output(2, 54) <= input(21);
output(2, 55) <= input(22);
output(2, 56) <= input(23);
output(2, 57) <= input(24);
output(2, 58) <= input(25);
output(2, 59) <= input(26);
output(2, 60) <= input(27);
output(2, 61) <= input(28);
output(2, 62) <= input(29);
output(2, 63) <= input(30);
output(2, 64) <= input(54);
output(2, 65) <= input(52);
output(2, 66) <= input(50);
output(2, 67) <= input(1);
output(2, 68) <= input(2);
output(2, 69) <= input(3);
output(2, 70) <= input(4);
output(2, 71) <= input(5);
output(2, 72) <= input(6);
output(2, 73) <= input(7);
output(2, 74) <= input(8);
output(2, 75) <= input(9);
output(2, 76) <= input(10);
output(2, 77) <= input(11);
output(2, 78) <= input(12);
output(2, 79) <= input(13);
output(2, 80) <= input(55);
output(2, 81) <= input(53);
output(2, 82) <= input(51);
output(2, 83) <= input(17);
output(2, 84) <= input(18);
output(2, 85) <= input(19);
output(2, 86) <= input(20);
output(2, 87) <= input(21);
output(2, 88) <= input(22);
output(2, 89) <= input(23);
output(2, 90) <= input(24);
output(2, 91) <= input(25);
output(2, 92) <= input(26);
output(2, 93) <= input(27);
output(2, 94) <= input(28);
output(2, 95) <= input(29);
output(2, 96) <= input(56);
output(2, 97) <= input(54);
output(2, 98) <= input(52);
output(2, 99) <= input(50);
output(2, 100) <= input(1);
output(2, 101) <= input(2);
output(2, 102) <= input(3);
output(2, 103) <= input(4);
output(2, 104) <= input(5);
output(2, 105) <= input(6);
output(2, 106) <= input(7);
output(2, 107) <= input(8);
output(2, 108) <= input(9);
output(2, 109) <= input(10);
output(2, 110) <= input(11);
output(2, 111) <= input(12);
output(2, 112) <= input(56);
output(2, 113) <= input(54);
output(2, 114) <= input(52);
output(2, 115) <= input(50);
output(2, 116) <= input(1);
output(2, 117) <= input(2);
output(2, 118) <= input(3);
output(2, 119) <= input(4);
output(2, 120) <= input(5);
output(2, 121) <= input(6);
output(2, 122) <= input(7);
output(2, 123) <= input(8);
output(2, 124) <= input(9);
output(2, 125) <= input(10);
output(2, 126) <= input(11);
output(2, 127) <= input(12);
output(2, 128) <= input(57);
output(2, 129) <= input(55);
output(2, 130) <= input(53);
output(2, 131) <= input(51);
output(2, 132) <= input(17);
output(2, 133) <= input(18);
output(2, 134) <= input(19);
output(2, 135) <= input(20);
output(2, 136) <= input(21);
output(2, 137) <= input(22);
output(2, 138) <= input(23);
output(2, 139) <= input(24);
output(2, 140) <= input(25);
output(2, 141) <= input(26);
output(2, 142) <= input(27);
output(2, 143) <= input(28);
output(2, 144) <= input(58);
output(2, 145) <= input(56);
output(2, 146) <= input(54);
output(2, 147) <= input(52);
output(2, 148) <= input(50);
output(2, 149) <= input(1);
output(2, 150) <= input(2);
output(2, 151) <= input(3);
output(2, 152) <= input(4);
output(2, 153) <= input(5);
output(2, 154) <= input(6);
output(2, 155) <= input(7);
output(2, 156) <= input(8);
output(2, 157) <= input(9);
output(2, 158) <= input(10);
output(2, 159) <= input(11);
output(2, 160) <= input(59);
output(2, 161) <= input(57);
output(2, 162) <= input(55);
output(2, 163) <= input(53);
output(2, 164) <= input(51);
output(2, 165) <= input(17);
output(2, 166) <= input(18);
output(2, 167) <= input(19);
output(2, 168) <= input(20);
output(2, 169) <= input(21);
output(2, 170) <= input(22);
output(2, 171) <= input(23);
output(2, 172) <= input(24);
output(2, 173) <= input(25);
output(2, 174) <= input(26);
output(2, 175) <= input(27);
output(2, 176) <= input(60);
output(2, 177) <= input(58);
output(2, 178) <= input(56);
output(2, 179) <= input(54);
output(2, 180) <= input(52);
output(2, 181) <= input(50);
output(2, 182) <= input(1);
output(2, 183) <= input(2);
output(2, 184) <= input(3);
output(2, 185) <= input(4);
output(2, 186) <= input(5);
output(2, 187) <= input(6);
output(2, 188) <= input(7);
output(2, 189) <= input(8);
output(2, 190) <= input(9);
output(2, 191) <= input(10);
output(2, 192) <= input(61);
output(2, 193) <= input(59);
output(2, 194) <= input(57);
output(2, 195) <= input(55);
output(2, 196) <= input(53);
output(2, 197) <= input(51);
output(2, 198) <= input(17);
output(2, 199) <= input(18);
output(2, 200) <= input(19);
output(2, 201) <= input(20);
output(2, 202) <= input(21);
output(2, 203) <= input(22);
output(2, 204) <= input(23);
output(2, 205) <= input(24);
output(2, 206) <= input(25);
output(2, 207) <= input(26);
output(2, 208) <= input(62);
output(2, 209) <= input(60);
output(2, 210) <= input(58);
output(2, 211) <= input(56);
output(2, 212) <= input(54);
output(2, 213) <= input(52);
output(2, 214) <= input(50);
output(2, 215) <= input(1);
output(2, 216) <= input(2);
output(2, 217) <= input(3);
output(2, 218) <= input(4);
output(2, 219) <= input(5);
output(2, 220) <= input(6);
output(2, 221) <= input(7);
output(2, 222) <= input(8);
output(2, 223) <= input(9);
output(2, 224) <= input(63);
output(2, 225) <= input(61);
output(2, 226) <= input(59);
output(2, 227) <= input(57);
output(2, 228) <= input(55);
output(2, 229) <= input(53);
output(2, 230) <= input(51);
output(2, 231) <= input(17);
output(2, 232) <= input(18);
output(2, 233) <= input(19);
output(2, 234) <= input(20);
output(2, 235) <= input(21);
output(2, 236) <= input(22);
output(2, 237) <= input(23);
output(2, 238) <= input(24);
output(2, 239) <= input(25);
output(2, 240) <= input(63);
output(2, 241) <= input(61);
output(2, 242) <= input(59);
output(2, 243) <= input(57);
output(2, 244) <= input(55);
output(2, 245) <= input(53);
output(2, 246) <= input(51);
output(2, 247) <= input(17);
output(2, 248) <= input(18);
output(2, 249) <= input(19);
output(2, 250) <= input(20);
output(2, 251) <= input(21);
output(2, 252) <= input(22);
output(2, 253) <= input(23);
output(2, 254) <= input(24);
output(2, 255) <= input(25);
when "0101" =>
output(0, 0) <= input(0);
output(0, 1) <= input(1);
output(0, 2) <= input(2);
output(0, 3) <= input(3);
output(0, 4) <= input(4);
output(0, 5) <= input(5);
output(0, 6) <= input(6);
output(0, 7) <= input(7);
output(0, 8) <= input(8);
output(0, 9) <= input(9);
output(0, 10) <= input(10);
output(0, 11) <= input(11);
output(0, 12) <= input(12);
output(0, 13) <= input(13);
output(0, 14) <= input(14);
output(0, 15) <= input(15);
output(0, 16) <= input(16);
output(0, 17) <= input(17);
output(0, 18) <= input(18);
output(0, 19) <= input(19);
output(0, 20) <= input(20);
output(0, 21) <= input(21);
output(0, 22) <= input(22);
output(0, 23) <= input(23);
output(0, 24) <= input(24);
output(0, 25) <= input(25);
output(0, 26) <= input(26);
output(0, 27) <= input(27);
output(0, 28) <= input(28);
output(0, 29) <= input(29);
output(0, 30) <= input(30);
output(0, 31) <= input(31);
output(0, 32) <= input(32);
output(0, 33) <= input(0);
output(0, 34) <= input(1);
output(0, 35) <= input(2);
output(0, 36) <= input(3);
output(0, 37) <= input(4);
output(0, 38) <= input(5);
output(0, 39) <= input(6);
output(0, 40) <= input(7);
output(0, 41) <= input(8);
output(0, 42) <= input(9);
output(0, 43) <= input(10);
output(0, 44) <= input(11);
output(0, 45) <= input(12);
output(0, 46) <= input(13);
output(0, 47) <= input(14);
output(0, 48) <= input(33);
output(0, 49) <= input(16);
output(0, 50) <= input(17);
output(0, 51) <= input(18);
output(0, 52) <= input(19);
output(0, 53) <= input(20);
output(0, 54) <= input(21);
output(0, 55) <= input(22);
output(0, 56) <= input(23);
output(0, 57) <= input(24);
output(0, 58) <= input(25);
output(0, 59) <= input(26);
output(0, 60) <= input(27);
output(0, 61) <= input(28);
output(0, 62) <= input(29);
output(0, 63) <= input(30);
output(0, 64) <= input(34);
output(0, 65) <= input(32);
output(0, 66) <= input(0);
output(0, 67) <= input(1);
output(0, 68) <= input(2);
output(0, 69) <= input(3);
output(0, 70) <= input(4);
output(0, 71) <= input(5);
output(0, 72) <= input(6);
output(0, 73) <= input(7);
output(0, 74) <= input(8);
output(0, 75) <= input(9);
output(0, 76) <= input(10);
output(0, 77) <= input(11);
output(0, 78) <= input(12);
output(0, 79) <= input(13);
output(0, 80) <= input(35);
output(0, 81) <= input(33);
output(0, 82) <= input(16);
output(0, 83) <= input(17);
output(0, 84) <= input(18);
output(0, 85) <= input(19);
output(0, 86) <= input(20);
output(0, 87) <= input(21);
output(0, 88) <= input(22);
output(0, 89) <= input(23);
output(0, 90) <= input(24);
output(0, 91) <= input(25);
output(0, 92) <= input(26);
output(0, 93) <= input(27);
output(0, 94) <= input(28);
output(0, 95) <= input(29);
output(0, 96) <= input(36);
output(0, 97) <= input(34);
output(0, 98) <= input(32);
output(0, 99) <= input(0);
output(0, 100) <= input(1);
output(0, 101) <= input(2);
output(0, 102) <= input(3);
output(0, 103) <= input(4);
output(0, 104) <= input(5);
output(0, 105) <= input(6);
output(0, 106) <= input(7);
output(0, 107) <= input(8);
output(0, 108) <= input(9);
output(0, 109) <= input(10);
output(0, 110) <= input(11);
output(0, 111) <= input(12);
output(0, 112) <= input(37);
output(0, 113) <= input(35);
output(0, 114) <= input(33);
output(0, 115) <= input(16);
output(0, 116) <= input(17);
output(0, 117) <= input(18);
output(0, 118) <= input(19);
output(0, 119) <= input(20);
output(0, 120) <= input(21);
output(0, 121) <= input(22);
output(0, 122) <= input(23);
output(0, 123) <= input(24);
output(0, 124) <= input(25);
output(0, 125) <= input(26);
output(0, 126) <= input(27);
output(0, 127) <= input(28);
output(0, 128) <= input(38);
output(0, 129) <= input(36);
output(0, 130) <= input(34);
output(0, 131) <= input(32);
output(0, 132) <= input(0);
output(0, 133) <= input(1);
output(0, 134) <= input(2);
output(0, 135) <= input(3);
output(0, 136) <= input(4);
output(0, 137) <= input(5);
output(0, 138) <= input(6);
output(0, 139) <= input(7);
output(0, 140) <= input(8);
output(0, 141) <= input(9);
output(0, 142) <= input(10);
output(0, 143) <= input(11);
output(0, 144) <= input(39);
output(0, 145) <= input(37);
output(0, 146) <= input(35);
output(0, 147) <= input(33);
output(0, 148) <= input(16);
output(0, 149) <= input(17);
output(0, 150) <= input(18);
output(0, 151) <= input(19);
output(0, 152) <= input(20);
output(0, 153) <= input(21);
output(0, 154) <= input(22);
output(0, 155) <= input(23);
output(0, 156) <= input(24);
output(0, 157) <= input(25);
output(0, 158) <= input(26);
output(0, 159) <= input(27);
output(0, 160) <= input(40);
output(0, 161) <= input(38);
output(0, 162) <= input(36);
output(0, 163) <= input(34);
output(0, 164) <= input(32);
output(0, 165) <= input(0);
output(0, 166) <= input(1);
output(0, 167) <= input(2);
output(0, 168) <= input(3);
output(0, 169) <= input(4);
output(0, 170) <= input(5);
output(0, 171) <= input(6);
output(0, 172) <= input(7);
output(0, 173) <= input(8);
output(0, 174) <= input(9);
output(0, 175) <= input(10);
output(0, 176) <= input(41);
output(0, 177) <= input(39);
output(0, 178) <= input(37);
output(0, 179) <= input(35);
output(0, 180) <= input(33);
output(0, 181) <= input(16);
output(0, 182) <= input(17);
output(0, 183) <= input(18);
output(0, 184) <= input(19);
output(0, 185) <= input(20);
output(0, 186) <= input(21);
output(0, 187) <= input(22);
output(0, 188) <= input(23);
output(0, 189) <= input(24);
output(0, 190) <= input(25);
output(0, 191) <= input(26);
output(0, 192) <= input(42);
output(0, 193) <= input(40);
output(0, 194) <= input(38);
output(0, 195) <= input(36);
output(0, 196) <= input(34);
output(0, 197) <= input(32);
output(0, 198) <= input(0);
output(0, 199) <= input(1);
output(0, 200) <= input(2);
output(0, 201) <= input(3);
output(0, 202) <= input(4);
output(0, 203) <= input(5);
output(0, 204) <= input(6);
output(0, 205) <= input(7);
output(0, 206) <= input(8);
output(0, 207) <= input(9);
output(0, 208) <= input(43);
output(0, 209) <= input(41);
output(0, 210) <= input(39);
output(0, 211) <= input(37);
output(0, 212) <= input(35);
output(0, 213) <= input(33);
output(0, 214) <= input(16);
output(0, 215) <= input(17);
output(0, 216) <= input(18);
output(0, 217) <= input(19);
output(0, 218) <= input(20);
output(0, 219) <= input(21);
output(0, 220) <= input(22);
output(0, 221) <= input(23);
output(0, 222) <= input(24);
output(0, 223) <= input(25);
output(0, 224) <= input(44);
output(0, 225) <= input(42);
output(0, 226) <= input(40);
output(0, 227) <= input(38);
output(0, 228) <= input(36);
output(0, 229) <= input(34);
output(0, 230) <= input(32);
output(0, 231) <= input(0);
output(0, 232) <= input(1);
output(0, 233) <= input(2);
output(0, 234) <= input(3);
output(0, 235) <= input(4);
output(0, 236) <= input(5);
output(0, 237) <= input(6);
output(0, 238) <= input(7);
output(0, 239) <= input(8);
output(0, 240) <= input(45);
output(0, 241) <= input(43);
output(0, 242) <= input(41);
output(0, 243) <= input(39);
output(0, 244) <= input(37);
output(0, 245) <= input(35);
output(0, 246) <= input(33);
output(0, 247) <= input(16);
output(0, 248) <= input(17);
output(0, 249) <= input(18);
output(0, 250) <= input(19);
output(0, 251) <= input(20);
output(0, 252) <= input(21);
output(0, 253) <= input(22);
output(0, 254) <= input(23);
output(0, 255) <= input(24);
output(1, 0) <= input(16);
output(1, 1) <= input(17);
output(1, 2) <= input(18);
output(1, 3) <= input(19);
output(1, 4) <= input(20);
output(1, 5) <= input(21);
output(1, 6) <= input(22);
output(1, 7) <= input(23);
output(1, 8) <= input(24);
output(1, 9) <= input(25);
output(1, 10) <= input(26);
output(1, 11) <= input(27);
output(1, 12) <= input(28);
output(1, 13) <= input(29);
output(1, 14) <= input(30);
output(1, 15) <= input(31);
output(1, 16) <= input(32);
output(1, 17) <= input(0);
output(1, 18) <= input(1);
output(1, 19) <= input(2);
output(1, 20) <= input(3);
output(1, 21) <= input(4);
output(1, 22) <= input(5);
output(1, 23) <= input(6);
output(1, 24) <= input(7);
output(1, 25) <= input(8);
output(1, 26) <= input(9);
output(1, 27) <= input(10);
output(1, 28) <= input(11);
output(1, 29) <= input(12);
output(1, 30) <= input(13);
output(1, 31) <= input(14);
output(1, 32) <= input(33);
output(1, 33) <= input(16);
output(1, 34) <= input(17);
output(1, 35) <= input(18);
output(1, 36) <= input(19);
output(1, 37) <= input(20);
output(1, 38) <= input(21);
output(1, 39) <= input(22);
output(1, 40) <= input(23);
output(1, 41) <= input(24);
output(1, 42) <= input(25);
output(1, 43) <= input(26);
output(1, 44) <= input(27);
output(1, 45) <= input(28);
output(1, 46) <= input(29);
output(1, 47) <= input(30);
output(1, 48) <= input(46);
output(1, 49) <= input(32);
output(1, 50) <= input(0);
output(1, 51) <= input(1);
output(1, 52) <= input(2);
output(1, 53) <= input(3);
output(1, 54) <= input(4);
output(1, 55) <= input(5);
output(1, 56) <= input(6);
output(1, 57) <= input(7);
output(1, 58) <= input(8);
output(1, 59) <= input(9);
output(1, 60) <= input(10);
output(1, 61) <= input(11);
output(1, 62) <= input(12);
output(1, 63) <= input(13);
output(1, 64) <= input(47);
output(1, 65) <= input(33);
output(1, 66) <= input(16);
output(1, 67) <= input(17);
output(1, 68) <= input(18);
output(1, 69) <= input(19);
output(1, 70) <= input(20);
output(1, 71) <= input(21);
output(1, 72) <= input(22);
output(1, 73) <= input(23);
output(1, 74) <= input(24);
output(1, 75) <= input(25);
output(1, 76) <= input(26);
output(1, 77) <= input(27);
output(1, 78) <= input(28);
output(1, 79) <= input(29);
output(1, 80) <= input(48);
output(1, 81) <= input(46);
output(1, 82) <= input(32);
output(1, 83) <= input(0);
output(1, 84) <= input(1);
output(1, 85) <= input(2);
output(1, 86) <= input(3);
output(1, 87) <= input(4);
output(1, 88) <= input(5);
output(1, 89) <= input(6);
output(1, 90) <= input(7);
output(1, 91) <= input(8);
output(1, 92) <= input(9);
output(1, 93) <= input(10);
output(1, 94) <= input(11);
output(1, 95) <= input(12);
output(1, 96) <= input(49);
output(1, 97) <= input(47);
output(1, 98) <= input(33);
output(1, 99) <= input(16);
output(1, 100) <= input(17);
output(1, 101) <= input(18);
output(1, 102) <= input(19);
output(1, 103) <= input(20);
output(1, 104) <= input(21);
output(1, 105) <= input(22);
output(1, 106) <= input(23);
output(1, 107) <= input(24);
output(1, 108) <= input(25);
output(1, 109) <= input(26);
output(1, 110) <= input(27);
output(1, 111) <= input(28);
output(1, 112) <= input(50);
output(1, 113) <= input(48);
output(1, 114) <= input(46);
output(1, 115) <= input(32);
output(1, 116) <= input(0);
output(1, 117) <= input(1);
output(1, 118) <= input(2);
output(1, 119) <= input(3);
output(1, 120) <= input(4);
output(1, 121) <= input(5);
output(1, 122) <= input(6);
output(1, 123) <= input(7);
output(1, 124) <= input(8);
output(1, 125) <= input(9);
output(1, 126) <= input(10);
output(1, 127) <= input(11);
output(1, 128) <= input(51);
output(1, 129) <= input(50);
output(1, 130) <= input(48);
output(1, 131) <= input(46);
output(1, 132) <= input(32);
output(1, 133) <= input(0);
output(1, 134) <= input(1);
output(1, 135) <= input(2);
output(1, 136) <= input(3);
output(1, 137) <= input(4);
output(1, 138) <= input(5);
output(1, 139) <= input(6);
output(1, 140) <= input(7);
output(1, 141) <= input(8);
output(1, 142) <= input(9);
output(1, 143) <= input(10);
output(1, 144) <= input(52);
output(1, 145) <= input(53);
output(1, 146) <= input(49);
output(1, 147) <= input(47);
output(1, 148) <= input(33);
output(1, 149) <= input(16);
output(1, 150) <= input(17);
output(1, 151) <= input(18);
output(1, 152) <= input(19);
output(1, 153) <= input(20);
output(1, 154) <= input(21);
output(1, 155) <= input(22);
output(1, 156) <= input(23);
output(1, 157) <= input(24);
output(1, 158) <= input(25);
output(1, 159) <= input(26);
output(1, 160) <= input(54);
output(1, 161) <= input(51);
output(1, 162) <= input(50);
output(1, 163) <= input(48);
output(1, 164) <= input(46);
output(1, 165) <= input(32);
output(1, 166) <= input(0);
output(1, 167) <= input(1);
output(1, 168) <= input(2);
output(1, 169) <= input(3);
output(1, 170) <= input(4);
output(1, 171) <= input(5);
output(1, 172) <= input(6);
output(1, 173) <= input(7);
output(1, 174) <= input(8);
output(1, 175) <= input(9);
output(1, 176) <= input(55);
output(1, 177) <= input(52);
output(1, 178) <= input(53);
output(1, 179) <= input(49);
output(1, 180) <= input(47);
output(1, 181) <= input(33);
output(1, 182) <= input(16);
output(1, 183) <= input(17);
output(1, 184) <= input(18);
output(1, 185) <= input(19);
output(1, 186) <= input(20);
output(1, 187) <= input(21);
output(1, 188) <= input(22);
output(1, 189) <= input(23);
output(1, 190) <= input(24);
output(1, 191) <= input(25);
output(1, 192) <= input(56);
output(1, 193) <= input(54);
output(1, 194) <= input(51);
output(1, 195) <= input(50);
output(1, 196) <= input(48);
output(1, 197) <= input(46);
output(1, 198) <= input(32);
output(1, 199) <= input(0);
output(1, 200) <= input(1);
output(1, 201) <= input(2);
output(1, 202) <= input(3);
output(1, 203) <= input(4);
output(1, 204) <= input(5);
output(1, 205) <= input(6);
output(1, 206) <= input(7);
output(1, 207) <= input(8);
output(1, 208) <= input(57);
output(1, 209) <= input(55);
output(1, 210) <= input(52);
output(1, 211) <= input(53);
output(1, 212) <= input(49);
output(1, 213) <= input(47);
output(1, 214) <= input(33);
output(1, 215) <= input(16);
output(1, 216) <= input(17);
output(1, 217) <= input(18);
output(1, 218) <= input(19);
output(1, 219) <= input(20);
output(1, 220) <= input(21);
output(1, 221) <= input(22);
output(1, 222) <= input(23);
output(1, 223) <= input(24);
output(1, 224) <= input(58);
output(1, 225) <= input(56);
output(1, 226) <= input(54);
output(1, 227) <= input(51);
output(1, 228) <= input(50);
output(1, 229) <= input(48);
output(1, 230) <= input(46);
output(1, 231) <= input(32);
output(1, 232) <= input(0);
output(1, 233) <= input(1);
output(1, 234) <= input(2);
output(1, 235) <= input(3);
output(1, 236) <= input(4);
output(1, 237) <= input(5);
output(1, 238) <= input(6);
output(1, 239) <= input(7);
output(1, 240) <= input(59);
output(1, 241) <= input(57);
output(1, 242) <= input(55);
output(1, 243) <= input(52);
output(1, 244) <= input(53);
output(1, 245) <= input(49);
output(1, 246) <= input(47);
output(1, 247) <= input(33);
output(1, 248) <= input(16);
output(1, 249) <= input(17);
output(1, 250) <= input(18);
output(1, 251) <= input(19);
output(1, 252) <= input(20);
output(1, 253) <= input(21);
output(1, 254) <= input(22);
output(1, 255) <= input(23);
when "0110" =>
output(0, 0) <= input(0);
output(0, 1) <= input(1);
output(0, 2) <= input(2);
output(0, 3) <= input(3);
output(0, 4) <= input(4);
output(0, 5) <= input(5);
output(0, 6) <= input(6);
output(0, 7) <= input(7);
output(0, 8) <= input(8);
output(0, 9) <= input(9);
output(0, 10) <= input(10);
output(0, 11) <= input(11);
output(0, 12) <= input(12);
output(0, 13) <= input(13);
output(0, 14) <= input(14);
output(0, 15) <= input(15);
output(0, 16) <= input(16);
output(0, 17) <= input(17);
output(0, 18) <= input(18);
output(0, 19) <= input(19);
output(0, 20) <= input(20);
output(0, 21) <= input(21);
output(0, 22) <= input(22);
output(0, 23) <= input(23);
output(0, 24) <= input(24);
output(0, 25) <= input(25);
output(0, 26) <= input(26);
output(0, 27) <= input(27);
output(0, 28) <= input(28);
output(0, 29) <= input(29);
output(0, 30) <= input(30);
output(0, 31) <= input(31);
output(0, 32) <= input(32);
output(0, 33) <= input(0);
output(0, 34) <= input(1);
output(0, 35) <= input(2);
output(0, 36) <= input(3);
output(0, 37) <= input(4);
output(0, 38) <= input(5);
output(0, 39) <= input(6);
output(0, 40) <= input(7);
output(0, 41) <= input(8);
output(0, 42) <= input(9);
output(0, 43) <= input(10);
output(0, 44) <= input(11);
output(0, 45) <= input(12);
output(0, 46) <= input(13);
output(0, 47) <= input(14);
output(0, 48) <= input(33);
output(0, 49) <= input(16);
output(0, 50) <= input(17);
output(0, 51) <= input(18);
output(0, 52) <= input(19);
output(0, 53) <= input(20);
output(0, 54) <= input(21);
output(0, 55) <= input(22);
output(0, 56) <= input(23);
output(0, 57) <= input(24);
output(0, 58) <= input(25);
output(0, 59) <= input(26);
output(0, 60) <= input(27);
output(0, 61) <= input(28);
output(0, 62) <= input(29);
output(0, 63) <= input(30);
output(0, 64) <= input(34);
output(0, 65) <= input(33);
output(0, 66) <= input(16);
output(0, 67) <= input(17);
output(0, 68) <= input(18);
output(0, 69) <= input(19);
output(0, 70) <= input(20);
output(0, 71) <= input(21);
output(0, 72) <= input(22);
output(0, 73) <= input(23);
output(0, 74) <= input(24);
output(0, 75) <= input(25);
output(0, 76) <= input(26);
output(0, 77) <= input(27);
output(0, 78) <= input(28);
output(0, 79) <= input(29);
output(0, 80) <= input(35);
output(0, 81) <= input(36);
output(0, 82) <= input(32);
output(0, 83) <= input(0);
output(0, 84) <= input(1);
output(0, 85) <= input(2);
output(0, 86) <= input(3);
output(0, 87) <= input(4);
output(0, 88) <= input(5);
output(0, 89) <= input(6);
output(0, 90) <= input(7);
output(0, 91) <= input(8);
output(0, 92) <= input(9);
output(0, 93) <= input(10);
output(0, 94) <= input(11);
output(0, 95) <= input(12);
output(0, 96) <= input(37);
output(0, 97) <= input(34);
output(0, 98) <= input(33);
output(0, 99) <= input(16);
output(0, 100) <= input(17);
output(0, 101) <= input(18);
output(0, 102) <= input(19);
output(0, 103) <= input(20);
output(0, 104) <= input(21);
output(0, 105) <= input(22);
output(0, 106) <= input(23);
output(0, 107) <= input(24);
output(0, 108) <= input(25);
output(0, 109) <= input(26);
output(0, 110) <= input(27);
output(0, 111) <= input(28);
output(0, 112) <= input(38);
output(0, 113) <= input(35);
output(0, 114) <= input(36);
output(0, 115) <= input(32);
output(0, 116) <= input(0);
output(0, 117) <= input(1);
output(0, 118) <= input(2);
output(0, 119) <= input(3);
output(0, 120) <= input(4);
output(0, 121) <= input(5);
output(0, 122) <= input(6);
output(0, 123) <= input(7);
output(0, 124) <= input(8);
output(0, 125) <= input(9);
output(0, 126) <= input(10);
output(0, 127) <= input(11);
output(0, 128) <= input(39);
output(0, 129) <= input(38);
output(0, 130) <= input(35);
output(0, 131) <= input(36);
output(0, 132) <= input(32);
output(0, 133) <= input(0);
output(0, 134) <= input(1);
output(0, 135) <= input(2);
output(0, 136) <= input(3);
output(0, 137) <= input(4);
output(0, 138) <= input(5);
output(0, 139) <= input(6);
output(0, 140) <= input(7);
output(0, 141) <= input(8);
output(0, 142) <= input(9);
output(0, 143) <= input(10);
output(0, 144) <= input(40);
output(0, 145) <= input(41);
output(0, 146) <= input(37);
output(0, 147) <= input(34);
output(0, 148) <= input(33);
output(0, 149) <= input(16);
output(0, 150) <= input(17);
output(0, 151) <= input(18);
output(0, 152) <= input(19);
output(0, 153) <= input(20);
output(0, 154) <= input(21);
output(0, 155) <= input(22);
output(0, 156) <= input(23);
output(0, 157) <= input(24);
output(0, 158) <= input(25);
output(0, 159) <= input(26);
output(0, 160) <= input(42);
output(0, 161) <= input(39);
output(0, 162) <= input(38);
output(0, 163) <= input(35);
output(0, 164) <= input(36);
output(0, 165) <= input(32);
output(0, 166) <= input(0);
output(0, 167) <= input(1);
output(0, 168) <= input(2);
output(0, 169) <= input(3);
output(0, 170) <= input(4);
output(0, 171) <= input(5);
output(0, 172) <= input(6);
output(0, 173) <= input(7);
output(0, 174) <= input(8);
output(0, 175) <= input(9);
output(0, 176) <= input(43);
output(0, 177) <= input(40);
output(0, 178) <= input(41);
output(0, 179) <= input(37);
output(0, 180) <= input(34);
output(0, 181) <= input(33);
output(0, 182) <= input(16);
output(0, 183) <= input(17);
output(0, 184) <= input(18);
output(0, 185) <= input(19);
output(0, 186) <= input(20);
output(0, 187) <= input(21);
output(0, 188) <= input(22);
output(0, 189) <= input(23);
output(0, 190) <= input(24);
output(0, 191) <= input(25);
output(0, 192) <= input(44);
output(0, 193) <= input(43);
output(0, 194) <= input(40);
output(0, 195) <= input(41);
output(0, 196) <= input(37);
output(0, 197) <= input(34);
output(0, 198) <= input(33);
output(0, 199) <= input(16);
output(0, 200) <= input(17);
output(0, 201) <= input(18);
output(0, 202) <= input(19);
output(0, 203) <= input(20);
output(0, 204) <= input(21);
output(0, 205) <= input(22);
output(0, 206) <= input(23);
output(0, 207) <= input(24);
output(0, 208) <= input(45);
output(0, 209) <= input(46);
output(0, 210) <= input(42);
output(0, 211) <= input(39);
output(0, 212) <= input(38);
output(0, 213) <= input(35);
output(0, 214) <= input(36);
output(0, 215) <= input(32);
output(0, 216) <= input(0);
output(0, 217) <= input(1);
output(0, 218) <= input(2);
output(0, 219) <= input(3);
output(0, 220) <= input(4);
output(0, 221) <= input(5);
output(0, 222) <= input(6);
output(0, 223) <= input(7);
output(0, 224) <= input(47);
output(0, 225) <= input(44);
output(0, 226) <= input(43);
output(0, 227) <= input(40);
output(0, 228) <= input(41);
output(0, 229) <= input(37);
output(0, 230) <= input(34);
output(0, 231) <= input(33);
output(0, 232) <= input(16);
output(0, 233) <= input(17);
output(0, 234) <= input(18);
output(0, 235) <= input(19);
output(0, 236) <= input(20);
output(0, 237) <= input(21);
output(0, 238) <= input(22);
output(0, 239) <= input(23);
output(0, 240) <= input(48);
output(0, 241) <= input(45);
output(0, 242) <= input(46);
output(0, 243) <= input(42);
output(0, 244) <= input(39);
output(0, 245) <= input(38);
output(0, 246) <= input(35);
output(0, 247) <= input(36);
output(0, 248) <= input(32);
output(0, 249) <= input(0);
output(0, 250) <= input(1);
output(0, 251) <= input(2);
output(0, 252) <= input(3);
output(0, 253) <= input(4);
output(0, 254) <= input(5);
output(0, 255) <= input(6);
output(1, 0) <= input(49);
output(1, 1) <= input(1);
output(1, 2) <= input(2);
output(1, 3) <= input(3);
output(1, 4) <= input(4);
output(1, 5) <= input(5);
output(1, 6) <= input(6);
output(1, 7) <= input(7);
output(1, 8) <= input(8);
output(1, 9) <= input(9);
output(1, 10) <= input(10);
output(1, 11) <= input(11);
output(1, 12) <= input(12);
output(1, 13) <= input(13);
output(1, 14) <= input(14);
output(1, 15) <= input(15);
output(1, 16) <= input(50);
output(1, 17) <= input(51);
output(1, 18) <= input(18);
output(1, 19) <= input(19);
output(1, 20) <= input(20);
output(1, 21) <= input(21);
output(1, 22) <= input(22);
output(1, 23) <= input(23);
output(1, 24) <= input(24);
output(1, 25) <= input(25);
output(1, 26) <= input(26);
output(1, 27) <= input(27);
output(1, 28) <= input(28);
output(1, 29) <= input(29);
output(1, 30) <= input(30);
output(1, 31) <= input(31);
output(1, 32) <= input(52);
output(1, 33) <= input(50);
output(1, 34) <= input(51);
output(1, 35) <= input(18);
output(1, 36) <= input(19);
output(1, 37) <= input(20);
output(1, 38) <= input(21);
output(1, 39) <= input(22);
output(1, 40) <= input(23);
output(1, 41) <= input(24);
output(1, 42) <= input(25);
output(1, 43) <= input(26);
output(1, 44) <= input(27);
output(1, 45) <= input(28);
output(1, 46) <= input(29);
output(1, 47) <= input(30);
output(1, 48) <= input(53);
output(1, 49) <= input(54);
output(1, 50) <= input(49);
output(1, 51) <= input(1);
output(1, 52) <= input(2);
output(1, 53) <= input(3);
output(1, 54) <= input(4);
output(1, 55) <= input(5);
output(1, 56) <= input(6);
output(1, 57) <= input(7);
output(1, 58) <= input(8);
output(1, 59) <= input(9);
output(1, 60) <= input(10);
output(1, 61) <= input(11);
output(1, 62) <= input(12);
output(1, 63) <= input(13);
output(1, 64) <= input(55);
output(1, 65) <= input(53);
output(1, 66) <= input(54);
output(1, 67) <= input(49);
output(1, 68) <= input(1);
output(1, 69) <= input(2);
output(1, 70) <= input(3);
output(1, 71) <= input(4);
output(1, 72) <= input(5);
output(1, 73) <= input(6);
output(1, 74) <= input(7);
output(1, 75) <= input(8);
output(1, 76) <= input(9);
output(1, 77) <= input(10);
output(1, 78) <= input(11);
output(1, 79) <= input(12);
output(1, 80) <= input(56);
output(1, 81) <= input(57);
output(1, 82) <= input(52);
output(1, 83) <= input(50);
output(1, 84) <= input(51);
output(1, 85) <= input(18);
output(1, 86) <= input(19);
output(1, 87) <= input(20);
output(1, 88) <= input(21);
output(1, 89) <= input(22);
output(1, 90) <= input(23);
output(1, 91) <= input(24);
output(1, 92) <= input(25);
output(1, 93) <= input(26);
output(1, 94) <= input(27);
output(1, 95) <= input(28);
output(1, 96) <= input(58);
output(1, 97) <= input(56);
output(1, 98) <= input(57);
output(1, 99) <= input(52);
output(1, 100) <= input(50);
output(1, 101) <= input(51);
output(1, 102) <= input(18);
output(1, 103) <= input(19);
output(1, 104) <= input(20);
output(1, 105) <= input(21);
output(1, 106) <= input(22);
output(1, 107) <= input(23);
output(1, 108) <= input(24);
output(1, 109) <= input(25);
output(1, 110) <= input(26);
output(1, 111) <= input(27);
output(1, 112) <= input(59);
output(1, 113) <= input(60);
output(1, 114) <= input(55);
output(1, 115) <= input(53);
output(1, 116) <= input(54);
output(1, 117) <= input(49);
output(1, 118) <= input(1);
output(1, 119) <= input(2);
output(1, 120) <= input(3);
output(1, 121) <= input(4);
output(1, 122) <= input(5);
output(1, 123) <= input(6);
output(1, 124) <= input(7);
output(1, 125) <= input(8);
output(1, 126) <= input(9);
output(1, 127) <= input(10);
output(1, 128) <= input(61);
output(1, 129) <= input(58);
output(1, 130) <= input(56);
output(1, 131) <= input(57);
output(1, 132) <= input(52);
output(1, 133) <= input(50);
output(1, 134) <= input(51);
output(1, 135) <= input(18);
output(1, 136) <= input(19);
output(1, 137) <= input(20);
output(1, 138) <= input(21);
output(1, 139) <= input(22);
output(1, 140) <= input(23);
output(1, 141) <= input(24);
output(1, 142) <= input(25);
output(1, 143) <= input(26);
output(1, 144) <= input(62);
output(1, 145) <= input(61);
output(1, 146) <= input(58);
output(1, 147) <= input(56);
output(1, 148) <= input(57);
output(1, 149) <= input(52);
output(1, 150) <= input(50);
output(1, 151) <= input(51);
output(1, 152) <= input(18);
output(1, 153) <= input(19);
output(1, 154) <= input(20);
output(1, 155) <= input(21);
output(1, 156) <= input(22);
output(1, 157) <= input(23);
output(1, 158) <= input(24);
output(1, 159) <= input(25);
output(1, 160) <= input(63);
output(1, 161) <= input(64);
output(1, 162) <= input(59);
output(1, 163) <= input(60);
output(1, 164) <= input(55);
output(1, 165) <= input(53);
output(1, 166) <= input(54);
output(1, 167) <= input(49);
output(1, 168) <= input(1);
output(1, 169) <= input(2);
output(1, 170) <= input(3);
output(1, 171) <= input(4);
output(1, 172) <= input(5);
output(1, 173) <= input(6);
output(1, 174) <= input(7);
output(1, 175) <= input(8);
output(1, 176) <= input(46);
output(1, 177) <= input(63);
output(1, 178) <= input(64);
output(1, 179) <= input(59);
output(1, 180) <= input(60);
output(1, 181) <= input(55);
output(1, 182) <= input(53);
output(1, 183) <= input(54);
output(1, 184) <= input(49);
output(1, 185) <= input(1);
output(1, 186) <= input(2);
output(1, 187) <= input(3);
output(1, 188) <= input(4);
output(1, 189) <= input(5);
output(1, 190) <= input(6);
output(1, 191) <= input(7);
output(1, 192) <= input(44);
output(1, 193) <= input(43);
output(1, 194) <= input(62);
output(1, 195) <= input(61);
output(1, 196) <= input(58);
output(1, 197) <= input(56);
output(1, 198) <= input(57);
output(1, 199) <= input(52);
output(1, 200) <= input(50);
output(1, 201) <= input(51);
output(1, 202) <= input(18);
output(1, 203) <= input(19);
output(1, 204) <= input(20);
output(1, 205) <= input(21);
output(1, 206) <= input(22);
output(1, 207) <= input(23);
output(1, 208) <= input(65);
output(1, 209) <= input(44);
output(1, 210) <= input(43);
output(1, 211) <= input(62);
output(1, 212) <= input(61);
output(1, 213) <= input(58);
output(1, 214) <= input(56);
output(1, 215) <= input(57);
output(1, 216) <= input(52);
output(1, 217) <= input(50);
output(1, 218) <= input(51);
output(1, 219) <= input(18);
output(1, 220) <= input(19);
output(1, 221) <= input(20);
output(1, 222) <= input(21);
output(1, 223) <= input(22);
output(1, 224) <= input(66);
output(1, 225) <= input(45);
output(1, 226) <= input(46);
output(1, 227) <= input(63);
output(1, 228) <= input(64);
output(1, 229) <= input(59);
output(1, 230) <= input(60);
output(1, 231) <= input(55);
output(1, 232) <= input(53);
output(1, 233) <= input(54);
output(1, 234) <= input(49);
output(1, 235) <= input(1);
output(1, 236) <= input(2);
output(1, 237) <= input(3);
output(1, 238) <= input(4);
output(1, 239) <= input(5);
output(1, 240) <= input(67);
output(1, 241) <= input(65);
output(1, 242) <= input(44);
output(1, 243) <= input(43);
output(1, 244) <= input(62);
output(1, 245) <= input(61);
output(1, 246) <= input(58);
output(1, 247) <= input(56);
output(1, 248) <= input(57);
output(1, 249) <= input(52);
output(1, 250) <= input(50);
output(1, 251) <= input(51);
output(1, 252) <= input(18);
output(1, 253) <= input(19);
output(1, 254) <= input(20);
output(1, 255) <= input(21);
output(2, 0) <= input(49);
output(2, 1) <= input(1);
output(2, 2) <= input(2);
output(2, 3) <= input(3);
output(2, 4) <= input(4);
output(2, 5) <= input(5);
output(2, 6) <= input(6);
output(2, 7) <= input(7);
output(2, 8) <= input(8);
output(2, 9) <= input(9);
output(2, 10) <= input(10);
output(2, 11) <= input(11);
output(2, 12) <= input(12);
output(2, 13) <= input(13);
output(2, 14) <= input(14);
output(2, 15) <= input(15);
output(2, 16) <= input(68);
output(2, 17) <= input(49);
output(2, 18) <= input(1);
output(2, 19) <= input(2);
output(2, 20) <= input(3);
output(2, 21) <= input(4);
output(2, 22) <= input(5);
output(2, 23) <= input(6);
output(2, 24) <= input(7);
output(2, 25) <= input(8);
output(2, 26) <= input(9);
output(2, 27) <= input(10);
output(2, 28) <= input(11);
output(2, 29) <= input(12);
output(2, 30) <= input(13);
output(2, 31) <= input(14);
output(2, 32) <= input(69);
output(2, 33) <= input(70);
output(2, 34) <= input(51);
output(2, 35) <= input(18);
output(2, 36) <= input(19);
output(2, 37) <= input(20);
output(2, 38) <= input(21);
output(2, 39) <= input(22);
output(2, 40) <= input(23);
output(2, 41) <= input(24);
output(2, 42) <= input(25);
output(2, 43) <= input(26);
output(2, 44) <= input(27);
output(2, 45) <= input(28);
output(2, 46) <= input(29);
output(2, 47) <= input(30);
output(2, 48) <= input(71);
output(2, 49) <= input(69);
output(2, 50) <= input(70);
output(2, 51) <= input(51);
output(2, 52) <= input(18);
output(2, 53) <= input(19);
output(2, 54) <= input(20);
output(2, 55) <= input(21);
output(2, 56) <= input(22);
output(2, 57) <= input(23);
output(2, 58) <= input(24);
output(2, 59) <= input(25);
output(2, 60) <= input(26);
output(2, 61) <= input(27);
output(2, 62) <= input(28);
output(2, 63) <= input(29);
output(2, 64) <= input(72);
output(2, 65) <= input(71);
output(2, 66) <= input(69);
output(2, 67) <= input(70);
output(2, 68) <= input(51);
output(2, 69) <= input(18);
output(2, 70) <= input(19);
output(2, 71) <= input(20);
output(2, 72) <= input(21);
output(2, 73) <= input(22);
output(2, 74) <= input(23);
output(2, 75) <= input(24);
output(2, 76) <= input(25);
output(2, 77) <= input(26);
output(2, 78) <= input(27);
output(2, 79) <= input(28);
output(2, 80) <= input(73);
output(2, 81) <= input(74);
output(2, 82) <= input(75);
output(2, 83) <= input(68);
output(2, 84) <= input(49);
output(2, 85) <= input(1);
output(2, 86) <= input(2);
output(2, 87) <= input(3);
output(2, 88) <= input(4);
output(2, 89) <= input(5);
output(2, 90) <= input(6);
output(2, 91) <= input(7);
output(2, 92) <= input(8);
output(2, 93) <= input(9);
output(2, 94) <= input(10);
output(2, 95) <= input(11);
output(2, 96) <= input(76);
output(2, 97) <= input(73);
output(2, 98) <= input(74);
output(2, 99) <= input(75);
output(2, 100) <= input(68);
output(2, 101) <= input(49);
output(2, 102) <= input(1);
output(2, 103) <= input(2);
output(2, 104) <= input(3);
output(2, 105) <= input(4);
output(2, 106) <= input(5);
output(2, 107) <= input(6);
output(2, 108) <= input(7);
output(2, 109) <= input(8);
output(2, 110) <= input(9);
output(2, 111) <= input(10);
output(2, 112) <= input(77);
output(2, 113) <= input(78);
output(2, 114) <= input(72);
output(2, 115) <= input(71);
output(2, 116) <= input(69);
output(2, 117) <= input(70);
output(2, 118) <= input(51);
output(2, 119) <= input(18);
output(2, 120) <= input(19);
output(2, 121) <= input(20);
output(2, 122) <= input(21);
output(2, 123) <= input(22);
output(2, 124) <= input(23);
output(2, 125) <= input(24);
output(2, 126) <= input(25);
output(2, 127) <= input(26);
output(2, 128) <= input(79);
output(2, 129) <= input(77);
output(2, 130) <= input(78);
output(2, 131) <= input(72);
output(2, 132) <= input(71);
output(2, 133) <= input(69);
output(2, 134) <= input(70);
output(2, 135) <= input(51);
output(2, 136) <= input(18);
output(2, 137) <= input(19);
output(2, 138) <= input(20);
output(2, 139) <= input(21);
output(2, 140) <= input(22);
output(2, 141) <= input(23);
output(2, 142) <= input(24);
output(2, 143) <= input(25);
output(2, 144) <= input(80);
output(2, 145) <= input(79);
output(2, 146) <= input(77);
output(2, 147) <= input(78);
output(2, 148) <= input(72);
output(2, 149) <= input(71);
output(2, 150) <= input(69);
output(2, 151) <= input(70);
output(2, 152) <= input(51);
output(2, 153) <= input(18);
output(2, 154) <= input(19);
output(2, 155) <= input(20);
output(2, 156) <= input(21);
output(2, 157) <= input(22);
output(2, 158) <= input(23);
output(2, 159) <= input(24);
output(2, 160) <= input(81);
output(2, 161) <= input(82);
output(2, 162) <= input(83);
output(2, 163) <= input(76);
output(2, 164) <= input(73);
output(2, 165) <= input(74);
output(2, 166) <= input(75);
output(2, 167) <= input(68);
output(2, 168) <= input(49);
output(2, 169) <= input(1);
output(2, 170) <= input(2);
output(2, 171) <= input(3);
output(2, 172) <= input(4);
output(2, 173) <= input(5);
output(2, 174) <= input(6);
output(2, 175) <= input(7);
output(2, 176) <= input(84);
output(2, 177) <= input(81);
output(2, 178) <= input(82);
output(2, 179) <= input(83);
output(2, 180) <= input(76);
output(2, 181) <= input(73);
output(2, 182) <= input(74);
output(2, 183) <= input(75);
output(2, 184) <= input(68);
output(2, 185) <= input(49);
output(2, 186) <= input(1);
output(2, 187) <= input(2);
output(2, 188) <= input(3);
output(2, 189) <= input(4);
output(2, 190) <= input(5);
output(2, 191) <= input(6);
output(2, 192) <= input(85);
output(2, 193) <= input(84);
output(2, 194) <= input(81);
output(2, 195) <= input(82);
output(2, 196) <= input(83);
output(2, 197) <= input(76);
output(2, 198) <= input(73);
output(2, 199) <= input(74);
output(2, 200) <= input(75);
output(2, 201) <= input(68);
output(2, 202) <= input(49);
output(2, 203) <= input(1);
output(2, 204) <= input(2);
output(2, 205) <= input(3);
output(2, 206) <= input(4);
output(2, 207) <= input(5);
output(2, 208) <= input(86);
output(2, 209) <= input(87);
output(2, 210) <= input(88);
output(2, 211) <= input(80);
output(2, 212) <= input(79);
output(2, 213) <= input(77);
output(2, 214) <= input(78);
output(2, 215) <= input(72);
output(2, 216) <= input(71);
output(2, 217) <= input(69);
output(2, 218) <= input(70);
output(2, 219) <= input(51);
output(2, 220) <= input(18);
output(2, 221) <= input(19);
output(2, 222) <= input(20);
output(2, 223) <= input(21);
output(2, 224) <= input(89);
output(2, 225) <= input(86);
output(2, 226) <= input(87);
output(2, 227) <= input(88);
output(2, 228) <= input(80);
output(2, 229) <= input(79);
output(2, 230) <= input(77);
output(2, 231) <= input(78);
output(2, 232) <= input(72);
output(2, 233) <= input(71);
output(2, 234) <= input(69);
output(2, 235) <= input(70);
output(2, 236) <= input(51);
output(2, 237) <= input(18);
output(2, 238) <= input(19);
output(2, 239) <= input(20);
output(2, 240) <= input(90);
output(2, 241) <= input(91);
output(2, 242) <= input(85);
output(2, 243) <= input(84);
output(2, 244) <= input(81);
output(2, 245) <= input(82);
output(2, 246) <= input(83);
output(2, 247) <= input(76);
output(2, 248) <= input(73);
output(2, 249) <= input(74);
output(2, 250) <= input(75);
output(2, 251) <= input(68);
output(2, 252) <= input(49);
output(2, 253) <= input(1);
output(2, 254) <= input(2);
output(2, 255) <= input(3);
when "0111" =>
output(0, 0) <= input(0);
output(0, 1) <= input(1);
output(0, 2) <= input(2);
output(0, 3) <= input(3);
output(0, 4) <= input(4);
output(0, 5) <= input(5);
output(0, 6) <= input(6);
output(0, 7) <= input(7);
output(0, 8) <= input(8);
output(0, 9) <= input(9);
output(0, 10) <= input(10);
output(0, 11) <= input(11);
output(0, 12) <= input(12);
output(0, 13) <= input(13);
output(0, 14) <= input(14);
output(0, 15) <= input(15);
output(0, 16) <= input(16);
output(0, 17) <= input(0);
output(0, 18) <= input(1);
output(0, 19) <= input(2);
output(0, 20) <= input(3);
output(0, 21) <= input(4);
output(0, 22) <= input(5);
output(0, 23) <= input(6);
output(0, 24) <= input(7);
output(0, 25) <= input(8);
output(0, 26) <= input(9);
output(0, 27) <= input(10);
output(0, 28) <= input(11);
output(0, 29) <= input(12);
output(0, 30) <= input(13);
output(0, 31) <= input(14);
output(0, 32) <= input(17);
output(0, 33) <= input(16);
output(0, 34) <= input(0);
output(0, 35) <= input(1);
output(0, 36) <= input(2);
output(0, 37) <= input(3);
output(0, 38) <= input(4);
output(0, 39) <= input(5);
output(0, 40) <= input(6);
output(0, 41) <= input(7);
output(0, 42) <= input(8);
output(0, 43) <= input(9);
output(0, 44) <= input(10);
output(0, 45) <= input(11);
output(0, 46) <= input(12);
output(0, 47) <= input(13);
output(0, 48) <= input(18);
output(0, 49) <= input(17);
output(0, 50) <= input(16);
output(0, 51) <= input(0);
output(0, 52) <= input(1);
output(0, 53) <= input(2);
output(0, 54) <= input(3);
output(0, 55) <= input(4);
output(0, 56) <= input(5);
output(0, 57) <= input(6);
output(0, 58) <= input(7);
output(0, 59) <= input(8);
output(0, 60) <= input(9);
output(0, 61) <= input(10);
output(0, 62) <= input(11);
output(0, 63) <= input(12);
output(0, 64) <= input(19);
output(0, 65) <= input(18);
output(0, 66) <= input(17);
output(0, 67) <= input(16);
output(0, 68) <= input(0);
output(0, 69) <= input(1);
output(0, 70) <= input(2);
output(0, 71) <= input(3);
output(0, 72) <= input(4);
output(0, 73) <= input(5);
output(0, 74) <= input(6);
output(0, 75) <= input(7);
output(0, 76) <= input(8);
output(0, 77) <= input(9);
output(0, 78) <= input(10);
output(0, 79) <= input(11);
output(0, 80) <= input(20);
output(0, 81) <= input(21);
output(0, 82) <= input(22);
output(0, 83) <= input(23);
output(0, 84) <= input(24);
output(0, 85) <= input(25);
output(0, 86) <= input(26);
output(0, 87) <= input(27);
output(0, 88) <= input(28);
output(0, 89) <= input(29);
output(0, 90) <= input(30);
output(0, 91) <= input(31);
output(0, 92) <= input(32);
output(0, 93) <= input(33);
output(0, 94) <= input(34);
output(0, 95) <= input(35);
output(0, 96) <= input(36);
output(0, 97) <= input(20);
output(0, 98) <= input(21);
output(0, 99) <= input(22);
output(0, 100) <= input(23);
output(0, 101) <= input(24);
output(0, 102) <= input(25);
output(0, 103) <= input(26);
output(0, 104) <= input(27);
output(0, 105) <= input(28);
output(0, 106) <= input(29);
output(0, 107) <= input(30);
output(0, 108) <= input(31);
output(0, 109) <= input(32);
output(0, 110) <= input(33);
output(0, 111) <= input(34);
output(0, 112) <= input(37);
output(0, 113) <= input(36);
output(0, 114) <= input(20);
output(0, 115) <= input(21);
output(0, 116) <= input(22);
output(0, 117) <= input(23);
output(0, 118) <= input(24);
output(0, 119) <= input(25);
output(0, 120) <= input(26);
output(0, 121) <= input(27);
output(0, 122) <= input(28);
output(0, 123) <= input(29);
output(0, 124) <= input(30);
output(0, 125) <= input(31);
output(0, 126) <= input(32);
output(0, 127) <= input(33);
output(0, 128) <= input(38);
output(0, 129) <= input(37);
output(0, 130) <= input(36);
output(0, 131) <= input(20);
output(0, 132) <= input(21);
output(0, 133) <= input(22);
output(0, 134) <= input(23);
output(0, 135) <= input(24);
output(0, 136) <= input(25);
output(0, 137) <= input(26);
output(0, 138) <= input(27);
output(0, 139) <= input(28);
output(0, 140) <= input(29);
output(0, 141) <= input(30);
output(0, 142) <= input(31);
output(0, 143) <= input(32);
output(0, 144) <= input(39);
output(0, 145) <= input(38);
output(0, 146) <= input(37);
output(0, 147) <= input(36);
output(0, 148) <= input(20);
output(0, 149) <= input(21);
output(0, 150) <= input(22);
output(0, 151) <= input(23);
output(0, 152) <= input(24);
output(0, 153) <= input(25);
output(0, 154) <= input(26);
output(0, 155) <= input(27);
output(0, 156) <= input(28);
output(0, 157) <= input(29);
output(0, 158) <= input(30);
output(0, 159) <= input(31);
output(0, 160) <= input(40);
output(0, 161) <= input(41);
output(0, 162) <= input(42);
output(0, 163) <= input(43);
output(0, 164) <= input(44);
output(0, 165) <= input(19);
output(0, 166) <= input(18);
output(0, 167) <= input(17);
output(0, 168) <= input(16);
output(0, 169) <= input(0);
output(0, 170) <= input(1);
output(0, 171) <= input(2);
output(0, 172) <= input(3);
output(0, 173) <= input(4);
output(0, 174) <= input(5);
output(0, 175) <= input(6);
output(0, 176) <= input(45);
output(0, 177) <= input(40);
output(0, 178) <= input(41);
output(0, 179) <= input(42);
output(0, 180) <= input(43);
output(0, 181) <= input(44);
output(0, 182) <= input(19);
output(0, 183) <= input(18);
output(0, 184) <= input(17);
output(0, 185) <= input(16);
output(0, 186) <= input(0);
output(0, 187) <= input(1);
output(0, 188) <= input(2);
output(0, 189) <= input(3);
output(0, 190) <= input(4);
output(0, 191) <= input(5);
output(0, 192) <= input(46);
output(0, 193) <= input(45);
output(0, 194) <= input(40);
output(0, 195) <= input(41);
output(0, 196) <= input(42);
output(0, 197) <= input(43);
output(0, 198) <= input(44);
output(0, 199) <= input(19);
output(0, 200) <= input(18);
output(0, 201) <= input(17);
output(0, 202) <= input(16);
output(0, 203) <= input(0);
output(0, 204) <= input(1);
output(0, 205) <= input(2);
output(0, 206) <= input(3);
output(0, 207) <= input(4);
output(0, 208) <= input(47);
output(0, 209) <= input(46);
output(0, 210) <= input(45);
output(0, 211) <= input(40);
output(0, 212) <= input(41);
output(0, 213) <= input(42);
output(0, 214) <= input(43);
output(0, 215) <= input(44);
output(0, 216) <= input(19);
output(0, 217) <= input(18);
output(0, 218) <= input(17);
output(0, 219) <= input(16);
output(0, 220) <= input(0);
output(0, 221) <= input(1);
output(0, 222) <= input(2);
output(0, 223) <= input(3);
output(0, 224) <= input(48);
output(0, 225) <= input(47);
output(0, 226) <= input(46);
output(0, 227) <= input(45);
output(0, 228) <= input(40);
output(0, 229) <= input(41);
output(0, 230) <= input(42);
output(0, 231) <= input(43);
output(0, 232) <= input(44);
output(0, 233) <= input(19);
output(0, 234) <= input(18);
output(0, 235) <= input(17);
output(0, 236) <= input(16);
output(0, 237) <= input(0);
output(0, 238) <= input(1);
output(0, 239) <= input(2);
output(0, 240) <= input(49);
output(0, 241) <= input(50);
output(0, 242) <= input(51);
output(0, 243) <= input(52);
output(0, 244) <= input(53);
output(0, 245) <= input(39);
output(0, 246) <= input(38);
output(0, 247) <= input(37);
output(0, 248) <= input(36);
output(0, 249) <= input(20);
output(0, 250) <= input(21);
output(0, 251) <= input(22);
output(0, 252) <= input(23);
output(0, 253) <= input(24);
output(0, 254) <= input(25);
output(0, 255) <= input(26);
output(1, 0) <= input(54);
output(1, 1) <= input(55);
output(1, 2) <= input(56);
output(1, 3) <= input(57);
output(1, 4) <= input(58);
output(1, 5) <= input(59);
output(1, 6) <= input(60);
output(1, 7) <= input(61);
output(1, 8) <= input(62);
output(1, 9) <= input(63);
output(1, 10) <= input(64);
output(1, 11) <= input(65);
output(1, 12) <= input(66);
output(1, 13) <= input(67);
output(1, 14) <= input(68);
output(1, 15) <= input(69);
output(1, 16) <= input(70);
output(1, 17) <= input(54);
output(1, 18) <= input(55);
output(1, 19) <= input(56);
output(1, 20) <= input(57);
output(1, 21) <= input(58);
output(1, 22) <= input(59);
output(1, 23) <= input(60);
output(1, 24) <= input(61);
output(1, 25) <= input(62);
output(1, 26) <= input(63);
output(1, 27) <= input(64);
output(1, 28) <= input(65);
output(1, 29) <= input(66);
output(1, 30) <= input(67);
output(1, 31) <= input(68);
output(1, 32) <= input(71);
output(1, 33) <= input(70);
output(1, 34) <= input(54);
output(1, 35) <= input(55);
output(1, 36) <= input(56);
output(1, 37) <= input(57);
output(1, 38) <= input(58);
output(1, 39) <= input(59);
output(1, 40) <= input(60);
output(1, 41) <= input(61);
output(1, 42) <= input(62);
output(1, 43) <= input(63);
output(1, 44) <= input(64);
output(1, 45) <= input(65);
output(1, 46) <= input(66);
output(1, 47) <= input(67);
output(1, 48) <= input(72);
output(1, 49) <= input(71);
output(1, 50) <= input(70);
output(1, 51) <= input(54);
output(1, 52) <= input(55);
output(1, 53) <= input(56);
output(1, 54) <= input(57);
output(1, 55) <= input(58);
output(1, 56) <= input(59);
output(1, 57) <= input(60);
output(1, 58) <= input(61);
output(1, 59) <= input(62);
output(1, 60) <= input(63);
output(1, 61) <= input(64);
output(1, 62) <= input(65);
output(1, 63) <= input(66);
output(1, 64) <= input(73);
output(1, 65) <= input(72);
output(1, 66) <= input(71);
output(1, 67) <= input(70);
output(1, 68) <= input(54);
output(1, 69) <= input(55);
output(1, 70) <= input(56);
output(1, 71) <= input(57);
output(1, 72) <= input(58);
output(1, 73) <= input(59);
output(1, 74) <= input(60);
output(1, 75) <= input(61);
output(1, 76) <= input(62);
output(1, 77) <= input(63);
output(1, 78) <= input(64);
output(1, 79) <= input(65);
output(1, 80) <= input(74);
output(1, 81) <= input(73);
output(1, 82) <= input(72);
output(1, 83) <= input(71);
output(1, 84) <= input(70);
output(1, 85) <= input(54);
output(1, 86) <= input(55);
output(1, 87) <= input(56);
output(1, 88) <= input(57);
output(1, 89) <= input(58);
output(1, 90) <= input(59);
output(1, 91) <= input(60);
output(1, 92) <= input(61);
output(1, 93) <= input(62);
output(1, 94) <= input(63);
output(1, 95) <= input(64);
output(1, 96) <= input(75);
output(1, 97) <= input(74);
output(1, 98) <= input(73);
output(1, 99) <= input(72);
output(1, 100) <= input(71);
output(1, 101) <= input(70);
output(1, 102) <= input(54);
output(1, 103) <= input(55);
output(1, 104) <= input(56);
output(1, 105) <= input(57);
output(1, 106) <= input(58);
output(1, 107) <= input(59);
output(1, 108) <= input(60);
output(1, 109) <= input(61);
output(1, 110) <= input(62);
output(1, 111) <= input(63);
output(1, 112) <= input(76);
output(1, 113) <= input(75);
output(1, 114) <= input(74);
output(1, 115) <= input(73);
output(1, 116) <= input(72);
output(1, 117) <= input(71);
output(1, 118) <= input(70);
output(1, 119) <= input(54);
output(1, 120) <= input(55);
output(1, 121) <= input(56);
output(1, 122) <= input(57);
output(1, 123) <= input(58);
output(1, 124) <= input(59);
output(1, 125) <= input(60);
output(1, 126) <= input(61);
output(1, 127) <= input(62);
output(1, 128) <= input(77);
output(1, 129) <= input(76);
output(1, 130) <= input(75);
output(1, 131) <= input(74);
output(1, 132) <= input(73);
output(1, 133) <= input(72);
output(1, 134) <= input(71);
output(1, 135) <= input(70);
output(1, 136) <= input(54);
output(1, 137) <= input(55);
output(1, 138) <= input(56);
output(1, 139) <= input(57);
output(1, 140) <= input(58);
output(1, 141) <= input(59);
output(1, 142) <= input(60);
output(1, 143) <= input(61);
output(1, 144) <= input(78);
output(1, 145) <= input(77);
output(1, 146) <= input(76);
output(1, 147) <= input(75);
output(1, 148) <= input(74);
output(1, 149) <= input(73);
output(1, 150) <= input(72);
output(1, 151) <= input(71);
output(1, 152) <= input(70);
output(1, 153) <= input(54);
output(1, 154) <= input(55);
output(1, 155) <= input(56);
output(1, 156) <= input(57);
output(1, 157) <= input(58);
output(1, 158) <= input(59);
output(1, 159) <= input(60);
output(1, 160) <= input(79);
output(1, 161) <= input(78);
output(1, 162) <= input(77);
output(1, 163) <= input(76);
output(1, 164) <= input(75);
output(1, 165) <= input(74);
output(1, 166) <= input(73);
output(1, 167) <= input(72);
output(1, 168) <= input(71);
output(1, 169) <= input(70);
output(1, 170) <= input(54);
output(1, 171) <= input(55);
output(1, 172) <= input(56);
output(1, 173) <= input(57);
output(1, 174) <= input(58);
output(1, 175) <= input(59);
output(1, 176) <= input(80);
output(1, 177) <= input(79);
output(1, 178) <= input(78);
output(1, 179) <= input(77);
output(1, 180) <= input(76);
output(1, 181) <= input(75);
output(1, 182) <= input(74);
output(1, 183) <= input(73);
output(1, 184) <= input(72);
output(1, 185) <= input(71);
output(1, 186) <= input(70);
output(1, 187) <= input(54);
output(1, 188) <= input(55);
output(1, 189) <= input(56);
output(1, 190) <= input(57);
output(1, 191) <= input(58);
output(1, 192) <= input(81);
output(1, 193) <= input(80);
output(1, 194) <= input(79);
output(1, 195) <= input(78);
output(1, 196) <= input(77);
output(1, 197) <= input(76);
output(1, 198) <= input(75);
output(1, 199) <= input(74);
output(1, 200) <= input(73);
output(1, 201) <= input(72);
output(1, 202) <= input(71);
output(1, 203) <= input(70);
output(1, 204) <= input(54);
output(1, 205) <= input(55);
output(1, 206) <= input(56);
output(1, 207) <= input(57);
output(1, 208) <= input(82);
output(1, 209) <= input(81);
output(1, 210) <= input(80);
output(1, 211) <= input(79);
output(1, 212) <= input(78);
output(1, 213) <= input(77);
output(1, 214) <= input(76);
output(1, 215) <= input(75);
output(1, 216) <= input(74);
output(1, 217) <= input(73);
output(1, 218) <= input(72);
output(1, 219) <= input(71);
output(1, 220) <= input(70);
output(1, 221) <= input(54);
output(1, 222) <= input(55);
output(1, 223) <= input(56);
output(1, 224) <= input(83);
output(1, 225) <= input(82);
output(1, 226) <= input(81);
output(1, 227) <= input(80);
output(1, 228) <= input(79);
output(1, 229) <= input(78);
output(1, 230) <= input(77);
output(1, 231) <= input(76);
output(1, 232) <= input(75);
output(1, 233) <= input(74);
output(1, 234) <= input(73);
output(1, 235) <= input(72);
output(1, 236) <= input(71);
output(1, 237) <= input(70);
output(1, 238) <= input(54);
output(1, 239) <= input(55);
output(1, 240) <= input(84);
output(1, 241) <= input(83);
output(1, 242) <= input(82);
output(1, 243) <= input(81);
output(1, 244) <= input(80);
output(1, 245) <= input(79);
output(1, 246) <= input(78);
output(1, 247) <= input(77);
output(1, 248) <= input(76);
output(1, 249) <= input(75);
output(1, 250) <= input(74);
output(1, 251) <= input(73);
output(1, 252) <= input(72);
output(1, 253) <= input(71);
output(1, 254) <= input(70);
output(1, 255) <= input(54);
when "1000" =>
output(0, 0) <= input(0);
output(0, 1) <= input(1);
output(0, 2) <= input(2);
output(0, 3) <= input(3);
output(0, 4) <= input(4);
output(0, 5) <= input(5);
output(0, 6) <= input(6);
output(0, 7) <= input(7);
output(0, 8) <= input(8);
output(0, 9) <= input(9);
output(0, 10) <= input(10);
output(0, 11) <= input(11);
output(0, 12) <= input(12);
output(0, 13) <= input(13);
output(0, 14) <= input(14);
output(0, 15) <= input(15);
output(0, 16) <= input(16);
output(0, 17) <= input(0);
output(0, 18) <= input(1);
output(0, 19) <= input(2);
output(0, 20) <= input(3);
output(0, 21) <= input(4);
output(0, 22) <= input(5);
output(0, 23) <= input(6);
output(0, 24) <= input(7);
output(0, 25) <= input(8);
output(0, 26) <= input(9);
output(0, 27) <= input(10);
output(0, 28) <= input(11);
output(0, 29) <= input(12);
output(0, 30) <= input(13);
output(0, 31) <= input(14);
output(0, 32) <= input(17);
output(0, 33) <= input(16);
output(0, 34) <= input(0);
output(0, 35) <= input(1);
output(0, 36) <= input(2);
output(0, 37) <= input(3);
output(0, 38) <= input(4);
output(0, 39) <= input(5);
output(0, 40) <= input(6);
output(0, 41) <= input(7);
output(0, 42) <= input(8);
output(0, 43) <= input(9);
output(0, 44) <= input(10);
output(0, 45) <= input(11);
output(0, 46) <= input(12);
output(0, 47) <= input(13);
output(0, 48) <= input(18);
output(0, 49) <= input(17);
output(0, 50) <= input(16);
output(0, 51) <= input(0);
output(0, 52) <= input(1);
output(0, 53) <= input(2);
output(0, 54) <= input(3);
output(0, 55) <= input(4);
output(0, 56) <= input(5);
output(0, 57) <= input(6);
output(0, 58) <= input(7);
output(0, 59) <= input(8);
output(0, 60) <= input(9);
output(0, 61) <= input(10);
output(0, 62) <= input(11);
output(0, 63) <= input(12);
output(0, 64) <= input(19);
output(0, 65) <= input(18);
output(0, 66) <= input(17);
output(0, 67) <= input(16);
output(0, 68) <= input(0);
output(0, 69) <= input(1);
output(0, 70) <= input(2);
output(0, 71) <= input(3);
output(0, 72) <= input(4);
output(0, 73) <= input(5);
output(0, 74) <= input(6);
output(0, 75) <= input(7);
output(0, 76) <= input(8);
output(0, 77) <= input(9);
output(0, 78) <= input(10);
output(0, 79) <= input(11);
output(0, 80) <= input(20);
output(0, 81) <= input(21);
output(0, 82) <= input(22);
output(0, 83) <= input(23);
output(0, 84) <= input(24);
output(0, 85) <= input(25);
output(0, 86) <= input(26);
output(0, 87) <= input(27);
output(0, 88) <= input(28);
output(0, 89) <= input(29);
output(0, 90) <= input(30);
output(0, 91) <= input(31);
output(0, 92) <= input(32);
output(0, 93) <= input(33);
output(0, 94) <= input(34);
output(0, 95) <= input(35);
output(0, 96) <= input(36);
output(0, 97) <= input(20);
output(0, 98) <= input(21);
output(0, 99) <= input(22);
output(0, 100) <= input(23);
output(0, 101) <= input(24);
output(0, 102) <= input(25);
output(0, 103) <= input(26);
output(0, 104) <= input(27);
output(0, 105) <= input(28);
output(0, 106) <= input(29);
output(0, 107) <= input(30);
output(0, 108) <= input(31);
output(0, 109) <= input(32);
output(0, 110) <= input(33);
output(0, 111) <= input(34);
output(0, 112) <= input(37);
output(0, 113) <= input(36);
output(0, 114) <= input(20);
output(0, 115) <= input(21);
output(0, 116) <= input(22);
output(0, 117) <= input(23);
output(0, 118) <= input(24);
output(0, 119) <= input(25);
output(0, 120) <= input(26);
output(0, 121) <= input(27);
output(0, 122) <= input(28);
output(0, 123) <= input(29);
output(0, 124) <= input(30);
output(0, 125) <= input(31);
output(0, 126) <= input(32);
output(0, 127) <= input(33);
output(0, 128) <= input(38);
output(0, 129) <= input(37);
output(0, 130) <= input(36);
output(0, 131) <= input(20);
output(0, 132) <= input(21);
output(0, 133) <= input(22);
output(0, 134) <= input(23);
output(0, 135) <= input(24);
output(0, 136) <= input(25);
output(0, 137) <= input(26);
output(0, 138) <= input(27);
output(0, 139) <= input(28);
output(0, 140) <= input(29);
output(0, 141) <= input(30);
output(0, 142) <= input(31);
output(0, 143) <= input(32);
output(0, 144) <= input(39);
output(0, 145) <= input(38);
output(0, 146) <= input(37);
output(0, 147) <= input(36);
output(0, 148) <= input(20);
output(0, 149) <= input(21);
output(0, 150) <= input(22);
output(0, 151) <= input(23);
output(0, 152) <= input(24);
output(0, 153) <= input(25);
output(0, 154) <= input(26);
output(0, 155) <= input(27);
output(0, 156) <= input(28);
output(0, 157) <= input(29);
output(0, 158) <= input(30);
output(0, 159) <= input(31);
output(0, 160) <= input(40);
output(0, 161) <= input(41);
output(0, 162) <= input(42);
output(0, 163) <= input(43);
output(0, 164) <= input(44);
output(0, 165) <= input(19);
output(0, 166) <= input(18);
output(0, 167) <= input(17);
output(0, 168) <= input(16);
output(0, 169) <= input(0);
output(0, 170) <= input(1);
output(0, 171) <= input(2);
output(0, 172) <= input(3);
output(0, 173) <= input(4);
output(0, 174) <= input(5);
output(0, 175) <= input(6);
output(0, 176) <= input(45);
output(0, 177) <= input(40);
output(0, 178) <= input(41);
output(0, 179) <= input(42);
output(0, 180) <= input(43);
output(0, 181) <= input(44);
output(0, 182) <= input(19);
output(0, 183) <= input(18);
output(0, 184) <= input(17);
output(0, 185) <= input(16);
output(0, 186) <= input(0);
output(0, 187) <= input(1);
output(0, 188) <= input(2);
output(0, 189) <= input(3);
output(0, 190) <= input(4);
output(0, 191) <= input(5);
output(0, 192) <= input(46);
output(0, 193) <= input(45);
output(0, 194) <= input(40);
output(0, 195) <= input(41);
output(0, 196) <= input(42);
output(0, 197) <= input(43);
output(0, 198) <= input(44);
output(0, 199) <= input(19);
output(0, 200) <= input(18);
output(0, 201) <= input(17);
output(0, 202) <= input(16);
output(0, 203) <= input(0);
output(0, 204) <= input(1);
output(0, 205) <= input(2);
output(0, 206) <= input(3);
output(0, 207) <= input(4);
output(0, 208) <= input(47);
output(0, 209) <= input(46);
output(0, 210) <= input(45);
output(0, 211) <= input(40);
output(0, 212) <= input(41);
output(0, 213) <= input(42);
output(0, 214) <= input(43);
output(0, 215) <= input(44);
output(0, 216) <= input(19);
output(0, 217) <= input(18);
output(0, 218) <= input(17);
output(0, 219) <= input(16);
output(0, 220) <= input(0);
output(0, 221) <= input(1);
output(0, 222) <= input(2);
output(0, 223) <= input(3);
output(0, 224) <= input(48);
output(0, 225) <= input(47);
output(0, 226) <= input(46);
output(0, 227) <= input(45);
output(0, 228) <= input(40);
output(0, 229) <= input(41);
output(0, 230) <= input(42);
output(0, 231) <= input(43);
output(0, 232) <= input(44);
output(0, 233) <= input(19);
output(0, 234) <= input(18);
output(0, 235) <= input(17);
output(0, 236) <= input(16);
output(0, 237) <= input(0);
output(0, 238) <= input(1);
output(0, 239) <= input(2);
output(0, 240) <= input(49);
output(0, 241) <= input(50);
output(0, 242) <= input(51);
output(0, 243) <= input(52);
output(0, 244) <= input(53);
output(0, 245) <= input(39);
output(0, 246) <= input(38);
output(0, 247) <= input(37);
output(0, 248) <= input(36);
output(0, 249) <= input(20);
output(0, 250) <= input(21);
output(0, 251) <= input(22);
output(0, 252) <= input(23);
output(0, 253) <= input(24);
output(0, 254) <= input(25);
output(0, 255) <= input(26);
when "1001" =>
output(0, 0) <= input(0);
output(0, 1) <= input(1);
output(0, 2) <= input(2);
output(0, 3) <= input(3);
output(0, 4) <= input(4);
output(0, 5) <= input(5);
output(0, 6) <= input(6);
output(0, 7) <= input(7);
output(0, 8) <= input(8);
output(0, 9) <= input(9);
output(0, 10) <= input(10);
output(0, 11) <= input(11);
output(0, 12) <= input(12);
output(0, 13) <= input(13);
output(0, 14) <= input(14);
output(0, 15) <= input(15);
output(0, 16) <= input(16);
output(0, 17) <= input(0);
output(0, 18) <= input(1);
output(0, 19) <= input(2);
output(0, 20) <= input(3);
output(0, 21) <= input(4);
output(0, 22) <= input(5);
output(0, 23) <= input(6);
output(0, 24) <= input(7);
output(0, 25) <= input(8);
output(0, 26) <= input(9);
output(0, 27) <= input(10);
output(0, 28) <= input(11);
output(0, 29) <= input(12);
output(0, 30) <= input(13);
output(0, 31) <= input(14);
output(0, 32) <= input(17);
output(0, 33) <= input(18);
output(0, 34) <= input(19);
output(0, 35) <= input(20);
output(0, 36) <= input(21);
output(0, 37) <= input(22);
output(0, 38) <= input(23);
output(0, 39) <= input(24);
output(0, 40) <= input(25);
output(0, 41) <= input(26);
output(0, 42) <= input(27);
output(0, 43) <= input(28);
output(0, 44) <= input(29);
output(0, 45) <= input(30);
output(0, 46) <= input(31);
output(0, 47) <= input(32);
output(0, 48) <= input(33);
output(0, 49) <= input(17);
output(0, 50) <= input(18);
output(0, 51) <= input(19);
output(0, 52) <= input(20);
output(0, 53) <= input(21);
output(0, 54) <= input(22);
output(0, 55) <= input(23);
output(0, 56) <= input(24);
output(0, 57) <= input(25);
output(0, 58) <= input(26);
output(0, 59) <= input(27);
output(0, 60) <= input(28);
output(0, 61) <= input(29);
output(0, 62) <= input(30);
output(0, 63) <= input(31);
output(0, 64) <= input(34);
output(0, 65) <= input(33);
output(0, 66) <= input(17);
output(0, 67) <= input(18);
output(0, 68) <= input(19);
output(0, 69) <= input(20);
output(0, 70) <= input(21);
output(0, 71) <= input(22);
output(0, 72) <= input(23);
output(0, 73) <= input(24);
output(0, 74) <= input(25);
output(0, 75) <= input(26);
output(0, 76) <= input(27);
output(0, 77) <= input(28);
output(0, 78) <= input(29);
output(0, 79) <= input(30);
output(0, 80) <= input(35);
output(0, 81) <= input(36);
output(0, 82) <= input(37);
output(0, 83) <= input(16);
output(0, 84) <= input(0);
output(0, 85) <= input(1);
output(0, 86) <= input(2);
output(0, 87) <= input(3);
output(0, 88) <= input(4);
output(0, 89) <= input(5);
output(0, 90) <= input(6);
output(0, 91) <= input(7);
output(0, 92) <= input(8);
output(0, 93) <= input(9);
output(0, 94) <= input(10);
output(0, 95) <= input(11);
output(0, 96) <= input(38);
output(0, 97) <= input(35);
output(0, 98) <= input(36);
output(0, 99) <= input(37);
output(0, 100) <= input(16);
output(0, 101) <= input(0);
output(0, 102) <= input(1);
output(0, 103) <= input(2);
output(0, 104) <= input(3);
output(0, 105) <= input(4);
output(0, 106) <= input(5);
output(0, 107) <= input(6);
output(0, 108) <= input(7);
output(0, 109) <= input(8);
output(0, 110) <= input(9);
output(0, 111) <= input(10);
output(0, 112) <= input(39);
output(0, 113) <= input(40);
output(0, 114) <= input(34);
output(0, 115) <= input(33);
output(0, 116) <= input(17);
output(0, 117) <= input(18);
output(0, 118) <= input(19);
output(0, 119) <= input(20);
output(0, 120) <= input(21);
output(0, 121) <= input(22);
output(0, 122) <= input(23);
output(0, 123) <= input(24);
output(0, 124) <= input(25);
output(0, 125) <= input(26);
output(0, 126) <= input(27);
output(0, 127) <= input(28);
output(0, 128) <= input(41);
output(0, 129) <= input(39);
output(0, 130) <= input(40);
output(0, 131) <= input(34);
output(0, 132) <= input(33);
output(0, 133) <= input(17);
output(0, 134) <= input(18);
output(0, 135) <= input(19);
output(0, 136) <= input(20);
output(0, 137) <= input(21);
output(0, 138) <= input(22);
output(0, 139) <= input(23);
output(0, 140) <= input(24);
output(0, 141) <= input(25);
output(0, 142) <= input(26);
output(0, 143) <= input(27);
output(0, 144) <= input(42);
output(0, 145) <= input(41);
output(0, 146) <= input(39);
output(0, 147) <= input(40);
output(0, 148) <= input(34);
output(0, 149) <= input(33);
output(0, 150) <= input(17);
output(0, 151) <= input(18);
output(0, 152) <= input(19);
output(0, 153) <= input(20);
output(0, 154) <= input(21);
output(0, 155) <= input(22);
output(0, 156) <= input(23);
output(0, 157) <= input(24);
output(0, 158) <= input(25);
output(0, 159) <= input(26);
output(0, 160) <= input(43);
output(0, 161) <= input(44);
output(0, 162) <= input(45);
output(0, 163) <= input(38);
output(0, 164) <= input(35);
output(0, 165) <= input(36);
output(0, 166) <= input(37);
output(0, 167) <= input(16);
output(0, 168) <= input(0);
output(0, 169) <= input(1);
output(0, 170) <= input(2);
output(0, 171) <= input(3);
output(0, 172) <= input(4);
output(0, 173) <= input(5);
output(0, 174) <= input(6);
output(0, 175) <= input(7);
output(0, 176) <= input(46);
output(0, 177) <= input(43);
output(0, 178) <= input(44);
output(0, 179) <= input(45);
output(0, 180) <= input(38);
output(0, 181) <= input(35);
output(0, 182) <= input(36);
output(0, 183) <= input(37);
output(0, 184) <= input(16);
output(0, 185) <= input(0);
output(0, 186) <= input(1);
output(0, 187) <= input(2);
output(0, 188) <= input(3);
output(0, 189) <= input(4);
output(0, 190) <= input(5);
output(0, 191) <= input(6);
output(0, 192) <= input(47);
output(0, 193) <= input(46);
output(0, 194) <= input(43);
output(0, 195) <= input(44);
output(0, 196) <= input(45);
output(0, 197) <= input(38);
output(0, 198) <= input(35);
output(0, 199) <= input(36);
output(0, 200) <= input(37);
output(0, 201) <= input(16);
output(0, 202) <= input(0);
output(0, 203) <= input(1);
output(0, 204) <= input(2);
output(0, 205) <= input(3);
output(0, 206) <= input(4);
output(0, 207) <= input(5);
output(0, 208) <= input(48);
output(0, 209) <= input(49);
output(0, 210) <= input(50);
output(0, 211) <= input(42);
output(0, 212) <= input(41);
output(0, 213) <= input(39);
output(0, 214) <= input(40);
output(0, 215) <= input(34);
output(0, 216) <= input(33);
output(0, 217) <= input(17);
output(0, 218) <= input(18);
output(0, 219) <= input(19);
output(0, 220) <= input(20);
output(0, 221) <= input(21);
output(0, 222) <= input(22);
output(0, 223) <= input(23);
output(0, 224) <= input(51);
output(0, 225) <= input(48);
output(0, 226) <= input(49);
output(0, 227) <= input(50);
output(0, 228) <= input(42);
output(0, 229) <= input(41);
output(0, 230) <= input(39);
output(0, 231) <= input(40);
output(0, 232) <= input(34);
output(0, 233) <= input(33);
output(0, 234) <= input(17);
output(0, 235) <= input(18);
output(0, 236) <= input(19);
output(0, 237) <= input(20);
output(0, 238) <= input(21);
output(0, 239) <= input(22);
output(0, 240) <= input(52);
output(0, 241) <= input(53);
output(0, 242) <= input(47);
output(0, 243) <= input(46);
output(0, 244) <= input(43);
output(0, 245) <= input(44);
output(0, 246) <= input(45);
output(0, 247) <= input(38);
output(0, 248) <= input(35);
output(0, 249) <= input(36);
output(0, 250) <= input(37);
output(0, 251) <= input(16);
output(0, 252) <= input(0);
output(0, 253) <= input(1);
output(0, 254) <= input(2);
output(0, 255) <= input(3);
output(1, 0) <= input(0);
output(1, 1) <= input(1);
output(1, 2) <= input(2);
output(1, 3) <= input(3);
output(1, 4) <= input(4);
output(1, 5) <= input(5);
output(1, 6) <= input(6);
output(1, 7) <= input(7);
output(1, 8) <= input(8);
output(1, 9) <= input(9);
output(1, 10) <= input(10);
output(1, 11) <= input(11);
output(1, 12) <= input(12);
output(1, 13) <= input(13);
output(1, 14) <= input(14);
output(1, 15) <= input(15);
output(1, 16) <= input(54);
output(1, 17) <= input(19);
output(1, 18) <= input(20);
output(1, 19) <= input(21);
output(1, 20) <= input(22);
output(1, 21) <= input(23);
output(1, 22) <= input(24);
output(1, 23) <= input(25);
output(1, 24) <= input(26);
output(1, 25) <= input(27);
output(1, 26) <= input(28);
output(1, 27) <= input(29);
output(1, 28) <= input(30);
output(1, 29) <= input(31);
output(1, 30) <= input(32);
output(1, 31) <= input(55);
output(1, 32) <= input(56);
output(1, 33) <= input(54);
output(1, 34) <= input(19);
output(1, 35) <= input(20);
output(1, 36) <= input(21);
output(1, 37) <= input(22);
output(1, 38) <= input(23);
output(1, 39) <= input(24);
output(1, 40) <= input(25);
output(1, 41) <= input(26);
output(1, 42) <= input(27);
output(1, 43) <= input(28);
output(1, 44) <= input(29);
output(1, 45) <= input(30);
output(1, 46) <= input(31);
output(1, 47) <= input(32);
output(1, 48) <= input(57);
output(1, 49) <= input(58);
output(1, 50) <= input(0);
output(1, 51) <= input(1);
output(1, 52) <= input(2);
output(1, 53) <= input(3);
output(1, 54) <= input(4);
output(1, 55) <= input(5);
output(1, 56) <= input(6);
output(1, 57) <= input(7);
output(1, 58) <= input(8);
output(1, 59) <= input(9);
output(1, 60) <= input(10);
output(1, 61) <= input(11);
output(1, 62) <= input(12);
output(1, 63) <= input(13);
output(1, 64) <= input(59);
output(1, 65) <= input(57);
output(1, 66) <= input(58);
output(1, 67) <= input(0);
output(1, 68) <= input(1);
output(1, 69) <= input(2);
output(1, 70) <= input(3);
output(1, 71) <= input(4);
output(1, 72) <= input(5);
output(1, 73) <= input(6);
output(1, 74) <= input(7);
output(1, 75) <= input(8);
output(1, 76) <= input(9);
output(1, 77) <= input(10);
output(1, 78) <= input(11);
output(1, 79) <= input(12);
output(1, 80) <= input(60);
output(1, 81) <= input(61);
output(1, 82) <= input(56);
output(1, 83) <= input(54);
output(1, 84) <= input(19);
output(1, 85) <= input(20);
output(1, 86) <= input(21);
output(1, 87) <= input(22);
output(1, 88) <= input(23);
output(1, 89) <= input(24);
output(1, 90) <= input(25);
output(1, 91) <= input(26);
output(1, 92) <= input(27);
output(1, 93) <= input(28);
output(1, 94) <= input(29);
output(1, 95) <= input(30);
output(1, 96) <= input(62);
output(1, 97) <= input(60);
output(1, 98) <= input(61);
output(1, 99) <= input(56);
output(1, 100) <= input(54);
output(1, 101) <= input(19);
output(1, 102) <= input(20);
output(1, 103) <= input(21);
output(1, 104) <= input(22);
output(1, 105) <= input(23);
output(1, 106) <= input(24);
output(1, 107) <= input(25);
output(1, 108) <= input(26);
output(1, 109) <= input(27);
output(1, 110) <= input(28);
output(1, 111) <= input(29);
output(1, 112) <= input(63);
output(1, 113) <= input(64);
output(1, 114) <= input(59);
output(1, 115) <= input(57);
output(1, 116) <= input(58);
output(1, 117) <= input(0);
output(1, 118) <= input(1);
output(1, 119) <= input(2);
output(1, 120) <= input(3);
output(1, 121) <= input(4);
output(1, 122) <= input(5);
output(1, 123) <= input(6);
output(1, 124) <= input(7);
output(1, 125) <= input(8);
output(1, 126) <= input(9);
output(1, 127) <= input(10);
output(1, 128) <= input(65);
output(1, 129) <= input(62);
output(1, 130) <= input(60);
output(1, 131) <= input(61);
output(1, 132) <= input(56);
output(1, 133) <= input(54);
output(1, 134) <= input(19);
output(1, 135) <= input(20);
output(1, 136) <= input(21);
output(1, 137) <= input(22);
output(1, 138) <= input(23);
output(1, 139) <= input(24);
output(1, 140) <= input(25);
output(1, 141) <= input(26);
output(1, 142) <= input(27);
output(1, 143) <= input(28);
output(1, 144) <= input(66);
output(1, 145) <= input(65);
output(1, 146) <= input(62);
output(1, 147) <= input(60);
output(1, 148) <= input(61);
output(1, 149) <= input(56);
output(1, 150) <= input(54);
output(1, 151) <= input(19);
output(1, 152) <= input(20);
output(1, 153) <= input(21);
output(1, 154) <= input(22);
output(1, 155) <= input(23);
output(1, 156) <= input(24);
output(1, 157) <= input(25);
output(1, 158) <= input(26);
output(1, 159) <= input(27);
output(1, 160) <= input(67);
output(1, 161) <= input(68);
output(1, 162) <= input(63);
output(1, 163) <= input(64);
output(1, 164) <= input(59);
output(1, 165) <= input(57);
output(1, 166) <= input(58);
output(1, 167) <= input(0);
output(1, 168) <= input(1);
output(1, 169) <= input(2);
output(1, 170) <= input(3);
output(1, 171) <= input(4);
output(1, 172) <= input(5);
output(1, 173) <= input(6);
output(1, 174) <= input(7);
output(1, 175) <= input(8);
output(1, 176) <= input(69);
output(1, 177) <= input(67);
output(1, 178) <= input(68);
output(1, 179) <= input(63);
output(1, 180) <= input(64);
output(1, 181) <= input(59);
output(1, 182) <= input(57);
output(1, 183) <= input(58);
output(1, 184) <= input(0);
output(1, 185) <= input(1);
output(1, 186) <= input(2);
output(1, 187) <= input(3);
output(1, 188) <= input(4);
output(1, 189) <= input(5);
output(1, 190) <= input(6);
output(1, 191) <= input(7);
output(1, 192) <= input(70);
output(1, 193) <= input(71);
output(1, 194) <= input(66);
output(1, 195) <= input(65);
output(1, 196) <= input(62);
output(1, 197) <= input(60);
output(1, 198) <= input(61);
output(1, 199) <= input(56);
output(1, 200) <= input(54);
output(1, 201) <= input(19);
output(1, 202) <= input(20);
output(1, 203) <= input(21);
output(1, 204) <= input(22);
output(1, 205) <= input(23);
output(1, 206) <= input(24);
output(1, 207) <= input(25);
output(1, 208) <= input(72);
output(1, 209) <= input(70);
output(1, 210) <= input(71);
output(1, 211) <= input(66);
output(1, 212) <= input(65);
output(1, 213) <= input(62);
output(1, 214) <= input(60);
output(1, 215) <= input(61);
output(1, 216) <= input(56);
output(1, 217) <= input(54);
output(1, 218) <= input(19);
output(1, 219) <= input(20);
output(1, 220) <= input(21);
output(1, 221) <= input(22);
output(1, 222) <= input(23);
output(1, 223) <= input(24);
output(1, 224) <= input(73);
output(1, 225) <= input(74);
output(1, 226) <= input(69);
output(1, 227) <= input(67);
output(1, 228) <= input(68);
output(1, 229) <= input(63);
output(1, 230) <= input(64);
output(1, 231) <= input(59);
output(1, 232) <= input(57);
output(1, 233) <= input(58);
output(1, 234) <= input(0);
output(1, 235) <= input(1);
output(1, 236) <= input(2);
output(1, 237) <= input(3);
output(1, 238) <= input(4);
output(1, 239) <= input(5);
output(1, 240) <= input(75);
output(1, 241) <= input(72);
output(1, 242) <= input(70);
output(1, 243) <= input(71);
output(1, 244) <= input(66);
output(1, 245) <= input(65);
output(1, 246) <= input(62);
output(1, 247) <= input(60);
output(1, 248) <= input(61);
output(1, 249) <= input(56);
output(1, 250) <= input(54);
output(1, 251) <= input(19);
output(1, 252) <= input(20);
output(1, 253) <= input(21);
output(1, 254) <= input(22);
output(1, 255) <= input(23);
output(2, 0) <= input(76);
output(2, 1) <= input(1);
output(2, 2) <= input(2);
output(2, 3) <= input(3);
output(2, 4) <= input(4);
output(2, 5) <= input(5);
output(2, 6) <= input(6);
output(2, 7) <= input(7);
output(2, 8) <= input(8);
output(2, 9) <= input(9);
output(2, 10) <= input(10);
output(2, 11) <= input(11);
output(2, 12) <= input(12);
output(2, 13) <= input(13);
output(2, 14) <= input(14);
output(2, 15) <= input(15);
output(2, 16) <= input(77);
output(2, 17) <= input(78);
output(2, 18) <= input(20);
output(2, 19) <= input(21);
output(2, 20) <= input(22);
output(2, 21) <= input(23);
output(2, 22) <= input(24);
output(2, 23) <= input(25);
output(2, 24) <= input(26);
output(2, 25) <= input(27);
output(2, 26) <= input(28);
output(2, 27) <= input(29);
output(2, 28) <= input(30);
output(2, 29) <= input(31);
output(2, 30) <= input(32);
output(2, 31) <= input(55);
output(2, 32) <= input(79);
output(2, 33) <= input(76);
output(2, 34) <= input(1);
output(2, 35) <= input(2);
output(2, 36) <= input(3);
output(2, 37) <= input(4);
output(2, 38) <= input(5);
output(2, 39) <= input(6);
output(2, 40) <= input(7);
output(2, 41) <= input(8);
output(2, 42) <= input(9);
output(2, 43) <= input(10);
output(2, 44) <= input(11);
output(2, 45) <= input(12);
output(2, 46) <= input(13);
output(2, 47) <= input(14);
output(2, 48) <= input(80);
output(2, 49) <= input(77);
output(2, 50) <= input(78);
output(2, 51) <= input(20);
output(2, 52) <= input(21);
output(2, 53) <= input(22);
output(2, 54) <= input(23);
output(2, 55) <= input(24);
output(2, 56) <= input(25);
output(2, 57) <= input(26);
output(2, 58) <= input(27);
output(2, 59) <= input(28);
output(2, 60) <= input(29);
output(2, 61) <= input(30);
output(2, 62) <= input(31);
output(2, 63) <= input(32);
output(2, 64) <= input(81);
output(2, 65) <= input(80);
output(2, 66) <= input(77);
output(2, 67) <= input(78);
output(2, 68) <= input(20);
output(2, 69) <= input(21);
output(2, 70) <= input(22);
output(2, 71) <= input(23);
output(2, 72) <= input(24);
output(2, 73) <= input(25);
output(2, 74) <= input(26);
output(2, 75) <= input(27);
output(2, 76) <= input(28);
output(2, 77) <= input(29);
output(2, 78) <= input(30);
output(2, 79) <= input(31);
output(2, 80) <= input(82);
output(2, 81) <= input(83);
output(2, 82) <= input(79);
output(2, 83) <= input(76);
output(2, 84) <= input(1);
output(2, 85) <= input(2);
output(2, 86) <= input(3);
output(2, 87) <= input(4);
output(2, 88) <= input(5);
output(2, 89) <= input(6);
output(2, 90) <= input(7);
output(2, 91) <= input(8);
output(2, 92) <= input(9);
output(2, 93) <= input(10);
output(2, 94) <= input(11);
output(2, 95) <= input(12);
output(2, 96) <= input(84);
output(2, 97) <= input(81);
output(2, 98) <= input(80);
output(2, 99) <= input(77);
output(2, 100) <= input(78);
output(2, 101) <= input(20);
output(2, 102) <= input(21);
output(2, 103) <= input(22);
output(2, 104) <= input(23);
output(2, 105) <= input(24);
output(2, 106) <= input(25);
output(2, 107) <= input(26);
output(2, 108) <= input(27);
output(2, 109) <= input(28);
output(2, 110) <= input(29);
output(2, 111) <= input(30);
output(2, 112) <= input(85);
output(2, 113) <= input(82);
output(2, 114) <= input(83);
output(2, 115) <= input(79);
output(2, 116) <= input(76);
output(2, 117) <= input(1);
output(2, 118) <= input(2);
output(2, 119) <= input(3);
output(2, 120) <= input(4);
output(2, 121) <= input(5);
output(2, 122) <= input(6);
output(2, 123) <= input(7);
output(2, 124) <= input(8);
output(2, 125) <= input(9);
output(2, 126) <= input(10);
output(2, 127) <= input(11);
output(2, 128) <= input(86);
output(2, 129) <= input(85);
output(2, 130) <= input(82);
output(2, 131) <= input(83);
output(2, 132) <= input(79);
output(2, 133) <= input(76);
output(2, 134) <= input(1);
output(2, 135) <= input(2);
output(2, 136) <= input(3);
output(2, 137) <= input(4);
output(2, 138) <= input(5);
output(2, 139) <= input(6);
output(2, 140) <= input(7);
output(2, 141) <= input(8);
output(2, 142) <= input(9);
output(2, 143) <= input(10);
output(2, 144) <= input(87);
output(2, 145) <= input(88);
output(2, 146) <= input(84);
output(2, 147) <= input(81);
output(2, 148) <= input(80);
output(2, 149) <= input(77);
output(2, 150) <= input(78);
output(2, 151) <= input(20);
output(2, 152) <= input(21);
output(2, 153) <= input(22);
output(2, 154) <= input(23);
output(2, 155) <= input(24);
output(2, 156) <= input(25);
output(2, 157) <= input(26);
output(2, 158) <= input(27);
output(2, 159) <= input(28);
output(2, 160) <= input(89);
output(2, 161) <= input(86);
output(2, 162) <= input(85);
output(2, 163) <= input(82);
output(2, 164) <= input(83);
output(2, 165) <= input(79);
output(2, 166) <= input(76);
output(2, 167) <= input(1);
output(2, 168) <= input(2);
output(2, 169) <= input(3);
output(2, 170) <= input(4);
output(2, 171) <= input(5);
output(2, 172) <= input(6);
output(2, 173) <= input(7);
output(2, 174) <= input(8);
output(2, 175) <= input(9);
output(2, 176) <= input(71);
output(2, 177) <= input(87);
output(2, 178) <= input(88);
output(2, 179) <= input(84);
output(2, 180) <= input(81);
output(2, 181) <= input(80);
output(2, 182) <= input(77);
output(2, 183) <= input(78);
output(2, 184) <= input(20);
output(2, 185) <= input(21);
output(2, 186) <= input(22);
output(2, 187) <= input(23);
output(2, 188) <= input(24);
output(2, 189) <= input(25);
output(2, 190) <= input(26);
output(2, 191) <= input(27);
output(2, 192) <= input(70);
output(2, 193) <= input(71);
output(2, 194) <= input(87);
output(2, 195) <= input(88);
output(2, 196) <= input(84);
output(2, 197) <= input(81);
output(2, 198) <= input(80);
output(2, 199) <= input(77);
output(2, 200) <= input(78);
output(2, 201) <= input(20);
output(2, 202) <= input(21);
output(2, 203) <= input(22);
output(2, 204) <= input(23);
output(2, 205) <= input(24);
output(2, 206) <= input(25);
output(2, 207) <= input(26);
output(2, 208) <= input(74);
output(2, 209) <= input(69);
output(2, 210) <= input(89);
output(2, 211) <= input(86);
output(2, 212) <= input(85);
output(2, 213) <= input(82);
output(2, 214) <= input(83);
output(2, 215) <= input(79);
output(2, 216) <= input(76);
output(2, 217) <= input(1);
output(2, 218) <= input(2);
output(2, 219) <= input(3);
output(2, 220) <= input(4);
output(2, 221) <= input(5);
output(2, 222) <= input(6);
output(2, 223) <= input(7);
output(2, 224) <= input(90);
output(2, 225) <= input(70);
output(2, 226) <= input(71);
output(2, 227) <= input(87);
output(2, 228) <= input(88);
output(2, 229) <= input(84);
output(2, 230) <= input(81);
output(2, 231) <= input(80);
output(2, 232) <= input(77);
output(2, 233) <= input(78);
output(2, 234) <= input(20);
output(2, 235) <= input(21);
output(2, 236) <= input(22);
output(2, 237) <= input(23);
output(2, 238) <= input(24);
output(2, 239) <= input(25);
output(2, 240) <= input(91);
output(2, 241) <= input(74);
output(2, 242) <= input(69);
output(2, 243) <= input(89);
output(2, 244) <= input(86);
output(2, 245) <= input(85);
output(2, 246) <= input(82);
output(2, 247) <= input(83);
output(2, 248) <= input(79);
output(2, 249) <= input(76);
output(2, 250) <= input(1);
output(2, 251) <= input(2);
output(2, 252) <= input(3);
output(2, 253) <= input(4);
output(2, 254) <= input(5);
output(2, 255) <= input(6);
when "1010" =>
output(0, 0) <= input(0);
output(0, 1) <= input(1);
output(0, 2) <= input(2);
output(0, 3) <= input(3);
output(0, 4) <= input(4);
output(0, 5) <= input(5);
output(0, 6) <= input(6);
output(0, 7) <= input(7);
output(0, 8) <= input(8);
output(0, 9) <= input(9);
output(0, 10) <= input(10);
output(0, 11) <= input(11);
output(0, 12) <= input(12);
output(0, 13) <= input(13);
output(0, 14) <= input(14);
output(0, 15) <= input(15);
output(0, 16) <= input(16);
output(0, 17) <= input(17);
output(0, 18) <= input(18);
output(0, 19) <= input(19);
output(0, 20) <= input(20);
output(0, 21) <= input(21);
output(0, 22) <= input(22);
output(0, 23) <= input(23);
output(0, 24) <= input(24);
output(0, 25) <= input(25);
output(0, 26) <= input(26);
output(0, 27) <= input(27);
output(0, 28) <= input(28);
output(0, 29) <= input(29);
output(0, 30) <= input(30);
output(0, 31) <= input(31);
output(0, 32) <= input(32);
output(0, 33) <= input(0);
output(0, 34) <= input(1);
output(0, 35) <= input(2);
output(0, 36) <= input(3);
output(0, 37) <= input(4);
output(0, 38) <= input(5);
output(0, 39) <= input(6);
output(0, 40) <= input(7);
output(0, 41) <= input(8);
output(0, 42) <= input(9);
output(0, 43) <= input(10);
output(0, 44) <= input(11);
output(0, 45) <= input(12);
output(0, 46) <= input(13);
output(0, 47) <= input(14);
output(0, 48) <= input(33);
output(0, 49) <= input(16);
output(0, 50) <= input(17);
output(0, 51) <= input(18);
output(0, 52) <= input(19);
output(0, 53) <= input(20);
output(0, 54) <= input(21);
output(0, 55) <= input(22);
output(0, 56) <= input(23);
output(0, 57) <= input(24);
output(0, 58) <= input(25);
output(0, 59) <= input(26);
output(0, 60) <= input(27);
output(0, 61) <= input(28);
output(0, 62) <= input(29);
output(0, 63) <= input(30);
output(0, 64) <= input(34);
output(0, 65) <= input(32);
output(0, 66) <= input(0);
output(0, 67) <= input(1);
output(0, 68) <= input(2);
output(0, 69) <= input(3);
output(0, 70) <= input(4);
output(0, 71) <= input(5);
output(0, 72) <= input(6);
output(0, 73) <= input(7);
output(0, 74) <= input(8);
output(0, 75) <= input(9);
output(0, 76) <= input(10);
output(0, 77) <= input(11);
output(0, 78) <= input(12);
output(0, 79) <= input(13);
output(0, 80) <= input(35);
output(0, 81) <= input(33);
output(0, 82) <= input(16);
output(0, 83) <= input(17);
output(0, 84) <= input(18);
output(0, 85) <= input(19);
output(0, 86) <= input(20);
output(0, 87) <= input(21);
output(0, 88) <= input(22);
output(0, 89) <= input(23);
output(0, 90) <= input(24);
output(0, 91) <= input(25);
output(0, 92) <= input(26);
output(0, 93) <= input(27);
output(0, 94) <= input(28);
output(0, 95) <= input(29);
output(0, 96) <= input(36);
output(0, 97) <= input(34);
output(0, 98) <= input(32);
output(0, 99) <= input(0);
output(0, 100) <= input(1);
output(0, 101) <= input(2);
output(0, 102) <= input(3);
output(0, 103) <= input(4);
output(0, 104) <= input(5);
output(0, 105) <= input(6);
output(0, 106) <= input(7);
output(0, 107) <= input(8);
output(0, 108) <= input(9);
output(0, 109) <= input(10);
output(0, 110) <= input(11);
output(0, 111) <= input(12);
output(0, 112) <= input(37);
output(0, 113) <= input(35);
output(0, 114) <= input(33);
output(0, 115) <= input(16);
output(0, 116) <= input(17);
output(0, 117) <= input(18);
output(0, 118) <= input(19);
output(0, 119) <= input(20);
output(0, 120) <= input(21);
output(0, 121) <= input(22);
output(0, 122) <= input(23);
output(0, 123) <= input(24);
output(0, 124) <= input(25);
output(0, 125) <= input(26);
output(0, 126) <= input(27);
output(0, 127) <= input(28);
output(0, 128) <= input(38);
output(0, 129) <= input(37);
output(0, 130) <= input(35);
output(0, 131) <= input(33);
output(0, 132) <= input(16);
output(0, 133) <= input(17);
output(0, 134) <= input(18);
output(0, 135) <= input(19);
output(0, 136) <= input(20);
output(0, 137) <= input(21);
output(0, 138) <= input(22);
output(0, 139) <= input(23);
output(0, 140) <= input(24);
output(0, 141) <= input(25);
output(0, 142) <= input(26);
output(0, 143) <= input(27);
output(0, 144) <= input(39);
output(0, 145) <= input(40);
output(0, 146) <= input(36);
output(0, 147) <= input(34);
output(0, 148) <= input(32);
output(0, 149) <= input(0);
output(0, 150) <= input(1);
output(0, 151) <= input(2);
output(0, 152) <= input(3);
output(0, 153) <= input(4);
output(0, 154) <= input(5);
output(0, 155) <= input(6);
output(0, 156) <= input(7);
output(0, 157) <= input(8);
output(0, 158) <= input(9);
output(0, 159) <= input(10);
output(0, 160) <= input(41);
output(0, 161) <= input(38);
output(0, 162) <= input(37);
output(0, 163) <= input(35);
output(0, 164) <= input(33);
output(0, 165) <= input(16);
output(0, 166) <= input(17);
output(0, 167) <= input(18);
output(0, 168) <= input(19);
output(0, 169) <= input(20);
output(0, 170) <= input(21);
output(0, 171) <= input(22);
output(0, 172) <= input(23);
output(0, 173) <= input(24);
output(0, 174) <= input(25);
output(0, 175) <= input(26);
output(0, 176) <= input(42);
output(0, 177) <= input(39);
output(0, 178) <= input(40);
output(0, 179) <= input(36);
output(0, 180) <= input(34);
output(0, 181) <= input(32);
output(0, 182) <= input(0);
output(0, 183) <= input(1);
output(0, 184) <= input(2);
output(0, 185) <= input(3);
output(0, 186) <= input(4);
output(0, 187) <= input(5);
output(0, 188) <= input(6);
output(0, 189) <= input(7);
output(0, 190) <= input(8);
output(0, 191) <= input(9);
output(0, 192) <= input(43);
output(0, 193) <= input(41);
output(0, 194) <= input(38);
output(0, 195) <= input(37);
output(0, 196) <= input(35);
output(0, 197) <= input(33);
output(0, 198) <= input(16);
output(0, 199) <= input(17);
output(0, 200) <= input(18);
output(0, 201) <= input(19);
output(0, 202) <= input(20);
output(0, 203) <= input(21);
output(0, 204) <= input(22);
output(0, 205) <= input(23);
output(0, 206) <= input(24);
output(0, 207) <= input(25);
output(0, 208) <= input(44);
output(0, 209) <= input(42);
output(0, 210) <= input(39);
output(0, 211) <= input(40);
output(0, 212) <= input(36);
output(0, 213) <= input(34);
output(0, 214) <= input(32);
output(0, 215) <= input(0);
output(0, 216) <= input(1);
output(0, 217) <= input(2);
output(0, 218) <= input(3);
output(0, 219) <= input(4);
output(0, 220) <= input(5);
output(0, 221) <= input(6);
output(0, 222) <= input(7);
output(0, 223) <= input(8);
output(0, 224) <= input(45);
output(0, 225) <= input(43);
output(0, 226) <= input(41);
output(0, 227) <= input(38);
output(0, 228) <= input(37);
output(0, 229) <= input(35);
output(0, 230) <= input(33);
output(0, 231) <= input(16);
output(0, 232) <= input(17);
output(0, 233) <= input(18);
output(0, 234) <= input(19);
output(0, 235) <= input(20);
output(0, 236) <= input(21);
output(0, 237) <= input(22);
output(0, 238) <= input(23);
output(0, 239) <= input(24);
output(0, 240) <= input(46);
output(0, 241) <= input(44);
output(0, 242) <= input(42);
output(0, 243) <= input(39);
output(0, 244) <= input(40);
output(0, 245) <= input(36);
output(0, 246) <= input(34);
output(0, 247) <= input(32);
output(0, 248) <= input(0);
output(0, 249) <= input(1);
output(0, 250) <= input(2);
output(0, 251) <= input(3);
output(0, 252) <= input(4);
output(0, 253) <= input(5);
output(0, 254) <= input(6);
output(0, 255) <= input(7);
output(1, 0) <= input(17);
output(1, 1) <= input(18);
output(1, 2) <= input(19);
output(1, 3) <= input(20);
output(1, 4) <= input(21);
output(1, 5) <= input(22);
output(1, 6) <= input(23);
output(1, 7) <= input(24);
output(1, 8) <= input(25);
output(1, 9) <= input(26);
output(1, 10) <= input(27);
output(1, 11) <= input(28);
output(1, 12) <= input(29);
output(1, 13) <= input(30);
output(1, 14) <= input(31);
output(1, 15) <= input(47);
output(1, 16) <= input(0);
output(1, 17) <= input(1);
output(1, 18) <= input(2);
output(1, 19) <= input(3);
output(1, 20) <= input(4);
output(1, 21) <= input(5);
output(1, 22) <= input(6);
output(1, 23) <= input(7);
output(1, 24) <= input(8);
output(1, 25) <= input(9);
output(1, 26) <= input(10);
output(1, 27) <= input(11);
output(1, 28) <= input(12);
output(1, 29) <= input(13);
output(1, 30) <= input(14);
output(1, 31) <= input(15);
output(1, 32) <= input(16);
output(1, 33) <= input(17);
output(1, 34) <= input(18);
output(1, 35) <= input(19);
output(1, 36) <= input(20);
output(1, 37) <= input(21);
output(1, 38) <= input(22);
output(1, 39) <= input(23);
output(1, 40) <= input(24);
output(1, 41) <= input(25);
output(1, 42) <= input(26);
output(1, 43) <= input(27);
output(1, 44) <= input(28);
output(1, 45) <= input(29);
output(1, 46) <= input(30);
output(1, 47) <= input(31);
output(1, 48) <= input(32);
output(1, 49) <= input(0);
output(1, 50) <= input(1);
output(1, 51) <= input(2);
output(1, 52) <= input(3);
output(1, 53) <= input(4);
output(1, 54) <= input(5);
output(1, 55) <= input(6);
output(1, 56) <= input(7);
output(1, 57) <= input(8);
output(1, 58) <= input(9);
output(1, 59) <= input(10);
output(1, 60) <= input(11);
output(1, 61) <= input(12);
output(1, 62) <= input(13);
output(1, 63) <= input(14);
output(1, 64) <= input(48);
output(1, 65) <= input(16);
output(1, 66) <= input(17);
output(1, 67) <= input(18);
output(1, 68) <= input(19);
output(1, 69) <= input(20);
output(1, 70) <= input(21);
output(1, 71) <= input(22);
output(1, 72) <= input(23);
output(1, 73) <= input(24);
output(1, 74) <= input(25);
output(1, 75) <= input(26);
output(1, 76) <= input(27);
output(1, 77) <= input(28);
output(1, 78) <= input(29);
output(1, 79) <= input(30);
output(1, 80) <= input(49);
output(1, 81) <= input(32);
output(1, 82) <= input(0);
output(1, 83) <= input(1);
output(1, 84) <= input(2);
output(1, 85) <= input(3);
output(1, 86) <= input(4);
output(1, 87) <= input(5);
output(1, 88) <= input(6);
output(1, 89) <= input(7);
output(1, 90) <= input(8);
output(1, 91) <= input(9);
output(1, 92) <= input(10);
output(1, 93) <= input(11);
output(1, 94) <= input(12);
output(1, 95) <= input(13);
output(1, 96) <= input(50);
output(1, 97) <= input(48);
output(1, 98) <= input(16);
output(1, 99) <= input(17);
output(1, 100) <= input(18);
output(1, 101) <= input(19);
output(1, 102) <= input(20);
output(1, 103) <= input(21);
output(1, 104) <= input(22);
output(1, 105) <= input(23);
output(1, 106) <= input(24);
output(1, 107) <= input(25);
output(1, 108) <= input(26);
output(1, 109) <= input(27);
output(1, 110) <= input(28);
output(1, 111) <= input(29);
output(1, 112) <= input(51);
output(1, 113) <= input(49);
output(1, 114) <= input(32);
output(1, 115) <= input(0);
output(1, 116) <= input(1);
output(1, 117) <= input(2);
output(1, 118) <= input(3);
output(1, 119) <= input(4);
output(1, 120) <= input(5);
output(1, 121) <= input(6);
output(1, 122) <= input(7);
output(1, 123) <= input(8);
output(1, 124) <= input(9);
output(1, 125) <= input(10);
output(1, 126) <= input(11);
output(1, 127) <= input(12);
output(1, 128) <= input(52);
output(1, 129) <= input(50);
output(1, 130) <= input(48);
output(1, 131) <= input(16);
output(1, 132) <= input(17);
output(1, 133) <= input(18);
output(1, 134) <= input(19);
output(1, 135) <= input(20);
output(1, 136) <= input(21);
output(1, 137) <= input(22);
output(1, 138) <= input(23);
output(1, 139) <= input(24);
output(1, 140) <= input(25);
output(1, 141) <= input(26);
output(1, 142) <= input(27);
output(1, 143) <= input(28);
output(1, 144) <= input(53);
output(1, 145) <= input(51);
output(1, 146) <= input(49);
output(1, 147) <= input(32);
output(1, 148) <= input(0);
output(1, 149) <= input(1);
output(1, 150) <= input(2);
output(1, 151) <= input(3);
output(1, 152) <= input(4);
output(1, 153) <= input(5);
output(1, 154) <= input(6);
output(1, 155) <= input(7);
output(1, 156) <= input(8);
output(1, 157) <= input(9);
output(1, 158) <= input(10);
output(1, 159) <= input(11);
output(1, 160) <= input(54);
output(1, 161) <= input(52);
output(1, 162) <= input(50);
output(1, 163) <= input(48);
output(1, 164) <= input(16);
output(1, 165) <= input(17);
output(1, 166) <= input(18);
output(1, 167) <= input(19);
output(1, 168) <= input(20);
output(1, 169) <= input(21);
output(1, 170) <= input(22);
output(1, 171) <= input(23);
output(1, 172) <= input(24);
output(1, 173) <= input(25);
output(1, 174) <= input(26);
output(1, 175) <= input(27);
output(1, 176) <= input(55);
output(1, 177) <= input(53);
output(1, 178) <= input(51);
output(1, 179) <= input(49);
output(1, 180) <= input(32);
output(1, 181) <= input(0);
output(1, 182) <= input(1);
output(1, 183) <= input(2);
output(1, 184) <= input(3);
output(1, 185) <= input(4);
output(1, 186) <= input(5);
output(1, 187) <= input(6);
output(1, 188) <= input(7);
output(1, 189) <= input(8);
output(1, 190) <= input(9);
output(1, 191) <= input(10);
output(1, 192) <= input(56);
output(1, 193) <= input(54);
output(1, 194) <= input(52);
output(1, 195) <= input(50);
output(1, 196) <= input(48);
output(1, 197) <= input(16);
output(1, 198) <= input(17);
output(1, 199) <= input(18);
output(1, 200) <= input(19);
output(1, 201) <= input(20);
output(1, 202) <= input(21);
output(1, 203) <= input(22);
output(1, 204) <= input(23);
output(1, 205) <= input(24);
output(1, 206) <= input(25);
output(1, 207) <= input(26);
output(1, 208) <= input(57);
output(1, 209) <= input(55);
output(1, 210) <= input(53);
output(1, 211) <= input(51);
output(1, 212) <= input(49);
output(1, 213) <= input(32);
output(1, 214) <= input(0);
output(1, 215) <= input(1);
output(1, 216) <= input(2);
output(1, 217) <= input(3);
output(1, 218) <= input(4);
output(1, 219) <= input(5);
output(1, 220) <= input(6);
output(1, 221) <= input(7);
output(1, 222) <= input(8);
output(1, 223) <= input(9);
output(1, 224) <= input(58);
output(1, 225) <= input(56);
output(1, 226) <= input(54);
output(1, 227) <= input(52);
output(1, 228) <= input(50);
output(1, 229) <= input(48);
output(1, 230) <= input(16);
output(1, 231) <= input(17);
output(1, 232) <= input(18);
output(1, 233) <= input(19);
output(1, 234) <= input(20);
output(1, 235) <= input(21);
output(1, 236) <= input(22);
output(1, 237) <= input(23);
output(1, 238) <= input(24);
output(1, 239) <= input(25);
output(1, 240) <= input(59);
output(1, 241) <= input(57);
output(1, 242) <= input(55);
output(1, 243) <= input(53);
output(1, 244) <= input(51);
output(1, 245) <= input(49);
output(1, 246) <= input(32);
output(1, 247) <= input(0);
output(1, 248) <= input(1);
output(1, 249) <= input(2);
output(1, 250) <= input(3);
output(1, 251) <= input(4);
output(1, 252) <= input(5);
output(1, 253) <= input(6);
output(1, 254) <= input(7);
output(1, 255) <= input(8);
when "1011" =>
output(0, 0) <= input(0);
output(0, 1) <= input(1);
output(0, 2) <= input(2);
output(0, 3) <= input(3);
output(0, 4) <= input(4);
output(0, 5) <= input(5);
output(0, 6) <= input(6);
output(0, 7) <= input(7);
output(0, 8) <= input(8);
output(0, 9) <= input(9);
output(0, 10) <= input(10);
output(0, 11) <= input(11);
output(0, 12) <= input(12);
output(0, 13) <= input(13);
output(0, 14) <= input(14);
output(0, 15) <= input(15);
output(0, 16) <= input(16);
output(0, 17) <= input(17);
output(0, 18) <= input(18);
output(0, 19) <= input(19);
output(0, 20) <= input(20);
output(0, 21) <= input(21);
output(0, 22) <= input(22);
output(0, 23) <= input(23);
output(0, 24) <= input(24);
output(0, 25) <= input(25);
output(0, 26) <= input(26);
output(0, 27) <= input(27);
output(0, 28) <= input(28);
output(0, 29) <= input(29);
output(0, 30) <= input(30);
output(0, 31) <= input(31);
output(0, 32) <= input(32);
output(0, 33) <= input(0);
output(0, 34) <= input(1);
output(0, 35) <= input(2);
output(0, 36) <= input(3);
output(0, 37) <= input(4);
output(0, 38) <= input(5);
output(0, 39) <= input(6);
output(0, 40) <= input(7);
output(0, 41) <= input(8);
output(0, 42) <= input(9);
output(0, 43) <= input(10);
output(0, 44) <= input(11);
output(0, 45) <= input(12);
output(0, 46) <= input(13);
output(0, 47) <= input(14);
output(0, 48) <= input(33);
output(0, 49) <= input(16);
output(0, 50) <= input(17);
output(0, 51) <= input(18);
output(0, 52) <= input(19);
output(0, 53) <= input(20);
output(0, 54) <= input(21);
output(0, 55) <= input(22);
output(0, 56) <= input(23);
output(0, 57) <= input(24);
output(0, 58) <= input(25);
output(0, 59) <= input(26);
output(0, 60) <= input(27);
output(0, 61) <= input(28);
output(0, 62) <= input(29);
output(0, 63) <= input(30);
output(0, 64) <= input(34);
output(0, 65) <= input(32);
output(0, 66) <= input(0);
output(0, 67) <= input(1);
output(0, 68) <= input(2);
output(0, 69) <= input(3);
output(0, 70) <= input(4);
output(0, 71) <= input(5);
output(0, 72) <= input(6);
output(0, 73) <= input(7);
output(0, 74) <= input(8);
output(0, 75) <= input(9);
output(0, 76) <= input(10);
output(0, 77) <= input(11);
output(0, 78) <= input(12);
output(0, 79) <= input(13);
output(0, 80) <= input(35);
output(0, 81) <= input(33);
output(0, 82) <= input(16);
output(0, 83) <= input(17);
output(0, 84) <= input(18);
output(0, 85) <= input(19);
output(0, 86) <= input(20);
output(0, 87) <= input(21);
output(0, 88) <= input(22);
output(0, 89) <= input(23);
output(0, 90) <= input(24);
output(0, 91) <= input(25);
output(0, 92) <= input(26);
output(0, 93) <= input(27);
output(0, 94) <= input(28);
output(0, 95) <= input(29);
output(0, 96) <= input(36);
output(0, 97) <= input(34);
output(0, 98) <= input(32);
output(0, 99) <= input(0);
output(0, 100) <= input(1);
output(0, 101) <= input(2);
output(0, 102) <= input(3);
output(0, 103) <= input(4);
output(0, 104) <= input(5);
output(0, 105) <= input(6);
output(0, 106) <= input(7);
output(0, 107) <= input(8);
output(0, 108) <= input(9);
output(0, 109) <= input(10);
output(0, 110) <= input(11);
output(0, 111) <= input(12);
output(0, 112) <= input(36);
output(0, 113) <= input(34);
output(0, 114) <= input(32);
output(0, 115) <= input(0);
output(0, 116) <= input(1);
output(0, 117) <= input(2);
output(0, 118) <= input(3);
output(0, 119) <= input(4);
output(0, 120) <= input(5);
output(0, 121) <= input(6);
output(0, 122) <= input(7);
output(0, 123) <= input(8);
output(0, 124) <= input(9);
output(0, 125) <= input(10);
output(0, 126) <= input(11);
output(0, 127) <= input(12);
output(0, 128) <= input(37);
output(0, 129) <= input(35);
output(0, 130) <= input(33);
output(0, 131) <= input(16);
output(0, 132) <= input(17);
output(0, 133) <= input(18);
output(0, 134) <= input(19);
output(0, 135) <= input(20);
output(0, 136) <= input(21);
output(0, 137) <= input(22);
output(0, 138) <= input(23);
output(0, 139) <= input(24);
output(0, 140) <= input(25);
output(0, 141) <= input(26);
output(0, 142) <= input(27);
output(0, 143) <= input(28);
output(0, 144) <= input(38);
output(0, 145) <= input(36);
output(0, 146) <= input(34);
output(0, 147) <= input(32);
output(0, 148) <= input(0);
output(0, 149) <= input(1);
output(0, 150) <= input(2);
output(0, 151) <= input(3);
output(0, 152) <= input(4);
output(0, 153) <= input(5);
output(0, 154) <= input(6);
output(0, 155) <= input(7);
output(0, 156) <= input(8);
output(0, 157) <= input(9);
output(0, 158) <= input(10);
output(0, 159) <= input(11);
output(0, 160) <= input(39);
output(0, 161) <= input(37);
output(0, 162) <= input(35);
output(0, 163) <= input(33);
output(0, 164) <= input(16);
output(0, 165) <= input(17);
output(0, 166) <= input(18);
output(0, 167) <= input(19);
output(0, 168) <= input(20);
output(0, 169) <= input(21);
output(0, 170) <= input(22);
output(0, 171) <= input(23);
output(0, 172) <= input(24);
output(0, 173) <= input(25);
output(0, 174) <= input(26);
output(0, 175) <= input(27);
output(0, 176) <= input(40);
output(0, 177) <= input(38);
output(0, 178) <= input(36);
output(0, 179) <= input(34);
output(0, 180) <= input(32);
output(0, 181) <= input(0);
output(0, 182) <= input(1);
output(0, 183) <= input(2);
output(0, 184) <= input(3);
output(0, 185) <= input(4);
output(0, 186) <= input(5);
output(0, 187) <= input(6);
output(0, 188) <= input(7);
output(0, 189) <= input(8);
output(0, 190) <= input(9);
output(0, 191) <= input(10);
output(0, 192) <= input(41);
output(0, 193) <= input(39);
output(0, 194) <= input(37);
output(0, 195) <= input(35);
output(0, 196) <= input(33);
output(0, 197) <= input(16);
output(0, 198) <= input(17);
output(0, 199) <= input(18);
output(0, 200) <= input(19);
output(0, 201) <= input(20);
output(0, 202) <= input(21);
output(0, 203) <= input(22);
output(0, 204) <= input(23);
output(0, 205) <= input(24);
output(0, 206) <= input(25);
output(0, 207) <= input(26);
output(0, 208) <= input(42);
output(0, 209) <= input(40);
output(0, 210) <= input(38);
output(0, 211) <= input(36);
output(0, 212) <= input(34);
output(0, 213) <= input(32);
output(0, 214) <= input(0);
output(0, 215) <= input(1);
output(0, 216) <= input(2);
output(0, 217) <= input(3);
output(0, 218) <= input(4);
output(0, 219) <= input(5);
output(0, 220) <= input(6);
output(0, 221) <= input(7);
output(0, 222) <= input(8);
output(0, 223) <= input(9);
output(0, 224) <= input(43);
output(0, 225) <= input(41);
output(0, 226) <= input(39);
output(0, 227) <= input(37);
output(0, 228) <= input(35);
output(0, 229) <= input(33);
output(0, 230) <= input(16);
output(0, 231) <= input(17);
output(0, 232) <= input(18);
output(0, 233) <= input(19);
output(0, 234) <= input(20);
output(0, 235) <= input(21);
output(0, 236) <= input(22);
output(0, 237) <= input(23);
output(0, 238) <= input(24);
output(0, 239) <= input(25);
output(0, 240) <= input(43);
output(0, 241) <= input(41);
output(0, 242) <= input(39);
output(0, 243) <= input(37);
output(0, 244) <= input(35);
output(0, 245) <= input(33);
output(0, 246) <= input(16);
output(0, 247) <= input(17);
output(0, 248) <= input(18);
output(0, 249) <= input(19);
output(0, 250) <= input(20);
output(0, 251) <= input(21);
output(0, 252) <= input(22);
output(0, 253) <= input(23);
output(0, 254) <= input(24);
output(0, 255) <= input(25);
output(1, 0) <= input(44);
output(1, 1) <= input(1);
output(1, 2) <= input(2);
output(1, 3) <= input(3);
output(1, 4) <= input(4);
output(1, 5) <= input(5);
output(1, 6) <= input(6);
output(1, 7) <= input(7);
output(1, 8) <= input(8);
output(1, 9) <= input(9);
output(1, 10) <= input(10);
output(1, 11) <= input(11);
output(1, 12) <= input(12);
output(1, 13) <= input(13);
output(1, 14) <= input(14);
output(1, 15) <= input(15);
output(1, 16) <= input(45);
output(1, 17) <= input(17);
output(1, 18) <= input(18);
output(1, 19) <= input(19);
output(1, 20) <= input(20);
output(1, 21) <= input(21);
output(1, 22) <= input(22);
output(1, 23) <= input(23);
output(1, 24) <= input(24);
output(1, 25) <= input(25);
output(1, 26) <= input(26);
output(1, 27) <= input(27);
output(1, 28) <= input(28);
output(1, 29) <= input(29);
output(1, 30) <= input(30);
output(1, 31) <= input(31);
output(1, 32) <= input(46);
output(1, 33) <= input(44);
output(1, 34) <= input(1);
output(1, 35) <= input(2);
output(1, 36) <= input(3);
output(1, 37) <= input(4);
output(1, 38) <= input(5);
output(1, 39) <= input(6);
output(1, 40) <= input(7);
output(1, 41) <= input(8);
output(1, 42) <= input(9);
output(1, 43) <= input(10);
output(1, 44) <= input(11);
output(1, 45) <= input(12);
output(1, 46) <= input(13);
output(1, 47) <= input(14);
output(1, 48) <= input(46);
output(1, 49) <= input(44);
output(1, 50) <= input(1);
output(1, 51) <= input(2);
output(1, 52) <= input(3);
output(1, 53) <= input(4);
output(1, 54) <= input(5);
output(1, 55) <= input(6);
output(1, 56) <= input(7);
output(1, 57) <= input(8);
output(1, 58) <= input(9);
output(1, 59) <= input(10);
output(1, 60) <= input(11);
output(1, 61) <= input(12);
output(1, 62) <= input(13);
output(1, 63) <= input(14);
output(1, 64) <= input(47);
output(1, 65) <= input(45);
output(1, 66) <= input(17);
output(1, 67) <= input(18);
output(1, 68) <= input(19);
output(1, 69) <= input(20);
output(1, 70) <= input(21);
output(1, 71) <= input(22);
output(1, 72) <= input(23);
output(1, 73) <= input(24);
output(1, 74) <= input(25);
output(1, 75) <= input(26);
output(1, 76) <= input(27);
output(1, 77) <= input(28);
output(1, 78) <= input(29);
output(1, 79) <= input(30);
output(1, 80) <= input(48);
output(1, 81) <= input(46);
output(1, 82) <= input(44);
output(1, 83) <= input(1);
output(1, 84) <= input(2);
output(1, 85) <= input(3);
output(1, 86) <= input(4);
output(1, 87) <= input(5);
output(1, 88) <= input(6);
output(1, 89) <= input(7);
output(1, 90) <= input(8);
output(1, 91) <= input(9);
output(1, 92) <= input(10);
output(1, 93) <= input(11);
output(1, 94) <= input(12);
output(1, 95) <= input(13);
output(1, 96) <= input(49);
output(1, 97) <= input(47);
output(1, 98) <= input(45);
output(1, 99) <= input(17);
output(1, 100) <= input(18);
output(1, 101) <= input(19);
output(1, 102) <= input(20);
output(1, 103) <= input(21);
output(1, 104) <= input(22);
output(1, 105) <= input(23);
output(1, 106) <= input(24);
output(1, 107) <= input(25);
output(1, 108) <= input(26);
output(1, 109) <= input(27);
output(1, 110) <= input(28);
output(1, 111) <= input(29);
output(1, 112) <= input(49);
output(1, 113) <= input(47);
output(1, 114) <= input(45);
output(1, 115) <= input(17);
output(1, 116) <= input(18);
output(1, 117) <= input(19);
output(1, 118) <= input(20);
output(1, 119) <= input(21);
output(1, 120) <= input(22);
output(1, 121) <= input(23);
output(1, 122) <= input(24);
output(1, 123) <= input(25);
output(1, 124) <= input(26);
output(1, 125) <= input(27);
output(1, 126) <= input(28);
output(1, 127) <= input(29);
output(1, 128) <= input(50);
output(1, 129) <= input(48);
output(1, 130) <= input(46);
output(1, 131) <= input(44);
output(1, 132) <= input(1);
output(1, 133) <= input(2);
output(1, 134) <= input(3);
output(1, 135) <= input(4);
output(1, 136) <= input(5);
output(1, 137) <= input(6);
output(1, 138) <= input(7);
output(1, 139) <= input(8);
output(1, 140) <= input(9);
output(1, 141) <= input(10);
output(1, 142) <= input(11);
output(1, 143) <= input(12);
output(1, 144) <= input(51);
output(1, 145) <= input(49);
output(1, 146) <= input(47);
output(1, 147) <= input(45);
output(1, 148) <= input(17);
output(1, 149) <= input(18);
output(1, 150) <= input(19);
output(1, 151) <= input(20);
output(1, 152) <= input(21);
output(1, 153) <= input(22);
output(1, 154) <= input(23);
output(1, 155) <= input(24);
output(1, 156) <= input(25);
output(1, 157) <= input(26);
output(1, 158) <= input(27);
output(1, 159) <= input(28);
output(1, 160) <= input(52);
output(1, 161) <= input(50);
output(1, 162) <= input(48);
output(1, 163) <= input(46);
output(1, 164) <= input(44);
output(1, 165) <= input(1);
output(1, 166) <= input(2);
output(1, 167) <= input(3);
output(1, 168) <= input(4);
output(1, 169) <= input(5);
output(1, 170) <= input(6);
output(1, 171) <= input(7);
output(1, 172) <= input(8);
output(1, 173) <= input(9);
output(1, 174) <= input(10);
output(1, 175) <= input(11);
output(1, 176) <= input(52);
output(1, 177) <= input(50);
output(1, 178) <= input(48);
output(1, 179) <= input(46);
output(1, 180) <= input(44);
output(1, 181) <= input(1);
output(1, 182) <= input(2);
output(1, 183) <= input(3);
output(1, 184) <= input(4);
output(1, 185) <= input(5);
output(1, 186) <= input(6);
output(1, 187) <= input(7);
output(1, 188) <= input(8);
output(1, 189) <= input(9);
output(1, 190) <= input(10);
output(1, 191) <= input(11);
output(1, 192) <= input(53);
output(1, 193) <= input(51);
output(1, 194) <= input(49);
output(1, 195) <= input(47);
output(1, 196) <= input(45);
output(1, 197) <= input(17);
output(1, 198) <= input(18);
output(1, 199) <= input(19);
output(1, 200) <= input(20);
output(1, 201) <= input(21);
output(1, 202) <= input(22);
output(1, 203) <= input(23);
output(1, 204) <= input(24);
output(1, 205) <= input(25);
output(1, 206) <= input(26);
output(1, 207) <= input(27);
output(1, 208) <= input(54);
output(1, 209) <= input(52);
output(1, 210) <= input(50);
output(1, 211) <= input(48);
output(1, 212) <= input(46);
output(1, 213) <= input(44);
output(1, 214) <= input(1);
output(1, 215) <= input(2);
output(1, 216) <= input(3);
output(1, 217) <= input(4);
output(1, 218) <= input(5);
output(1, 219) <= input(6);
output(1, 220) <= input(7);
output(1, 221) <= input(8);
output(1, 222) <= input(9);
output(1, 223) <= input(10);
output(1, 224) <= input(55);
output(1, 225) <= input(53);
output(1, 226) <= input(51);
output(1, 227) <= input(49);
output(1, 228) <= input(47);
output(1, 229) <= input(45);
output(1, 230) <= input(17);
output(1, 231) <= input(18);
output(1, 232) <= input(19);
output(1, 233) <= input(20);
output(1, 234) <= input(21);
output(1, 235) <= input(22);
output(1, 236) <= input(23);
output(1, 237) <= input(24);
output(1, 238) <= input(25);
output(1, 239) <= input(26);
output(1, 240) <= input(55);
output(1, 241) <= input(53);
output(1, 242) <= input(51);
output(1, 243) <= input(49);
output(1, 244) <= input(47);
output(1, 245) <= input(45);
output(1, 246) <= input(17);
output(1, 247) <= input(18);
output(1, 248) <= input(19);
output(1, 249) <= input(20);
output(1, 250) <= input(21);
output(1, 251) <= input(22);
output(1, 252) <= input(23);
output(1, 253) <= input(24);
output(1, 254) <= input(25);
output(1, 255) <= input(26);
output(2, 0) <= input(44);
output(2, 1) <= input(1);
output(2, 2) <= input(2);
output(2, 3) <= input(3);
output(2, 4) <= input(4);
output(2, 5) <= input(5);
output(2, 6) <= input(6);
output(2, 7) <= input(7);
output(2, 8) <= input(8);
output(2, 9) <= input(9);
output(2, 10) <= input(10);
output(2, 11) <= input(11);
output(2, 12) <= input(12);
output(2, 13) <= input(13);
output(2, 14) <= input(14);
output(2, 15) <= input(15);
output(2, 16) <= input(45);
output(2, 17) <= input(17);
output(2, 18) <= input(18);
output(2, 19) <= input(19);
output(2, 20) <= input(20);
output(2, 21) <= input(21);
output(2, 22) <= input(22);
output(2, 23) <= input(23);
output(2, 24) <= input(24);
output(2, 25) <= input(25);
output(2, 26) <= input(26);
output(2, 27) <= input(27);
output(2, 28) <= input(28);
output(2, 29) <= input(29);
output(2, 30) <= input(30);
output(2, 31) <= input(31);
output(2, 32) <= input(45);
output(2, 33) <= input(17);
output(2, 34) <= input(18);
output(2, 35) <= input(19);
output(2, 36) <= input(20);
output(2, 37) <= input(21);
output(2, 38) <= input(22);
output(2, 39) <= input(23);
output(2, 40) <= input(24);
output(2, 41) <= input(25);
output(2, 42) <= input(26);
output(2, 43) <= input(27);
output(2, 44) <= input(28);
output(2, 45) <= input(29);
output(2, 46) <= input(30);
output(2, 47) <= input(31);
output(2, 48) <= input(56);
output(2, 49) <= input(44);
output(2, 50) <= input(1);
output(2, 51) <= input(2);
output(2, 52) <= input(3);
output(2, 53) <= input(4);
output(2, 54) <= input(5);
output(2, 55) <= input(6);
output(2, 56) <= input(7);
output(2, 57) <= input(8);
output(2, 58) <= input(9);
output(2, 59) <= input(10);
output(2, 60) <= input(11);
output(2, 61) <= input(12);
output(2, 62) <= input(13);
output(2, 63) <= input(14);
output(2, 64) <= input(57);
output(2, 65) <= input(45);
output(2, 66) <= input(17);
output(2, 67) <= input(18);
output(2, 68) <= input(19);
output(2, 69) <= input(20);
output(2, 70) <= input(21);
output(2, 71) <= input(22);
output(2, 72) <= input(23);
output(2, 73) <= input(24);
output(2, 74) <= input(25);
output(2, 75) <= input(26);
output(2, 76) <= input(27);
output(2, 77) <= input(28);
output(2, 78) <= input(29);
output(2, 79) <= input(30);
output(2, 80) <= input(57);
output(2, 81) <= input(45);
output(2, 82) <= input(17);
output(2, 83) <= input(18);
output(2, 84) <= input(19);
output(2, 85) <= input(20);
output(2, 86) <= input(21);
output(2, 87) <= input(22);
output(2, 88) <= input(23);
output(2, 89) <= input(24);
output(2, 90) <= input(25);
output(2, 91) <= input(26);
output(2, 92) <= input(27);
output(2, 93) <= input(28);
output(2, 94) <= input(29);
output(2, 95) <= input(30);
output(2, 96) <= input(58);
output(2, 97) <= input(56);
output(2, 98) <= input(44);
output(2, 99) <= input(1);
output(2, 100) <= input(2);
output(2, 101) <= input(3);
output(2, 102) <= input(4);
output(2, 103) <= input(5);
output(2, 104) <= input(6);
output(2, 105) <= input(7);
output(2, 106) <= input(8);
output(2, 107) <= input(9);
output(2, 108) <= input(10);
output(2, 109) <= input(11);
output(2, 110) <= input(12);
output(2, 111) <= input(13);
output(2, 112) <= input(58);
output(2, 113) <= input(56);
output(2, 114) <= input(44);
output(2, 115) <= input(1);
output(2, 116) <= input(2);
output(2, 117) <= input(3);
output(2, 118) <= input(4);
output(2, 119) <= input(5);
output(2, 120) <= input(6);
output(2, 121) <= input(7);
output(2, 122) <= input(8);
output(2, 123) <= input(9);
output(2, 124) <= input(10);
output(2, 125) <= input(11);
output(2, 126) <= input(12);
output(2, 127) <= input(13);
output(2, 128) <= input(59);
output(2, 129) <= input(57);
output(2, 130) <= input(45);
output(2, 131) <= input(17);
output(2, 132) <= input(18);
output(2, 133) <= input(19);
output(2, 134) <= input(20);
output(2, 135) <= input(21);
output(2, 136) <= input(22);
output(2, 137) <= input(23);
output(2, 138) <= input(24);
output(2, 139) <= input(25);
output(2, 140) <= input(26);
output(2, 141) <= input(27);
output(2, 142) <= input(28);
output(2, 143) <= input(29);
output(2, 144) <= input(60);
output(2, 145) <= input(58);
output(2, 146) <= input(56);
output(2, 147) <= input(44);
output(2, 148) <= input(1);
output(2, 149) <= input(2);
output(2, 150) <= input(3);
output(2, 151) <= input(4);
output(2, 152) <= input(5);
output(2, 153) <= input(6);
output(2, 154) <= input(7);
output(2, 155) <= input(8);
output(2, 156) <= input(9);
output(2, 157) <= input(10);
output(2, 158) <= input(11);
output(2, 159) <= input(12);
output(2, 160) <= input(60);
output(2, 161) <= input(58);
output(2, 162) <= input(56);
output(2, 163) <= input(44);
output(2, 164) <= input(1);
output(2, 165) <= input(2);
output(2, 166) <= input(3);
output(2, 167) <= input(4);
output(2, 168) <= input(5);
output(2, 169) <= input(6);
output(2, 170) <= input(7);
output(2, 171) <= input(8);
output(2, 172) <= input(9);
output(2, 173) <= input(10);
output(2, 174) <= input(11);
output(2, 175) <= input(12);
output(2, 176) <= input(61);
output(2, 177) <= input(59);
output(2, 178) <= input(57);
output(2, 179) <= input(45);
output(2, 180) <= input(17);
output(2, 181) <= input(18);
output(2, 182) <= input(19);
output(2, 183) <= input(20);
output(2, 184) <= input(21);
output(2, 185) <= input(22);
output(2, 186) <= input(23);
output(2, 187) <= input(24);
output(2, 188) <= input(25);
output(2, 189) <= input(26);
output(2, 190) <= input(27);
output(2, 191) <= input(28);
output(2, 192) <= input(62);
output(2, 193) <= input(60);
output(2, 194) <= input(58);
output(2, 195) <= input(56);
output(2, 196) <= input(44);
output(2, 197) <= input(1);
output(2, 198) <= input(2);
output(2, 199) <= input(3);
output(2, 200) <= input(4);
output(2, 201) <= input(5);
output(2, 202) <= input(6);
output(2, 203) <= input(7);
output(2, 204) <= input(8);
output(2, 205) <= input(9);
output(2, 206) <= input(10);
output(2, 207) <= input(11);
output(2, 208) <= input(62);
output(2, 209) <= input(60);
output(2, 210) <= input(58);
output(2, 211) <= input(56);
output(2, 212) <= input(44);
output(2, 213) <= input(1);
output(2, 214) <= input(2);
output(2, 215) <= input(3);
output(2, 216) <= input(4);
output(2, 217) <= input(5);
output(2, 218) <= input(6);
output(2, 219) <= input(7);
output(2, 220) <= input(8);
output(2, 221) <= input(9);
output(2, 222) <= input(10);
output(2, 223) <= input(11);
output(2, 224) <= input(63);
output(2, 225) <= input(61);
output(2, 226) <= input(59);
output(2, 227) <= input(57);
output(2, 228) <= input(45);
output(2, 229) <= input(17);
output(2, 230) <= input(18);
output(2, 231) <= input(19);
output(2, 232) <= input(20);
output(2, 233) <= input(21);
output(2, 234) <= input(22);
output(2, 235) <= input(23);
output(2, 236) <= input(24);
output(2, 237) <= input(25);
output(2, 238) <= input(26);
output(2, 239) <= input(27);
output(2, 240) <= input(63);
output(2, 241) <= input(61);
output(2, 242) <= input(59);
output(2, 243) <= input(57);
output(2, 244) <= input(45);
output(2, 245) <= input(17);
output(2, 246) <= input(18);
output(2, 247) <= input(19);
output(2, 248) <= input(20);
output(2, 249) <= input(21);
output(2, 250) <= input(22);
output(2, 251) <= input(23);
output(2, 252) <= input(24);
output(2, 253) <= input(25);
output(2, 254) <= input(26);
output(2, 255) <= input(27);
when "1100" =>
output(0, 0) <= input(0);
output(0, 1) <= input(1);
output(0, 2) <= input(2);
output(0, 3) <= input(3);
output(0, 4) <= input(4);
output(0, 5) <= input(5);
output(0, 6) <= input(6);
output(0, 7) <= input(7);
output(0, 8) <= input(8);
output(0, 9) <= input(9);
output(0, 10) <= input(10);
output(0, 11) <= input(11);
output(0, 12) <= input(12);
output(0, 13) <= input(13);
output(0, 14) <= input(14);
output(0, 15) <= input(15);
output(0, 16) <= input(0);
output(0, 17) <= input(1);
output(0, 18) <= input(2);
output(0, 19) <= input(3);
output(0, 20) <= input(4);
output(0, 21) <= input(5);
output(0, 22) <= input(6);
output(0, 23) <= input(7);
output(0, 24) <= input(8);
output(0, 25) <= input(9);
output(0, 26) <= input(10);
output(0, 27) <= input(11);
output(0, 28) <= input(12);
output(0, 29) <= input(13);
output(0, 30) <= input(14);
output(0, 31) <= input(15);
output(0, 32) <= input(16);
output(0, 33) <= input(17);
output(0, 34) <= input(18);
output(0, 35) <= input(19);
output(0, 36) <= input(20);
output(0, 37) <= input(21);
output(0, 38) <= input(22);
output(0, 39) <= input(23);
output(0, 40) <= input(24);
output(0, 41) <= input(25);
output(0, 42) <= input(26);
output(0, 43) <= input(27);
output(0, 44) <= input(28);
output(0, 45) <= input(29);
output(0, 46) <= input(30);
output(0, 47) <= input(31);
output(0, 48) <= input(16);
output(0, 49) <= input(17);
output(0, 50) <= input(18);
output(0, 51) <= input(19);
output(0, 52) <= input(20);
output(0, 53) <= input(21);
output(0, 54) <= input(22);
output(0, 55) <= input(23);
output(0, 56) <= input(24);
output(0, 57) <= input(25);
output(0, 58) <= input(26);
output(0, 59) <= input(27);
output(0, 60) <= input(28);
output(0, 61) <= input(29);
output(0, 62) <= input(30);
output(0, 63) <= input(31);
output(0, 64) <= input(32);
output(0, 65) <= input(0);
output(0, 66) <= input(1);
output(0, 67) <= input(2);
output(0, 68) <= input(3);
output(0, 69) <= input(4);
output(0, 70) <= input(5);
output(0, 71) <= input(6);
output(0, 72) <= input(7);
output(0, 73) <= input(8);
output(0, 74) <= input(9);
output(0, 75) <= input(10);
output(0, 76) <= input(11);
output(0, 77) <= input(12);
output(0, 78) <= input(13);
output(0, 79) <= input(14);
output(0, 80) <= input(32);
output(0, 81) <= input(0);
output(0, 82) <= input(1);
output(0, 83) <= input(2);
output(0, 84) <= input(3);
output(0, 85) <= input(4);
output(0, 86) <= input(5);
output(0, 87) <= input(6);
output(0, 88) <= input(7);
output(0, 89) <= input(8);
output(0, 90) <= input(9);
output(0, 91) <= input(10);
output(0, 92) <= input(11);
output(0, 93) <= input(12);
output(0, 94) <= input(13);
output(0, 95) <= input(14);
output(0, 96) <= input(33);
output(0, 97) <= input(16);
output(0, 98) <= input(17);
output(0, 99) <= input(18);
output(0, 100) <= input(19);
output(0, 101) <= input(20);
output(0, 102) <= input(21);
output(0, 103) <= input(22);
output(0, 104) <= input(23);
output(0, 105) <= input(24);
output(0, 106) <= input(25);
output(0, 107) <= input(26);
output(0, 108) <= input(27);
output(0, 109) <= input(28);
output(0, 110) <= input(29);
output(0, 111) <= input(30);
output(0, 112) <= input(33);
output(0, 113) <= input(16);
output(0, 114) <= input(17);
output(0, 115) <= input(18);
output(0, 116) <= input(19);
output(0, 117) <= input(20);
output(0, 118) <= input(21);
output(0, 119) <= input(22);
output(0, 120) <= input(23);
output(0, 121) <= input(24);
output(0, 122) <= input(25);
output(0, 123) <= input(26);
output(0, 124) <= input(27);
output(0, 125) <= input(28);
output(0, 126) <= input(29);
output(0, 127) <= input(30);
output(0, 128) <= input(34);
output(0, 129) <= input(32);
output(0, 130) <= input(0);
output(0, 131) <= input(1);
output(0, 132) <= input(2);
output(0, 133) <= input(3);
output(0, 134) <= input(4);
output(0, 135) <= input(5);
output(0, 136) <= input(6);
output(0, 137) <= input(7);
output(0, 138) <= input(8);
output(0, 139) <= input(9);
output(0, 140) <= input(10);
output(0, 141) <= input(11);
output(0, 142) <= input(12);
output(0, 143) <= input(13);
output(0, 144) <= input(34);
output(0, 145) <= input(32);
output(0, 146) <= input(0);
output(0, 147) <= input(1);
output(0, 148) <= input(2);
output(0, 149) <= input(3);
output(0, 150) <= input(4);
output(0, 151) <= input(5);
output(0, 152) <= input(6);
output(0, 153) <= input(7);
output(0, 154) <= input(8);
output(0, 155) <= input(9);
output(0, 156) <= input(10);
output(0, 157) <= input(11);
output(0, 158) <= input(12);
output(0, 159) <= input(13);
output(0, 160) <= input(35);
output(0, 161) <= input(33);
output(0, 162) <= input(16);
output(0, 163) <= input(17);
output(0, 164) <= input(18);
output(0, 165) <= input(19);
output(0, 166) <= input(20);
output(0, 167) <= input(21);
output(0, 168) <= input(22);
output(0, 169) <= input(23);
output(0, 170) <= input(24);
output(0, 171) <= input(25);
output(0, 172) <= input(26);
output(0, 173) <= input(27);
output(0, 174) <= input(28);
output(0, 175) <= input(29);
output(0, 176) <= input(35);
output(0, 177) <= input(33);
output(0, 178) <= input(16);
output(0, 179) <= input(17);
output(0, 180) <= input(18);
output(0, 181) <= input(19);
output(0, 182) <= input(20);
output(0, 183) <= input(21);
output(0, 184) <= input(22);
output(0, 185) <= input(23);
output(0, 186) <= input(24);
output(0, 187) <= input(25);
output(0, 188) <= input(26);
output(0, 189) <= input(27);
output(0, 190) <= input(28);
output(0, 191) <= input(29);
output(0, 192) <= input(36);
output(0, 193) <= input(34);
output(0, 194) <= input(32);
output(0, 195) <= input(0);
output(0, 196) <= input(1);
output(0, 197) <= input(2);
output(0, 198) <= input(3);
output(0, 199) <= input(4);
output(0, 200) <= input(5);
output(0, 201) <= input(6);
output(0, 202) <= input(7);
output(0, 203) <= input(8);
output(0, 204) <= input(9);
output(0, 205) <= input(10);
output(0, 206) <= input(11);
output(0, 207) <= input(12);
output(0, 208) <= input(36);
output(0, 209) <= input(34);
output(0, 210) <= input(32);
output(0, 211) <= input(0);
output(0, 212) <= input(1);
output(0, 213) <= input(2);
output(0, 214) <= input(3);
output(0, 215) <= input(4);
output(0, 216) <= input(5);
output(0, 217) <= input(6);
output(0, 218) <= input(7);
output(0, 219) <= input(8);
output(0, 220) <= input(9);
output(0, 221) <= input(10);
output(0, 222) <= input(11);
output(0, 223) <= input(12);
output(0, 224) <= input(37);
output(0, 225) <= input(35);
output(0, 226) <= input(33);
output(0, 227) <= input(16);
output(0, 228) <= input(17);
output(0, 229) <= input(18);
output(0, 230) <= input(19);
output(0, 231) <= input(20);
output(0, 232) <= input(21);
output(0, 233) <= input(22);
output(0, 234) <= input(23);
output(0, 235) <= input(24);
output(0, 236) <= input(25);
output(0, 237) <= input(26);
output(0, 238) <= input(27);
output(0, 239) <= input(28);
output(0, 240) <= input(37);
output(0, 241) <= input(35);
output(0, 242) <= input(33);
output(0, 243) <= input(16);
output(0, 244) <= input(17);
output(0, 245) <= input(18);
output(0, 246) <= input(19);
output(0, 247) <= input(20);
output(0, 248) <= input(21);
output(0, 249) <= input(22);
output(0, 250) <= input(23);
output(0, 251) <= input(24);
output(0, 252) <= input(25);
output(0, 253) <= input(26);
output(0, 254) <= input(27);
output(0, 255) <= input(28);
output(1, 0) <= input(38);
output(1, 1) <= input(1);
output(1, 2) <= input(2);
output(1, 3) <= input(3);
output(1, 4) <= input(4);
output(1, 5) <= input(5);
output(1, 6) <= input(6);
output(1, 7) <= input(7);
output(1, 8) <= input(8);
output(1, 9) <= input(9);
output(1, 10) <= input(10);
output(1, 11) <= input(11);
output(1, 12) <= input(12);
output(1, 13) <= input(13);
output(1, 14) <= input(14);
output(1, 15) <= input(15);
output(1, 16) <= input(38);
output(1, 17) <= input(1);
output(1, 18) <= input(2);
output(1, 19) <= input(3);
output(1, 20) <= input(4);
output(1, 21) <= input(5);
output(1, 22) <= input(6);
output(1, 23) <= input(7);
output(1, 24) <= input(8);
output(1, 25) <= input(9);
output(1, 26) <= input(10);
output(1, 27) <= input(11);
output(1, 28) <= input(12);
output(1, 29) <= input(13);
output(1, 30) <= input(14);
output(1, 31) <= input(15);
output(1, 32) <= input(39);
output(1, 33) <= input(17);
output(1, 34) <= input(18);
output(1, 35) <= input(19);
output(1, 36) <= input(20);
output(1, 37) <= input(21);
output(1, 38) <= input(22);
output(1, 39) <= input(23);
output(1, 40) <= input(24);
output(1, 41) <= input(25);
output(1, 42) <= input(26);
output(1, 43) <= input(27);
output(1, 44) <= input(28);
output(1, 45) <= input(29);
output(1, 46) <= input(30);
output(1, 47) <= input(31);
output(1, 48) <= input(39);
output(1, 49) <= input(17);
output(1, 50) <= input(18);
output(1, 51) <= input(19);
output(1, 52) <= input(20);
output(1, 53) <= input(21);
output(1, 54) <= input(22);
output(1, 55) <= input(23);
output(1, 56) <= input(24);
output(1, 57) <= input(25);
output(1, 58) <= input(26);
output(1, 59) <= input(27);
output(1, 60) <= input(28);
output(1, 61) <= input(29);
output(1, 62) <= input(30);
output(1, 63) <= input(31);
output(1, 64) <= input(39);
output(1, 65) <= input(17);
output(1, 66) <= input(18);
output(1, 67) <= input(19);
output(1, 68) <= input(20);
output(1, 69) <= input(21);
output(1, 70) <= input(22);
output(1, 71) <= input(23);
output(1, 72) <= input(24);
output(1, 73) <= input(25);
output(1, 74) <= input(26);
output(1, 75) <= input(27);
output(1, 76) <= input(28);
output(1, 77) <= input(29);
output(1, 78) <= input(30);
output(1, 79) <= input(31);
output(1, 80) <= input(40);
output(1, 81) <= input(38);
output(1, 82) <= input(1);
output(1, 83) <= input(2);
output(1, 84) <= input(3);
output(1, 85) <= input(4);
output(1, 86) <= input(5);
output(1, 87) <= input(6);
output(1, 88) <= input(7);
output(1, 89) <= input(8);
output(1, 90) <= input(9);
output(1, 91) <= input(10);
output(1, 92) <= input(11);
output(1, 93) <= input(12);
output(1, 94) <= input(13);
output(1, 95) <= input(14);
output(1, 96) <= input(40);
output(1, 97) <= input(38);
output(1, 98) <= input(1);
output(1, 99) <= input(2);
output(1, 100) <= input(3);
output(1, 101) <= input(4);
output(1, 102) <= input(5);
output(1, 103) <= input(6);
output(1, 104) <= input(7);
output(1, 105) <= input(8);
output(1, 106) <= input(9);
output(1, 107) <= input(10);
output(1, 108) <= input(11);
output(1, 109) <= input(12);
output(1, 110) <= input(13);
output(1, 111) <= input(14);
output(1, 112) <= input(40);
output(1, 113) <= input(38);
output(1, 114) <= input(1);
output(1, 115) <= input(2);
output(1, 116) <= input(3);
output(1, 117) <= input(4);
output(1, 118) <= input(5);
output(1, 119) <= input(6);
output(1, 120) <= input(7);
output(1, 121) <= input(8);
output(1, 122) <= input(9);
output(1, 123) <= input(10);
output(1, 124) <= input(11);
output(1, 125) <= input(12);
output(1, 126) <= input(13);
output(1, 127) <= input(14);
output(1, 128) <= input(41);
output(1, 129) <= input(39);
output(1, 130) <= input(17);
output(1, 131) <= input(18);
output(1, 132) <= input(19);
output(1, 133) <= input(20);
output(1, 134) <= input(21);
output(1, 135) <= input(22);
output(1, 136) <= input(23);
output(1, 137) <= input(24);
output(1, 138) <= input(25);
output(1, 139) <= input(26);
output(1, 140) <= input(27);
output(1, 141) <= input(28);
output(1, 142) <= input(29);
output(1, 143) <= input(30);
output(1, 144) <= input(41);
output(1, 145) <= input(39);
output(1, 146) <= input(17);
output(1, 147) <= input(18);
output(1, 148) <= input(19);
output(1, 149) <= input(20);
output(1, 150) <= input(21);
output(1, 151) <= input(22);
output(1, 152) <= input(23);
output(1, 153) <= input(24);
output(1, 154) <= input(25);
output(1, 155) <= input(26);
output(1, 156) <= input(27);
output(1, 157) <= input(28);
output(1, 158) <= input(29);
output(1, 159) <= input(30);
output(1, 160) <= input(42);
output(1, 161) <= input(40);
output(1, 162) <= input(38);
output(1, 163) <= input(1);
output(1, 164) <= input(2);
output(1, 165) <= input(3);
output(1, 166) <= input(4);
output(1, 167) <= input(5);
output(1, 168) <= input(6);
output(1, 169) <= input(7);
output(1, 170) <= input(8);
output(1, 171) <= input(9);
output(1, 172) <= input(10);
output(1, 173) <= input(11);
output(1, 174) <= input(12);
output(1, 175) <= input(13);
output(1, 176) <= input(42);
output(1, 177) <= input(40);
output(1, 178) <= input(38);
output(1, 179) <= input(1);
output(1, 180) <= input(2);
output(1, 181) <= input(3);
output(1, 182) <= input(4);
output(1, 183) <= input(5);
output(1, 184) <= input(6);
output(1, 185) <= input(7);
output(1, 186) <= input(8);
output(1, 187) <= input(9);
output(1, 188) <= input(10);
output(1, 189) <= input(11);
output(1, 190) <= input(12);
output(1, 191) <= input(13);
output(1, 192) <= input(42);
output(1, 193) <= input(40);
output(1, 194) <= input(38);
output(1, 195) <= input(1);
output(1, 196) <= input(2);
output(1, 197) <= input(3);
output(1, 198) <= input(4);
output(1, 199) <= input(5);
output(1, 200) <= input(6);
output(1, 201) <= input(7);
output(1, 202) <= input(8);
output(1, 203) <= input(9);
output(1, 204) <= input(10);
output(1, 205) <= input(11);
output(1, 206) <= input(12);
output(1, 207) <= input(13);
output(1, 208) <= input(43);
output(1, 209) <= input(41);
output(1, 210) <= input(39);
output(1, 211) <= input(17);
output(1, 212) <= input(18);
output(1, 213) <= input(19);
output(1, 214) <= input(20);
output(1, 215) <= input(21);
output(1, 216) <= input(22);
output(1, 217) <= input(23);
output(1, 218) <= input(24);
output(1, 219) <= input(25);
output(1, 220) <= input(26);
output(1, 221) <= input(27);
output(1, 222) <= input(28);
output(1, 223) <= input(29);
output(1, 224) <= input(43);
output(1, 225) <= input(41);
output(1, 226) <= input(39);
output(1, 227) <= input(17);
output(1, 228) <= input(18);
output(1, 229) <= input(19);
output(1, 230) <= input(20);
output(1, 231) <= input(21);
output(1, 232) <= input(22);
output(1, 233) <= input(23);
output(1, 234) <= input(24);
output(1, 235) <= input(25);
output(1, 236) <= input(26);
output(1, 237) <= input(27);
output(1, 238) <= input(28);
output(1, 239) <= input(29);
output(1, 240) <= input(43);
output(1, 241) <= input(41);
output(1, 242) <= input(39);
output(1, 243) <= input(17);
output(1, 244) <= input(18);
output(1, 245) <= input(19);
output(1, 246) <= input(20);
output(1, 247) <= input(21);
output(1, 248) <= input(22);
output(1, 249) <= input(23);
output(1, 250) <= input(24);
output(1, 251) <= input(25);
output(1, 252) <= input(26);
output(1, 253) <= input(27);
output(1, 254) <= input(28);
output(1, 255) <= input(29);
output(2, 0) <= input(44);
output(2, 1) <= input(1);
output(2, 2) <= input(2);
output(2, 3) <= input(3);
output(2, 4) <= input(4);
output(2, 5) <= input(5);
output(2, 6) <= input(6);
output(2, 7) <= input(7);
output(2, 8) <= input(8);
output(2, 9) <= input(9);
output(2, 10) <= input(10);
output(2, 11) <= input(11);
output(2, 12) <= input(12);
output(2, 13) <= input(13);
output(2, 14) <= input(14);
output(2, 15) <= input(15);
output(2, 16) <= input(44);
output(2, 17) <= input(1);
output(2, 18) <= input(2);
output(2, 19) <= input(3);
output(2, 20) <= input(4);
output(2, 21) <= input(5);
output(2, 22) <= input(6);
output(2, 23) <= input(7);
output(2, 24) <= input(8);
output(2, 25) <= input(9);
output(2, 26) <= input(10);
output(2, 27) <= input(11);
output(2, 28) <= input(12);
output(2, 29) <= input(13);
output(2, 30) <= input(14);
output(2, 31) <= input(15);
output(2, 32) <= input(44);
output(2, 33) <= input(1);
output(2, 34) <= input(2);
output(2, 35) <= input(3);
output(2, 36) <= input(4);
output(2, 37) <= input(5);
output(2, 38) <= input(6);
output(2, 39) <= input(7);
output(2, 40) <= input(8);
output(2, 41) <= input(9);
output(2, 42) <= input(10);
output(2, 43) <= input(11);
output(2, 44) <= input(12);
output(2, 45) <= input(13);
output(2, 46) <= input(14);
output(2, 47) <= input(15);
output(2, 48) <= input(44);
output(2, 49) <= input(1);
output(2, 50) <= input(2);
output(2, 51) <= input(3);
output(2, 52) <= input(4);
output(2, 53) <= input(5);
output(2, 54) <= input(6);
output(2, 55) <= input(7);
output(2, 56) <= input(8);
output(2, 57) <= input(9);
output(2, 58) <= input(10);
output(2, 59) <= input(11);
output(2, 60) <= input(12);
output(2, 61) <= input(13);
output(2, 62) <= input(14);
output(2, 63) <= input(15);
output(2, 64) <= input(45);
output(2, 65) <= input(17);
output(2, 66) <= input(18);
output(2, 67) <= input(19);
output(2, 68) <= input(20);
output(2, 69) <= input(21);
output(2, 70) <= input(22);
output(2, 71) <= input(23);
output(2, 72) <= input(24);
output(2, 73) <= input(25);
output(2, 74) <= input(26);
output(2, 75) <= input(27);
output(2, 76) <= input(28);
output(2, 77) <= input(29);
output(2, 78) <= input(30);
output(2, 79) <= input(31);
output(2, 80) <= input(45);
output(2, 81) <= input(17);
output(2, 82) <= input(18);
output(2, 83) <= input(19);
output(2, 84) <= input(20);
output(2, 85) <= input(21);
output(2, 86) <= input(22);
output(2, 87) <= input(23);
output(2, 88) <= input(24);
output(2, 89) <= input(25);
output(2, 90) <= input(26);
output(2, 91) <= input(27);
output(2, 92) <= input(28);
output(2, 93) <= input(29);
output(2, 94) <= input(30);
output(2, 95) <= input(31);
output(2, 96) <= input(45);
output(2, 97) <= input(17);
output(2, 98) <= input(18);
output(2, 99) <= input(19);
output(2, 100) <= input(20);
output(2, 101) <= input(21);
output(2, 102) <= input(22);
output(2, 103) <= input(23);
output(2, 104) <= input(24);
output(2, 105) <= input(25);
output(2, 106) <= input(26);
output(2, 107) <= input(27);
output(2, 108) <= input(28);
output(2, 109) <= input(29);
output(2, 110) <= input(30);
output(2, 111) <= input(31);
output(2, 112) <= input(45);
output(2, 113) <= input(17);
output(2, 114) <= input(18);
output(2, 115) <= input(19);
output(2, 116) <= input(20);
output(2, 117) <= input(21);
output(2, 118) <= input(22);
output(2, 119) <= input(23);
output(2, 120) <= input(24);
output(2, 121) <= input(25);
output(2, 122) <= input(26);
output(2, 123) <= input(27);
output(2, 124) <= input(28);
output(2, 125) <= input(29);
output(2, 126) <= input(30);
output(2, 127) <= input(31);
output(2, 128) <= input(46);
output(2, 129) <= input(44);
output(2, 130) <= input(1);
output(2, 131) <= input(2);
output(2, 132) <= input(3);
output(2, 133) <= input(4);
output(2, 134) <= input(5);
output(2, 135) <= input(6);
output(2, 136) <= input(7);
output(2, 137) <= input(8);
output(2, 138) <= input(9);
output(2, 139) <= input(10);
output(2, 140) <= input(11);
output(2, 141) <= input(12);
output(2, 142) <= input(13);
output(2, 143) <= input(14);
output(2, 144) <= input(46);
output(2, 145) <= input(44);
output(2, 146) <= input(1);
output(2, 147) <= input(2);
output(2, 148) <= input(3);
output(2, 149) <= input(4);
output(2, 150) <= input(5);
output(2, 151) <= input(6);
output(2, 152) <= input(7);
output(2, 153) <= input(8);
output(2, 154) <= input(9);
output(2, 155) <= input(10);
output(2, 156) <= input(11);
output(2, 157) <= input(12);
output(2, 158) <= input(13);
output(2, 159) <= input(14);
output(2, 160) <= input(46);
output(2, 161) <= input(44);
output(2, 162) <= input(1);
output(2, 163) <= input(2);
output(2, 164) <= input(3);
output(2, 165) <= input(4);
output(2, 166) <= input(5);
output(2, 167) <= input(6);
output(2, 168) <= input(7);
output(2, 169) <= input(8);
output(2, 170) <= input(9);
output(2, 171) <= input(10);
output(2, 172) <= input(11);
output(2, 173) <= input(12);
output(2, 174) <= input(13);
output(2, 175) <= input(14);
output(2, 176) <= input(46);
output(2, 177) <= input(44);
output(2, 178) <= input(1);
output(2, 179) <= input(2);
output(2, 180) <= input(3);
output(2, 181) <= input(4);
output(2, 182) <= input(5);
output(2, 183) <= input(6);
output(2, 184) <= input(7);
output(2, 185) <= input(8);
output(2, 186) <= input(9);
output(2, 187) <= input(10);
output(2, 188) <= input(11);
output(2, 189) <= input(12);
output(2, 190) <= input(13);
output(2, 191) <= input(14);
output(2, 192) <= input(47);
output(2, 193) <= input(45);
output(2, 194) <= input(17);
output(2, 195) <= input(18);
output(2, 196) <= input(19);
output(2, 197) <= input(20);
output(2, 198) <= input(21);
output(2, 199) <= input(22);
output(2, 200) <= input(23);
output(2, 201) <= input(24);
output(2, 202) <= input(25);
output(2, 203) <= input(26);
output(2, 204) <= input(27);
output(2, 205) <= input(28);
output(2, 206) <= input(29);
output(2, 207) <= input(30);
output(2, 208) <= input(47);
output(2, 209) <= input(45);
output(2, 210) <= input(17);
output(2, 211) <= input(18);
output(2, 212) <= input(19);
output(2, 213) <= input(20);
output(2, 214) <= input(21);
output(2, 215) <= input(22);
output(2, 216) <= input(23);
output(2, 217) <= input(24);
output(2, 218) <= input(25);
output(2, 219) <= input(26);
output(2, 220) <= input(27);
output(2, 221) <= input(28);
output(2, 222) <= input(29);
output(2, 223) <= input(30);
output(2, 224) <= input(47);
output(2, 225) <= input(45);
output(2, 226) <= input(17);
output(2, 227) <= input(18);
output(2, 228) <= input(19);
output(2, 229) <= input(20);
output(2, 230) <= input(21);
output(2, 231) <= input(22);
output(2, 232) <= input(23);
output(2, 233) <= input(24);
output(2, 234) <= input(25);
output(2, 235) <= input(26);
output(2, 236) <= input(27);
output(2, 237) <= input(28);
output(2, 238) <= input(29);
output(2, 239) <= input(30);
output(2, 240) <= input(47);
output(2, 241) <= input(45);
output(2, 242) <= input(17);
output(2, 243) <= input(18);
output(2, 244) <= input(19);
output(2, 245) <= input(20);
output(2, 246) <= input(21);
output(2, 247) <= input(22);
output(2, 248) <= input(23);
output(2, 249) <= input(24);
output(2, 250) <= input(25);
output(2, 251) <= input(26);
output(2, 252) <= input(27);
output(2, 253) <= input(28);
output(2, 254) <= input(29);
output(2, 255) <= input(30);
when "1101" =>
output(0, 0) <= input(0);
output(0, 1) <= input(1);
output(0, 2) <= input(2);
output(0, 3) <= input(3);
output(0, 4) <= input(4);
output(0, 5) <= input(5);
output(0, 6) <= input(6);
output(0, 7) <= input(7);
output(0, 8) <= input(8);
output(0, 9) <= input(9);
output(0, 10) <= input(10);
output(0, 11) <= input(11);
output(0, 12) <= input(12);
output(0, 13) <= input(13);
output(0, 14) <= input(14);
output(0, 15) <= input(15);
output(0, 16) <= input(0);
output(0, 17) <= input(1);
output(0, 18) <= input(2);
output(0, 19) <= input(3);
output(0, 20) <= input(4);
output(0, 21) <= input(5);
output(0, 22) <= input(6);
output(0, 23) <= input(7);
output(0, 24) <= input(8);
output(0, 25) <= input(9);
output(0, 26) <= input(10);
output(0, 27) <= input(11);
output(0, 28) <= input(12);
output(0, 29) <= input(13);
output(0, 30) <= input(14);
output(0, 31) <= input(15);
output(0, 32) <= input(0);
output(0, 33) <= input(1);
output(0, 34) <= input(2);
output(0, 35) <= input(3);
output(0, 36) <= input(4);
output(0, 37) <= input(5);
output(0, 38) <= input(6);
output(0, 39) <= input(7);
output(0, 40) <= input(8);
output(0, 41) <= input(9);
output(0, 42) <= input(10);
output(0, 43) <= input(11);
output(0, 44) <= input(12);
output(0, 45) <= input(13);
output(0, 46) <= input(14);
output(0, 47) <= input(15);
output(0, 48) <= input(0);
output(0, 49) <= input(1);
output(0, 50) <= input(2);
output(0, 51) <= input(3);
output(0, 52) <= input(4);
output(0, 53) <= input(5);
output(0, 54) <= input(6);
output(0, 55) <= input(7);
output(0, 56) <= input(8);
output(0, 57) <= input(9);
output(0, 58) <= input(10);
output(0, 59) <= input(11);
output(0, 60) <= input(12);
output(0, 61) <= input(13);
output(0, 62) <= input(14);
output(0, 63) <= input(15);
output(0, 64) <= input(0);
output(0, 65) <= input(1);
output(0, 66) <= input(2);
output(0, 67) <= input(3);
output(0, 68) <= input(4);
output(0, 69) <= input(5);
output(0, 70) <= input(6);
output(0, 71) <= input(7);
output(0, 72) <= input(8);
output(0, 73) <= input(9);
output(0, 74) <= input(10);
output(0, 75) <= input(11);
output(0, 76) <= input(12);
output(0, 77) <= input(13);
output(0, 78) <= input(14);
output(0, 79) <= input(15);
output(0, 80) <= input(16);
output(0, 81) <= input(17);
output(0, 82) <= input(18);
output(0, 83) <= input(19);
output(0, 84) <= input(20);
output(0, 85) <= input(21);
output(0, 86) <= input(22);
output(0, 87) <= input(23);
output(0, 88) <= input(24);
output(0, 89) <= input(25);
output(0, 90) <= input(26);
output(0, 91) <= input(27);
output(0, 92) <= input(28);
output(0, 93) <= input(29);
output(0, 94) <= input(30);
output(0, 95) <= input(31);
output(0, 96) <= input(16);
output(0, 97) <= input(17);
output(0, 98) <= input(18);
output(0, 99) <= input(19);
output(0, 100) <= input(20);
output(0, 101) <= input(21);
output(0, 102) <= input(22);
output(0, 103) <= input(23);
output(0, 104) <= input(24);
output(0, 105) <= input(25);
output(0, 106) <= input(26);
output(0, 107) <= input(27);
output(0, 108) <= input(28);
output(0, 109) <= input(29);
output(0, 110) <= input(30);
output(0, 111) <= input(31);
output(0, 112) <= input(16);
output(0, 113) <= input(17);
output(0, 114) <= input(18);
output(0, 115) <= input(19);
output(0, 116) <= input(20);
output(0, 117) <= input(21);
output(0, 118) <= input(22);
output(0, 119) <= input(23);
output(0, 120) <= input(24);
output(0, 121) <= input(25);
output(0, 122) <= input(26);
output(0, 123) <= input(27);
output(0, 124) <= input(28);
output(0, 125) <= input(29);
output(0, 126) <= input(30);
output(0, 127) <= input(31);
output(0, 128) <= input(16);
output(0, 129) <= input(17);
output(0, 130) <= input(18);
output(0, 131) <= input(19);
output(0, 132) <= input(20);
output(0, 133) <= input(21);
output(0, 134) <= input(22);
output(0, 135) <= input(23);
output(0, 136) <= input(24);
output(0, 137) <= input(25);
output(0, 138) <= input(26);
output(0, 139) <= input(27);
output(0, 140) <= input(28);
output(0, 141) <= input(29);
output(0, 142) <= input(30);
output(0, 143) <= input(31);
output(0, 144) <= input(16);
output(0, 145) <= input(17);
output(0, 146) <= input(18);
output(0, 147) <= input(19);
output(0, 148) <= input(20);
output(0, 149) <= input(21);
output(0, 150) <= input(22);
output(0, 151) <= input(23);
output(0, 152) <= input(24);
output(0, 153) <= input(25);
output(0, 154) <= input(26);
output(0, 155) <= input(27);
output(0, 156) <= input(28);
output(0, 157) <= input(29);
output(0, 158) <= input(30);
output(0, 159) <= input(31);
output(0, 160) <= input(32);
output(0, 161) <= input(0);
output(0, 162) <= input(1);
output(0, 163) <= input(2);
output(0, 164) <= input(3);
output(0, 165) <= input(4);
output(0, 166) <= input(5);
output(0, 167) <= input(6);
output(0, 168) <= input(7);
output(0, 169) <= input(8);
output(0, 170) <= input(9);
output(0, 171) <= input(10);
output(0, 172) <= input(11);
output(0, 173) <= input(12);
output(0, 174) <= input(13);
output(0, 175) <= input(14);
output(0, 176) <= input(32);
output(0, 177) <= input(0);
output(0, 178) <= input(1);
output(0, 179) <= input(2);
output(0, 180) <= input(3);
output(0, 181) <= input(4);
output(0, 182) <= input(5);
output(0, 183) <= input(6);
output(0, 184) <= input(7);
output(0, 185) <= input(8);
output(0, 186) <= input(9);
output(0, 187) <= input(10);
output(0, 188) <= input(11);
output(0, 189) <= input(12);
output(0, 190) <= input(13);
output(0, 191) <= input(14);
output(0, 192) <= input(32);
output(0, 193) <= input(0);
output(0, 194) <= input(1);
output(0, 195) <= input(2);
output(0, 196) <= input(3);
output(0, 197) <= input(4);
output(0, 198) <= input(5);
output(0, 199) <= input(6);
output(0, 200) <= input(7);
output(0, 201) <= input(8);
output(0, 202) <= input(9);
output(0, 203) <= input(10);
output(0, 204) <= input(11);
output(0, 205) <= input(12);
output(0, 206) <= input(13);
output(0, 207) <= input(14);
output(0, 208) <= input(32);
output(0, 209) <= input(0);
output(0, 210) <= input(1);
output(0, 211) <= input(2);
output(0, 212) <= input(3);
output(0, 213) <= input(4);
output(0, 214) <= input(5);
output(0, 215) <= input(6);
output(0, 216) <= input(7);
output(0, 217) <= input(8);
output(0, 218) <= input(9);
output(0, 219) <= input(10);
output(0, 220) <= input(11);
output(0, 221) <= input(12);
output(0, 222) <= input(13);
output(0, 223) <= input(14);
output(0, 224) <= input(32);
output(0, 225) <= input(0);
output(0, 226) <= input(1);
output(0, 227) <= input(2);
output(0, 228) <= input(3);
output(0, 229) <= input(4);
output(0, 230) <= input(5);
output(0, 231) <= input(6);
output(0, 232) <= input(7);
output(0, 233) <= input(8);
output(0, 234) <= input(9);
output(0, 235) <= input(10);
output(0, 236) <= input(11);
output(0, 237) <= input(12);
output(0, 238) <= input(13);
output(0, 239) <= input(14);
output(0, 240) <= input(32);
output(0, 241) <= input(0);
output(0, 242) <= input(1);
output(0, 243) <= input(2);
output(0, 244) <= input(3);
output(0, 245) <= input(4);
output(0, 246) <= input(5);
output(0, 247) <= input(6);
output(0, 248) <= input(7);
output(0, 249) <= input(8);
output(0, 250) <= input(9);
output(0, 251) <= input(10);
output(0, 252) <= input(11);
output(0, 253) <= input(12);
output(0, 254) <= input(13);
output(0, 255) <= input(14);
output(1, 0) <= input(33);
output(1, 1) <= input(1);
output(1, 2) <= input(2);
output(1, 3) <= input(3);
output(1, 4) <= input(4);
output(1, 5) <= input(5);
output(1, 6) <= input(6);
output(1, 7) <= input(7);
output(1, 8) <= input(8);
output(1, 9) <= input(9);
output(1, 10) <= input(10);
output(1, 11) <= input(11);
output(1, 12) <= input(12);
output(1, 13) <= input(13);
output(1, 14) <= input(14);
output(1, 15) <= input(15);
output(1, 16) <= input(33);
output(1, 17) <= input(1);
output(1, 18) <= input(2);
output(1, 19) <= input(3);
output(1, 20) <= input(4);
output(1, 21) <= input(5);
output(1, 22) <= input(6);
output(1, 23) <= input(7);
output(1, 24) <= input(8);
output(1, 25) <= input(9);
output(1, 26) <= input(10);
output(1, 27) <= input(11);
output(1, 28) <= input(12);
output(1, 29) <= input(13);
output(1, 30) <= input(14);
output(1, 31) <= input(15);
output(1, 32) <= input(33);
output(1, 33) <= input(1);
output(1, 34) <= input(2);
output(1, 35) <= input(3);
output(1, 36) <= input(4);
output(1, 37) <= input(5);
output(1, 38) <= input(6);
output(1, 39) <= input(7);
output(1, 40) <= input(8);
output(1, 41) <= input(9);
output(1, 42) <= input(10);
output(1, 43) <= input(11);
output(1, 44) <= input(12);
output(1, 45) <= input(13);
output(1, 46) <= input(14);
output(1, 47) <= input(15);
output(1, 48) <= input(33);
output(1, 49) <= input(1);
output(1, 50) <= input(2);
output(1, 51) <= input(3);
output(1, 52) <= input(4);
output(1, 53) <= input(5);
output(1, 54) <= input(6);
output(1, 55) <= input(7);
output(1, 56) <= input(8);
output(1, 57) <= input(9);
output(1, 58) <= input(10);
output(1, 59) <= input(11);
output(1, 60) <= input(12);
output(1, 61) <= input(13);
output(1, 62) <= input(14);
output(1, 63) <= input(15);
output(1, 64) <= input(33);
output(1, 65) <= input(1);
output(1, 66) <= input(2);
output(1, 67) <= input(3);
output(1, 68) <= input(4);
output(1, 69) <= input(5);
output(1, 70) <= input(6);
output(1, 71) <= input(7);
output(1, 72) <= input(8);
output(1, 73) <= input(9);
output(1, 74) <= input(10);
output(1, 75) <= input(11);
output(1, 76) <= input(12);
output(1, 77) <= input(13);
output(1, 78) <= input(14);
output(1, 79) <= input(15);
output(1, 80) <= input(33);
output(1, 81) <= input(1);
output(1, 82) <= input(2);
output(1, 83) <= input(3);
output(1, 84) <= input(4);
output(1, 85) <= input(5);
output(1, 86) <= input(6);
output(1, 87) <= input(7);
output(1, 88) <= input(8);
output(1, 89) <= input(9);
output(1, 90) <= input(10);
output(1, 91) <= input(11);
output(1, 92) <= input(12);
output(1, 93) <= input(13);
output(1, 94) <= input(14);
output(1, 95) <= input(15);
output(1, 96) <= input(33);
output(1, 97) <= input(1);
output(1, 98) <= input(2);
output(1, 99) <= input(3);
output(1, 100) <= input(4);
output(1, 101) <= input(5);
output(1, 102) <= input(6);
output(1, 103) <= input(7);
output(1, 104) <= input(8);
output(1, 105) <= input(9);
output(1, 106) <= input(10);
output(1, 107) <= input(11);
output(1, 108) <= input(12);
output(1, 109) <= input(13);
output(1, 110) <= input(14);
output(1, 111) <= input(15);
output(1, 112) <= input(33);
output(1, 113) <= input(1);
output(1, 114) <= input(2);
output(1, 115) <= input(3);
output(1, 116) <= input(4);
output(1, 117) <= input(5);
output(1, 118) <= input(6);
output(1, 119) <= input(7);
output(1, 120) <= input(8);
output(1, 121) <= input(9);
output(1, 122) <= input(10);
output(1, 123) <= input(11);
output(1, 124) <= input(12);
output(1, 125) <= input(13);
output(1, 126) <= input(14);
output(1, 127) <= input(15);
output(1, 128) <= input(34);
output(1, 129) <= input(17);
output(1, 130) <= input(18);
output(1, 131) <= input(19);
output(1, 132) <= input(20);
output(1, 133) <= input(21);
output(1, 134) <= input(22);
output(1, 135) <= input(23);
output(1, 136) <= input(24);
output(1, 137) <= input(25);
output(1, 138) <= input(26);
output(1, 139) <= input(27);
output(1, 140) <= input(28);
output(1, 141) <= input(29);
output(1, 142) <= input(30);
output(1, 143) <= input(31);
output(1, 144) <= input(34);
output(1, 145) <= input(17);
output(1, 146) <= input(18);
output(1, 147) <= input(19);
output(1, 148) <= input(20);
output(1, 149) <= input(21);
output(1, 150) <= input(22);
output(1, 151) <= input(23);
output(1, 152) <= input(24);
output(1, 153) <= input(25);
output(1, 154) <= input(26);
output(1, 155) <= input(27);
output(1, 156) <= input(28);
output(1, 157) <= input(29);
output(1, 158) <= input(30);
output(1, 159) <= input(31);
output(1, 160) <= input(34);
output(1, 161) <= input(17);
output(1, 162) <= input(18);
output(1, 163) <= input(19);
output(1, 164) <= input(20);
output(1, 165) <= input(21);
output(1, 166) <= input(22);
output(1, 167) <= input(23);
output(1, 168) <= input(24);
output(1, 169) <= input(25);
output(1, 170) <= input(26);
output(1, 171) <= input(27);
output(1, 172) <= input(28);
output(1, 173) <= input(29);
output(1, 174) <= input(30);
output(1, 175) <= input(31);
output(1, 176) <= input(34);
output(1, 177) <= input(17);
output(1, 178) <= input(18);
output(1, 179) <= input(19);
output(1, 180) <= input(20);
output(1, 181) <= input(21);
output(1, 182) <= input(22);
output(1, 183) <= input(23);
output(1, 184) <= input(24);
output(1, 185) <= input(25);
output(1, 186) <= input(26);
output(1, 187) <= input(27);
output(1, 188) <= input(28);
output(1, 189) <= input(29);
output(1, 190) <= input(30);
output(1, 191) <= input(31);
output(1, 192) <= input(34);
output(1, 193) <= input(17);
output(1, 194) <= input(18);
output(1, 195) <= input(19);
output(1, 196) <= input(20);
output(1, 197) <= input(21);
output(1, 198) <= input(22);
output(1, 199) <= input(23);
output(1, 200) <= input(24);
output(1, 201) <= input(25);
output(1, 202) <= input(26);
output(1, 203) <= input(27);
output(1, 204) <= input(28);
output(1, 205) <= input(29);
output(1, 206) <= input(30);
output(1, 207) <= input(31);
output(1, 208) <= input(34);
output(1, 209) <= input(17);
output(1, 210) <= input(18);
output(1, 211) <= input(19);
output(1, 212) <= input(20);
output(1, 213) <= input(21);
output(1, 214) <= input(22);
output(1, 215) <= input(23);
output(1, 216) <= input(24);
output(1, 217) <= input(25);
output(1, 218) <= input(26);
output(1, 219) <= input(27);
output(1, 220) <= input(28);
output(1, 221) <= input(29);
output(1, 222) <= input(30);
output(1, 223) <= input(31);
output(1, 224) <= input(34);
output(1, 225) <= input(17);
output(1, 226) <= input(18);
output(1, 227) <= input(19);
output(1, 228) <= input(20);
output(1, 229) <= input(21);
output(1, 230) <= input(22);
output(1, 231) <= input(23);
output(1, 232) <= input(24);
output(1, 233) <= input(25);
output(1, 234) <= input(26);
output(1, 235) <= input(27);
output(1, 236) <= input(28);
output(1, 237) <= input(29);
output(1, 238) <= input(30);
output(1, 239) <= input(31);
output(1, 240) <= input(34);
output(1, 241) <= input(17);
output(1, 242) <= input(18);
output(1, 243) <= input(19);
output(1, 244) <= input(20);
output(1, 245) <= input(21);
output(1, 246) <= input(22);
output(1, 247) <= input(23);
output(1, 248) <= input(24);
output(1, 249) <= input(25);
output(1, 250) <= input(26);
output(1, 251) <= input(27);
output(1, 252) <= input(28);
output(1, 253) <= input(29);
output(1, 254) <= input(30);
output(1, 255) <= input(31);
output(2, 0) <= input(35);
output(2, 1) <= input(1);
output(2, 2) <= input(2);
output(2, 3) <= input(3);
output(2, 4) <= input(4);
output(2, 5) <= input(5);
output(2, 6) <= input(6);
output(2, 7) <= input(7);
output(2, 8) <= input(8);
output(2, 9) <= input(9);
output(2, 10) <= input(10);
output(2, 11) <= input(11);
output(2, 12) <= input(12);
output(2, 13) <= input(13);
output(2, 14) <= input(14);
output(2, 15) <= input(15);
output(2, 16) <= input(35);
output(2, 17) <= input(1);
output(2, 18) <= input(2);
output(2, 19) <= input(3);
output(2, 20) <= input(4);
output(2, 21) <= input(5);
output(2, 22) <= input(6);
output(2, 23) <= input(7);
output(2, 24) <= input(8);
output(2, 25) <= input(9);
output(2, 26) <= input(10);
output(2, 27) <= input(11);
output(2, 28) <= input(12);
output(2, 29) <= input(13);
output(2, 30) <= input(14);
output(2, 31) <= input(15);
output(2, 32) <= input(35);
output(2, 33) <= input(1);
output(2, 34) <= input(2);
output(2, 35) <= input(3);
output(2, 36) <= input(4);
output(2, 37) <= input(5);
output(2, 38) <= input(6);
output(2, 39) <= input(7);
output(2, 40) <= input(8);
output(2, 41) <= input(9);
output(2, 42) <= input(10);
output(2, 43) <= input(11);
output(2, 44) <= input(12);
output(2, 45) <= input(13);
output(2, 46) <= input(14);
output(2, 47) <= input(15);
output(2, 48) <= input(35);
output(2, 49) <= input(1);
output(2, 50) <= input(2);
output(2, 51) <= input(3);
output(2, 52) <= input(4);
output(2, 53) <= input(5);
output(2, 54) <= input(6);
output(2, 55) <= input(7);
output(2, 56) <= input(8);
output(2, 57) <= input(9);
output(2, 58) <= input(10);
output(2, 59) <= input(11);
output(2, 60) <= input(12);
output(2, 61) <= input(13);
output(2, 62) <= input(14);
output(2, 63) <= input(15);
output(2, 64) <= input(35);
output(2, 65) <= input(1);
output(2, 66) <= input(2);
output(2, 67) <= input(3);
output(2, 68) <= input(4);
output(2, 69) <= input(5);
output(2, 70) <= input(6);
output(2, 71) <= input(7);
output(2, 72) <= input(8);
output(2, 73) <= input(9);
output(2, 74) <= input(10);
output(2, 75) <= input(11);
output(2, 76) <= input(12);
output(2, 77) <= input(13);
output(2, 78) <= input(14);
output(2, 79) <= input(15);
output(2, 80) <= input(35);
output(2, 81) <= input(1);
output(2, 82) <= input(2);
output(2, 83) <= input(3);
output(2, 84) <= input(4);
output(2, 85) <= input(5);
output(2, 86) <= input(6);
output(2, 87) <= input(7);
output(2, 88) <= input(8);
output(2, 89) <= input(9);
output(2, 90) <= input(10);
output(2, 91) <= input(11);
output(2, 92) <= input(12);
output(2, 93) <= input(13);
output(2, 94) <= input(14);
output(2, 95) <= input(15);
output(2, 96) <= input(35);
output(2, 97) <= input(1);
output(2, 98) <= input(2);
output(2, 99) <= input(3);
output(2, 100) <= input(4);
output(2, 101) <= input(5);
output(2, 102) <= input(6);
output(2, 103) <= input(7);
output(2, 104) <= input(8);
output(2, 105) <= input(9);
output(2, 106) <= input(10);
output(2, 107) <= input(11);
output(2, 108) <= input(12);
output(2, 109) <= input(13);
output(2, 110) <= input(14);
output(2, 111) <= input(15);
output(2, 112) <= input(35);
output(2, 113) <= input(1);
output(2, 114) <= input(2);
output(2, 115) <= input(3);
output(2, 116) <= input(4);
output(2, 117) <= input(5);
output(2, 118) <= input(6);
output(2, 119) <= input(7);
output(2, 120) <= input(8);
output(2, 121) <= input(9);
output(2, 122) <= input(10);
output(2, 123) <= input(11);
output(2, 124) <= input(12);
output(2, 125) <= input(13);
output(2, 126) <= input(14);
output(2, 127) <= input(15);
output(2, 128) <= input(35);
output(2, 129) <= input(1);
output(2, 130) <= input(2);
output(2, 131) <= input(3);
output(2, 132) <= input(4);
output(2, 133) <= input(5);
output(2, 134) <= input(6);
output(2, 135) <= input(7);
output(2, 136) <= input(8);
output(2, 137) <= input(9);
output(2, 138) <= input(10);
output(2, 139) <= input(11);
output(2, 140) <= input(12);
output(2, 141) <= input(13);
output(2, 142) <= input(14);
output(2, 143) <= input(15);
output(2, 144) <= input(35);
output(2, 145) <= input(1);
output(2, 146) <= input(2);
output(2, 147) <= input(3);
output(2, 148) <= input(4);
output(2, 149) <= input(5);
output(2, 150) <= input(6);
output(2, 151) <= input(7);
output(2, 152) <= input(8);
output(2, 153) <= input(9);
output(2, 154) <= input(10);
output(2, 155) <= input(11);
output(2, 156) <= input(12);
output(2, 157) <= input(13);
output(2, 158) <= input(14);
output(2, 159) <= input(15);
output(2, 160) <= input(35);
output(2, 161) <= input(1);
output(2, 162) <= input(2);
output(2, 163) <= input(3);
output(2, 164) <= input(4);
output(2, 165) <= input(5);
output(2, 166) <= input(6);
output(2, 167) <= input(7);
output(2, 168) <= input(8);
output(2, 169) <= input(9);
output(2, 170) <= input(10);
output(2, 171) <= input(11);
output(2, 172) <= input(12);
output(2, 173) <= input(13);
output(2, 174) <= input(14);
output(2, 175) <= input(15);
output(2, 176) <= input(35);
output(2, 177) <= input(1);
output(2, 178) <= input(2);
output(2, 179) <= input(3);
output(2, 180) <= input(4);
output(2, 181) <= input(5);
output(2, 182) <= input(6);
output(2, 183) <= input(7);
output(2, 184) <= input(8);
output(2, 185) <= input(9);
output(2, 186) <= input(10);
output(2, 187) <= input(11);
output(2, 188) <= input(12);
output(2, 189) <= input(13);
output(2, 190) <= input(14);
output(2, 191) <= input(15);
output(2, 192) <= input(35);
output(2, 193) <= input(1);
output(2, 194) <= input(2);
output(2, 195) <= input(3);
output(2, 196) <= input(4);
output(2, 197) <= input(5);
output(2, 198) <= input(6);
output(2, 199) <= input(7);
output(2, 200) <= input(8);
output(2, 201) <= input(9);
output(2, 202) <= input(10);
output(2, 203) <= input(11);
output(2, 204) <= input(12);
output(2, 205) <= input(13);
output(2, 206) <= input(14);
output(2, 207) <= input(15);
output(2, 208) <= input(35);
output(2, 209) <= input(1);
output(2, 210) <= input(2);
output(2, 211) <= input(3);
output(2, 212) <= input(4);
output(2, 213) <= input(5);
output(2, 214) <= input(6);
output(2, 215) <= input(7);
output(2, 216) <= input(8);
output(2, 217) <= input(9);
output(2, 218) <= input(10);
output(2, 219) <= input(11);
output(2, 220) <= input(12);
output(2, 221) <= input(13);
output(2, 222) <= input(14);
output(2, 223) <= input(15);
output(2, 224) <= input(35);
output(2, 225) <= input(1);
output(2, 226) <= input(2);
output(2, 227) <= input(3);
output(2, 228) <= input(4);
output(2, 229) <= input(5);
output(2, 230) <= input(6);
output(2, 231) <= input(7);
output(2, 232) <= input(8);
output(2, 233) <= input(9);
output(2, 234) <= input(10);
output(2, 235) <= input(11);
output(2, 236) <= input(12);
output(2, 237) <= input(13);
output(2, 238) <= input(14);
output(2, 239) <= input(15);
output(2, 240) <= input(35);
output(2, 241) <= input(1);
output(2, 242) <= input(2);
output(2, 243) <= input(3);
output(2, 244) <= input(4);
output(2, 245) <= input(5);
output(2, 246) <= input(6);
output(2, 247) <= input(7);
output(2, 248) <= input(8);
output(2, 249) <= input(9);
output(2, 250) <= input(10);
output(2, 251) <= input(11);
output(2, 252) <= input(12);
output(2, 253) <= input(13);
output(2, 254) <= input(14);
output(2, 255) <= input(15);
output(3, 0) <= input(17);
output(3, 1) <= input(18);
output(3, 2) <= input(19);
output(3, 3) <= input(20);
output(3, 4) <= input(21);
output(3, 5) <= input(22);
output(3, 6) <= input(23);
output(3, 7) <= input(24);
output(3, 8) <= input(25);
output(3, 9) <= input(26);
output(3, 10) <= input(27);
output(3, 11) <= input(28);
output(3, 12) <= input(29);
output(3, 13) <= input(30);
output(3, 14) <= input(31);
output(3, 15) <= input(36);
output(3, 16) <= input(17);
output(3, 17) <= input(18);
output(3, 18) <= input(19);
output(3, 19) <= input(20);
output(3, 20) <= input(21);
output(3, 21) <= input(22);
output(3, 22) <= input(23);
output(3, 23) <= input(24);
output(3, 24) <= input(25);
output(3, 25) <= input(26);
output(3, 26) <= input(27);
output(3, 27) <= input(28);
output(3, 28) <= input(29);
output(3, 29) <= input(30);
output(3, 30) <= input(31);
output(3, 31) <= input(36);
output(3, 32) <= input(17);
output(3, 33) <= input(18);
output(3, 34) <= input(19);
output(3, 35) <= input(20);
output(3, 36) <= input(21);
output(3, 37) <= input(22);
output(3, 38) <= input(23);
output(3, 39) <= input(24);
output(3, 40) <= input(25);
output(3, 41) <= input(26);
output(3, 42) <= input(27);
output(3, 43) <= input(28);
output(3, 44) <= input(29);
output(3, 45) <= input(30);
output(3, 46) <= input(31);
output(3, 47) <= input(36);
output(3, 48) <= input(17);
output(3, 49) <= input(18);
output(3, 50) <= input(19);
output(3, 51) <= input(20);
output(3, 52) <= input(21);
output(3, 53) <= input(22);
output(3, 54) <= input(23);
output(3, 55) <= input(24);
output(3, 56) <= input(25);
output(3, 57) <= input(26);
output(3, 58) <= input(27);
output(3, 59) <= input(28);
output(3, 60) <= input(29);
output(3, 61) <= input(30);
output(3, 62) <= input(31);
output(3, 63) <= input(36);
output(3, 64) <= input(17);
output(3, 65) <= input(18);
output(3, 66) <= input(19);
output(3, 67) <= input(20);
output(3, 68) <= input(21);
output(3, 69) <= input(22);
output(3, 70) <= input(23);
output(3, 71) <= input(24);
output(3, 72) <= input(25);
output(3, 73) <= input(26);
output(3, 74) <= input(27);
output(3, 75) <= input(28);
output(3, 76) <= input(29);
output(3, 77) <= input(30);
output(3, 78) <= input(31);
output(3, 79) <= input(36);
output(3, 80) <= input(17);
output(3, 81) <= input(18);
output(3, 82) <= input(19);
output(3, 83) <= input(20);
output(3, 84) <= input(21);
output(3, 85) <= input(22);
output(3, 86) <= input(23);
output(3, 87) <= input(24);
output(3, 88) <= input(25);
output(3, 89) <= input(26);
output(3, 90) <= input(27);
output(3, 91) <= input(28);
output(3, 92) <= input(29);
output(3, 93) <= input(30);
output(3, 94) <= input(31);
output(3, 95) <= input(36);
output(3, 96) <= input(17);
output(3, 97) <= input(18);
output(3, 98) <= input(19);
output(3, 99) <= input(20);
output(3, 100) <= input(21);
output(3, 101) <= input(22);
output(3, 102) <= input(23);
output(3, 103) <= input(24);
output(3, 104) <= input(25);
output(3, 105) <= input(26);
output(3, 106) <= input(27);
output(3, 107) <= input(28);
output(3, 108) <= input(29);
output(3, 109) <= input(30);
output(3, 110) <= input(31);
output(3, 111) <= input(36);
output(3, 112) <= input(17);
output(3, 113) <= input(18);
output(3, 114) <= input(19);
output(3, 115) <= input(20);
output(3, 116) <= input(21);
output(3, 117) <= input(22);
output(3, 118) <= input(23);
output(3, 119) <= input(24);
output(3, 120) <= input(25);
output(3, 121) <= input(26);
output(3, 122) <= input(27);
output(3, 123) <= input(28);
output(3, 124) <= input(29);
output(3, 125) <= input(30);
output(3, 126) <= input(31);
output(3, 127) <= input(36);
output(3, 128) <= input(17);
output(3, 129) <= input(18);
output(3, 130) <= input(19);
output(3, 131) <= input(20);
output(3, 132) <= input(21);
output(3, 133) <= input(22);
output(3, 134) <= input(23);
output(3, 135) <= input(24);
output(3, 136) <= input(25);
output(3, 137) <= input(26);
output(3, 138) <= input(27);
output(3, 139) <= input(28);
output(3, 140) <= input(29);
output(3, 141) <= input(30);
output(3, 142) <= input(31);
output(3, 143) <= input(36);
output(3, 144) <= input(17);
output(3, 145) <= input(18);
output(3, 146) <= input(19);
output(3, 147) <= input(20);
output(3, 148) <= input(21);
output(3, 149) <= input(22);
output(3, 150) <= input(23);
output(3, 151) <= input(24);
output(3, 152) <= input(25);
output(3, 153) <= input(26);
output(3, 154) <= input(27);
output(3, 155) <= input(28);
output(3, 156) <= input(29);
output(3, 157) <= input(30);
output(3, 158) <= input(31);
output(3, 159) <= input(36);
output(3, 160) <= input(17);
output(3, 161) <= input(18);
output(3, 162) <= input(19);
output(3, 163) <= input(20);
output(3, 164) <= input(21);
output(3, 165) <= input(22);
output(3, 166) <= input(23);
output(3, 167) <= input(24);
output(3, 168) <= input(25);
output(3, 169) <= input(26);
output(3, 170) <= input(27);
output(3, 171) <= input(28);
output(3, 172) <= input(29);
output(3, 173) <= input(30);
output(3, 174) <= input(31);
output(3, 175) <= input(36);
output(3, 176) <= input(17);
output(3, 177) <= input(18);
output(3, 178) <= input(19);
output(3, 179) <= input(20);
output(3, 180) <= input(21);
output(3, 181) <= input(22);
output(3, 182) <= input(23);
output(3, 183) <= input(24);
output(3, 184) <= input(25);
output(3, 185) <= input(26);
output(3, 186) <= input(27);
output(3, 187) <= input(28);
output(3, 188) <= input(29);
output(3, 189) <= input(30);
output(3, 190) <= input(31);
output(3, 191) <= input(36);
output(3, 192) <= input(17);
output(3, 193) <= input(18);
output(3, 194) <= input(19);
output(3, 195) <= input(20);
output(3, 196) <= input(21);
output(3, 197) <= input(22);
output(3, 198) <= input(23);
output(3, 199) <= input(24);
output(3, 200) <= input(25);
output(3, 201) <= input(26);
output(3, 202) <= input(27);
output(3, 203) <= input(28);
output(3, 204) <= input(29);
output(3, 205) <= input(30);
output(3, 206) <= input(31);
output(3, 207) <= input(36);
output(3, 208) <= input(17);
output(3, 209) <= input(18);
output(3, 210) <= input(19);
output(3, 211) <= input(20);
output(3, 212) <= input(21);
output(3, 213) <= input(22);
output(3, 214) <= input(23);
output(3, 215) <= input(24);
output(3, 216) <= input(25);
output(3, 217) <= input(26);
output(3, 218) <= input(27);
output(3, 219) <= input(28);
output(3, 220) <= input(29);
output(3, 221) <= input(30);
output(3, 222) <= input(31);
output(3, 223) <= input(36);
output(3, 224) <= input(17);
output(3, 225) <= input(18);
output(3, 226) <= input(19);
output(3, 227) <= input(20);
output(3, 228) <= input(21);
output(3, 229) <= input(22);
output(3, 230) <= input(23);
output(3, 231) <= input(24);
output(3, 232) <= input(25);
output(3, 233) <= input(26);
output(3, 234) <= input(27);
output(3, 235) <= input(28);
output(3, 236) <= input(29);
output(3, 237) <= input(30);
output(3, 238) <= input(31);
output(3, 239) <= input(36);
output(3, 240) <= input(17);
output(3, 241) <= input(18);
output(3, 242) <= input(19);
output(3, 243) <= input(20);
output(3, 244) <= input(21);
output(3, 245) <= input(22);
output(3, 246) <= input(23);
output(3, 247) <= input(24);
output(3, 248) <= input(25);
output(3, 249) <= input(26);
output(3, 250) <= input(27);
output(3, 251) <= input(28);
output(3, 252) <= input(29);
output(3, 253) <= input(30);
output(3, 254) <= input(31);
output(3, 255) <= input(36);
output(4, 0) <= input(17);
output(4, 1) <= input(18);
output(4, 2) <= input(19);
output(4, 3) <= input(20);
output(4, 4) <= input(21);
output(4, 5) <= input(22);
output(4, 6) <= input(23);
output(4, 7) <= input(24);
output(4, 8) <= input(25);
output(4, 9) <= input(26);
output(4, 10) <= input(27);
output(4, 11) <= input(28);
output(4, 12) <= input(29);
output(4, 13) <= input(30);
output(4, 14) <= input(31);
output(4, 15) <= input(36);
output(4, 16) <= input(17);
output(4, 17) <= input(18);
output(4, 18) <= input(19);
output(4, 19) <= input(20);
output(4, 20) <= input(21);
output(4, 21) <= input(22);
output(4, 22) <= input(23);
output(4, 23) <= input(24);
output(4, 24) <= input(25);
output(4, 25) <= input(26);
output(4, 26) <= input(27);
output(4, 27) <= input(28);
output(4, 28) <= input(29);
output(4, 29) <= input(30);
output(4, 30) <= input(31);
output(4, 31) <= input(36);
output(4, 32) <= input(17);
output(4, 33) <= input(18);
output(4, 34) <= input(19);
output(4, 35) <= input(20);
output(4, 36) <= input(21);
output(4, 37) <= input(22);
output(4, 38) <= input(23);
output(4, 39) <= input(24);
output(4, 40) <= input(25);
output(4, 41) <= input(26);
output(4, 42) <= input(27);
output(4, 43) <= input(28);
output(4, 44) <= input(29);
output(4, 45) <= input(30);
output(4, 46) <= input(31);
output(4, 47) <= input(36);
output(4, 48) <= input(17);
output(4, 49) <= input(18);
output(4, 50) <= input(19);
output(4, 51) <= input(20);
output(4, 52) <= input(21);
output(4, 53) <= input(22);
output(4, 54) <= input(23);
output(4, 55) <= input(24);
output(4, 56) <= input(25);
output(4, 57) <= input(26);
output(4, 58) <= input(27);
output(4, 59) <= input(28);
output(4, 60) <= input(29);
output(4, 61) <= input(30);
output(4, 62) <= input(31);
output(4, 63) <= input(36);
output(4, 64) <= input(17);
output(4, 65) <= input(18);
output(4, 66) <= input(19);
output(4, 67) <= input(20);
output(4, 68) <= input(21);
output(4, 69) <= input(22);
output(4, 70) <= input(23);
output(4, 71) <= input(24);
output(4, 72) <= input(25);
output(4, 73) <= input(26);
output(4, 74) <= input(27);
output(4, 75) <= input(28);
output(4, 76) <= input(29);
output(4, 77) <= input(30);
output(4, 78) <= input(31);
output(4, 79) <= input(36);
output(4, 80) <= input(17);
output(4, 81) <= input(18);
output(4, 82) <= input(19);
output(4, 83) <= input(20);
output(4, 84) <= input(21);
output(4, 85) <= input(22);
output(4, 86) <= input(23);
output(4, 87) <= input(24);
output(4, 88) <= input(25);
output(4, 89) <= input(26);
output(4, 90) <= input(27);
output(4, 91) <= input(28);
output(4, 92) <= input(29);
output(4, 93) <= input(30);
output(4, 94) <= input(31);
output(4, 95) <= input(36);
output(4, 96) <= input(17);
output(4, 97) <= input(18);
output(4, 98) <= input(19);
output(4, 99) <= input(20);
output(4, 100) <= input(21);
output(4, 101) <= input(22);
output(4, 102) <= input(23);
output(4, 103) <= input(24);
output(4, 104) <= input(25);
output(4, 105) <= input(26);
output(4, 106) <= input(27);
output(4, 107) <= input(28);
output(4, 108) <= input(29);
output(4, 109) <= input(30);
output(4, 110) <= input(31);
output(4, 111) <= input(36);
output(4, 112) <= input(17);
output(4, 113) <= input(18);
output(4, 114) <= input(19);
output(4, 115) <= input(20);
output(4, 116) <= input(21);
output(4, 117) <= input(22);
output(4, 118) <= input(23);
output(4, 119) <= input(24);
output(4, 120) <= input(25);
output(4, 121) <= input(26);
output(4, 122) <= input(27);
output(4, 123) <= input(28);
output(4, 124) <= input(29);
output(4, 125) <= input(30);
output(4, 126) <= input(31);
output(4, 127) <= input(36);
output(4, 128) <= input(17);
output(4, 129) <= input(18);
output(4, 130) <= input(19);
output(4, 131) <= input(20);
output(4, 132) <= input(21);
output(4, 133) <= input(22);
output(4, 134) <= input(23);
output(4, 135) <= input(24);
output(4, 136) <= input(25);
output(4, 137) <= input(26);
output(4, 138) <= input(27);
output(4, 139) <= input(28);
output(4, 140) <= input(29);
output(4, 141) <= input(30);
output(4, 142) <= input(31);
output(4, 143) <= input(36);
output(4, 144) <= input(17);
output(4, 145) <= input(18);
output(4, 146) <= input(19);
output(4, 147) <= input(20);
output(4, 148) <= input(21);
output(4, 149) <= input(22);
output(4, 150) <= input(23);
output(4, 151) <= input(24);
output(4, 152) <= input(25);
output(4, 153) <= input(26);
output(4, 154) <= input(27);
output(4, 155) <= input(28);
output(4, 156) <= input(29);
output(4, 157) <= input(30);
output(4, 158) <= input(31);
output(4, 159) <= input(36);
output(4, 160) <= input(17);
output(4, 161) <= input(18);
output(4, 162) <= input(19);
output(4, 163) <= input(20);
output(4, 164) <= input(21);
output(4, 165) <= input(22);
output(4, 166) <= input(23);
output(4, 167) <= input(24);
output(4, 168) <= input(25);
output(4, 169) <= input(26);
output(4, 170) <= input(27);
output(4, 171) <= input(28);
output(4, 172) <= input(29);
output(4, 173) <= input(30);
output(4, 174) <= input(31);
output(4, 175) <= input(36);
output(4, 176) <= input(17);
output(4, 177) <= input(18);
output(4, 178) <= input(19);
output(4, 179) <= input(20);
output(4, 180) <= input(21);
output(4, 181) <= input(22);
output(4, 182) <= input(23);
output(4, 183) <= input(24);
output(4, 184) <= input(25);
output(4, 185) <= input(26);
output(4, 186) <= input(27);
output(4, 187) <= input(28);
output(4, 188) <= input(29);
output(4, 189) <= input(30);
output(4, 190) <= input(31);
output(4, 191) <= input(36);
output(4, 192) <= input(17);
output(4, 193) <= input(18);
output(4, 194) <= input(19);
output(4, 195) <= input(20);
output(4, 196) <= input(21);
output(4, 197) <= input(22);
output(4, 198) <= input(23);
output(4, 199) <= input(24);
output(4, 200) <= input(25);
output(4, 201) <= input(26);
output(4, 202) <= input(27);
output(4, 203) <= input(28);
output(4, 204) <= input(29);
output(4, 205) <= input(30);
output(4, 206) <= input(31);
output(4, 207) <= input(36);
output(4, 208) <= input(17);
output(4, 209) <= input(18);
output(4, 210) <= input(19);
output(4, 211) <= input(20);
output(4, 212) <= input(21);
output(4, 213) <= input(22);
output(4, 214) <= input(23);
output(4, 215) <= input(24);
output(4, 216) <= input(25);
output(4, 217) <= input(26);
output(4, 218) <= input(27);
output(4, 219) <= input(28);
output(4, 220) <= input(29);
output(4, 221) <= input(30);
output(4, 222) <= input(31);
output(4, 223) <= input(36);
output(4, 224) <= input(17);
output(4, 225) <= input(18);
output(4, 226) <= input(19);
output(4, 227) <= input(20);
output(4, 228) <= input(21);
output(4, 229) <= input(22);
output(4, 230) <= input(23);
output(4, 231) <= input(24);
output(4, 232) <= input(25);
output(4, 233) <= input(26);
output(4, 234) <= input(27);
output(4, 235) <= input(28);
output(4, 236) <= input(29);
output(4, 237) <= input(30);
output(4, 238) <= input(31);
output(4, 239) <= input(36);
output(4, 240) <= input(1);
output(4, 241) <= input(2);
output(4, 242) <= input(3);
output(4, 243) <= input(4);
output(4, 244) <= input(5);
output(4, 245) <= input(6);
output(4, 246) <= input(7);
output(4, 247) <= input(8);
output(4, 248) <= input(9);
output(4, 249) <= input(10);
output(4, 250) <= input(11);
output(4, 251) <= input(12);
output(4, 252) <= input(13);
output(4, 253) <= input(14);
output(4, 254) <= input(15);
output(4, 255) <= input(37);
output(5, 0) <= input(17);
output(5, 1) <= input(18);
output(5, 2) <= input(19);
output(5, 3) <= input(20);
output(5, 4) <= input(21);
output(5, 5) <= input(22);
output(5, 6) <= input(23);
output(5, 7) <= input(24);
output(5, 8) <= input(25);
output(5, 9) <= input(26);
output(5, 10) <= input(27);
output(5, 11) <= input(28);
output(5, 12) <= input(29);
output(5, 13) <= input(30);
output(5, 14) <= input(31);
output(5, 15) <= input(36);
output(5, 16) <= input(17);
output(5, 17) <= input(18);
output(5, 18) <= input(19);
output(5, 19) <= input(20);
output(5, 20) <= input(21);
output(5, 21) <= input(22);
output(5, 22) <= input(23);
output(5, 23) <= input(24);
output(5, 24) <= input(25);
output(5, 25) <= input(26);
output(5, 26) <= input(27);
output(5, 27) <= input(28);
output(5, 28) <= input(29);
output(5, 29) <= input(30);
output(5, 30) <= input(31);
output(5, 31) <= input(36);
output(5, 32) <= input(17);
output(5, 33) <= input(18);
output(5, 34) <= input(19);
output(5, 35) <= input(20);
output(5, 36) <= input(21);
output(5, 37) <= input(22);
output(5, 38) <= input(23);
output(5, 39) <= input(24);
output(5, 40) <= input(25);
output(5, 41) <= input(26);
output(5, 42) <= input(27);
output(5, 43) <= input(28);
output(5, 44) <= input(29);
output(5, 45) <= input(30);
output(5, 46) <= input(31);
output(5, 47) <= input(36);
output(5, 48) <= input(17);
output(5, 49) <= input(18);
output(5, 50) <= input(19);
output(5, 51) <= input(20);
output(5, 52) <= input(21);
output(5, 53) <= input(22);
output(5, 54) <= input(23);
output(5, 55) <= input(24);
output(5, 56) <= input(25);
output(5, 57) <= input(26);
output(5, 58) <= input(27);
output(5, 59) <= input(28);
output(5, 60) <= input(29);
output(5, 61) <= input(30);
output(5, 62) <= input(31);
output(5, 63) <= input(36);
output(5, 64) <= input(17);
output(5, 65) <= input(18);
output(5, 66) <= input(19);
output(5, 67) <= input(20);
output(5, 68) <= input(21);
output(5, 69) <= input(22);
output(5, 70) <= input(23);
output(5, 71) <= input(24);
output(5, 72) <= input(25);
output(5, 73) <= input(26);
output(5, 74) <= input(27);
output(5, 75) <= input(28);
output(5, 76) <= input(29);
output(5, 77) <= input(30);
output(5, 78) <= input(31);
output(5, 79) <= input(36);
output(5, 80) <= input(17);
output(5, 81) <= input(18);
output(5, 82) <= input(19);
output(5, 83) <= input(20);
output(5, 84) <= input(21);
output(5, 85) <= input(22);
output(5, 86) <= input(23);
output(5, 87) <= input(24);
output(5, 88) <= input(25);
output(5, 89) <= input(26);
output(5, 90) <= input(27);
output(5, 91) <= input(28);
output(5, 92) <= input(29);
output(5, 93) <= input(30);
output(5, 94) <= input(31);
output(5, 95) <= input(36);
output(5, 96) <= input(17);
output(5, 97) <= input(18);
output(5, 98) <= input(19);
output(5, 99) <= input(20);
output(5, 100) <= input(21);
output(5, 101) <= input(22);
output(5, 102) <= input(23);
output(5, 103) <= input(24);
output(5, 104) <= input(25);
output(5, 105) <= input(26);
output(5, 106) <= input(27);
output(5, 107) <= input(28);
output(5, 108) <= input(29);
output(5, 109) <= input(30);
output(5, 110) <= input(31);
output(5, 111) <= input(36);
output(5, 112) <= input(1);
output(5, 113) <= input(2);
output(5, 114) <= input(3);
output(5, 115) <= input(4);
output(5, 116) <= input(5);
output(5, 117) <= input(6);
output(5, 118) <= input(7);
output(5, 119) <= input(8);
output(5, 120) <= input(9);
output(5, 121) <= input(10);
output(5, 122) <= input(11);
output(5, 123) <= input(12);
output(5, 124) <= input(13);
output(5, 125) <= input(14);
output(5, 126) <= input(15);
output(5, 127) <= input(37);
output(5, 128) <= input(1);
output(5, 129) <= input(2);
output(5, 130) <= input(3);
output(5, 131) <= input(4);
output(5, 132) <= input(5);
output(5, 133) <= input(6);
output(5, 134) <= input(7);
output(5, 135) <= input(8);
output(5, 136) <= input(9);
output(5, 137) <= input(10);
output(5, 138) <= input(11);
output(5, 139) <= input(12);
output(5, 140) <= input(13);
output(5, 141) <= input(14);
output(5, 142) <= input(15);
output(5, 143) <= input(37);
output(5, 144) <= input(1);
output(5, 145) <= input(2);
output(5, 146) <= input(3);
output(5, 147) <= input(4);
output(5, 148) <= input(5);
output(5, 149) <= input(6);
output(5, 150) <= input(7);
output(5, 151) <= input(8);
output(5, 152) <= input(9);
output(5, 153) <= input(10);
output(5, 154) <= input(11);
output(5, 155) <= input(12);
output(5, 156) <= input(13);
output(5, 157) <= input(14);
output(5, 158) <= input(15);
output(5, 159) <= input(37);
output(5, 160) <= input(1);
output(5, 161) <= input(2);
output(5, 162) <= input(3);
output(5, 163) <= input(4);
output(5, 164) <= input(5);
output(5, 165) <= input(6);
output(5, 166) <= input(7);
output(5, 167) <= input(8);
output(5, 168) <= input(9);
output(5, 169) <= input(10);
output(5, 170) <= input(11);
output(5, 171) <= input(12);
output(5, 172) <= input(13);
output(5, 173) <= input(14);
output(5, 174) <= input(15);
output(5, 175) <= input(37);
output(5, 176) <= input(1);
output(5, 177) <= input(2);
output(5, 178) <= input(3);
output(5, 179) <= input(4);
output(5, 180) <= input(5);
output(5, 181) <= input(6);
output(5, 182) <= input(7);
output(5, 183) <= input(8);
output(5, 184) <= input(9);
output(5, 185) <= input(10);
output(5, 186) <= input(11);
output(5, 187) <= input(12);
output(5, 188) <= input(13);
output(5, 189) <= input(14);
output(5, 190) <= input(15);
output(5, 191) <= input(37);
output(5, 192) <= input(1);
output(5, 193) <= input(2);
output(5, 194) <= input(3);
output(5, 195) <= input(4);
output(5, 196) <= input(5);
output(5, 197) <= input(6);
output(5, 198) <= input(7);
output(5, 199) <= input(8);
output(5, 200) <= input(9);
output(5, 201) <= input(10);
output(5, 202) <= input(11);
output(5, 203) <= input(12);
output(5, 204) <= input(13);
output(5, 205) <= input(14);
output(5, 206) <= input(15);
output(5, 207) <= input(37);
output(5, 208) <= input(1);
output(5, 209) <= input(2);
output(5, 210) <= input(3);
output(5, 211) <= input(4);
output(5, 212) <= input(5);
output(5, 213) <= input(6);
output(5, 214) <= input(7);
output(5, 215) <= input(8);
output(5, 216) <= input(9);
output(5, 217) <= input(10);
output(5, 218) <= input(11);
output(5, 219) <= input(12);
output(5, 220) <= input(13);
output(5, 221) <= input(14);
output(5, 222) <= input(15);
output(5, 223) <= input(37);
output(5, 224) <= input(1);
output(5, 225) <= input(2);
output(5, 226) <= input(3);
output(5, 227) <= input(4);
output(5, 228) <= input(5);
output(5, 229) <= input(6);
output(5, 230) <= input(7);
output(5, 231) <= input(8);
output(5, 232) <= input(9);
output(5, 233) <= input(10);
output(5, 234) <= input(11);
output(5, 235) <= input(12);
output(5, 236) <= input(13);
output(5, 237) <= input(14);
output(5, 238) <= input(15);
output(5, 239) <= input(37);
output(5, 240) <= input(18);
output(5, 241) <= input(19);
output(5, 242) <= input(20);
output(5, 243) <= input(21);
output(5, 244) <= input(22);
output(5, 245) <= input(23);
output(5, 246) <= input(24);
output(5, 247) <= input(25);
output(5, 248) <= input(26);
output(5, 249) <= input(27);
output(5, 250) <= input(28);
output(5, 251) <= input(29);
output(5, 252) <= input(30);
output(5, 253) <= input(31);
output(5, 254) <= input(36);
output(5, 255) <= input(38);
output(6, 0) <= input(17);
output(6, 1) <= input(18);
output(6, 2) <= input(19);
output(6, 3) <= input(20);
output(6, 4) <= input(21);
output(6, 5) <= input(22);
output(6, 6) <= input(23);
output(6, 7) <= input(24);
output(6, 8) <= input(25);
output(6, 9) <= input(26);
output(6, 10) <= input(27);
output(6, 11) <= input(28);
output(6, 12) <= input(29);
output(6, 13) <= input(30);
output(6, 14) <= input(31);
output(6, 15) <= input(36);
output(6, 16) <= input(17);
output(6, 17) <= input(18);
output(6, 18) <= input(19);
output(6, 19) <= input(20);
output(6, 20) <= input(21);
output(6, 21) <= input(22);
output(6, 22) <= input(23);
output(6, 23) <= input(24);
output(6, 24) <= input(25);
output(6, 25) <= input(26);
output(6, 26) <= input(27);
output(6, 27) <= input(28);
output(6, 28) <= input(29);
output(6, 29) <= input(30);
output(6, 30) <= input(31);
output(6, 31) <= input(36);
output(6, 32) <= input(17);
output(6, 33) <= input(18);
output(6, 34) <= input(19);
output(6, 35) <= input(20);
output(6, 36) <= input(21);
output(6, 37) <= input(22);
output(6, 38) <= input(23);
output(6, 39) <= input(24);
output(6, 40) <= input(25);
output(6, 41) <= input(26);
output(6, 42) <= input(27);
output(6, 43) <= input(28);
output(6, 44) <= input(29);
output(6, 45) <= input(30);
output(6, 46) <= input(31);
output(6, 47) <= input(36);
output(6, 48) <= input(17);
output(6, 49) <= input(18);
output(6, 50) <= input(19);
output(6, 51) <= input(20);
output(6, 52) <= input(21);
output(6, 53) <= input(22);
output(6, 54) <= input(23);
output(6, 55) <= input(24);
output(6, 56) <= input(25);
output(6, 57) <= input(26);
output(6, 58) <= input(27);
output(6, 59) <= input(28);
output(6, 60) <= input(29);
output(6, 61) <= input(30);
output(6, 62) <= input(31);
output(6, 63) <= input(36);
output(6, 64) <= input(17);
output(6, 65) <= input(18);
output(6, 66) <= input(19);
output(6, 67) <= input(20);
output(6, 68) <= input(21);
output(6, 69) <= input(22);
output(6, 70) <= input(23);
output(6, 71) <= input(24);
output(6, 72) <= input(25);
output(6, 73) <= input(26);
output(6, 74) <= input(27);
output(6, 75) <= input(28);
output(6, 76) <= input(29);
output(6, 77) <= input(30);
output(6, 78) <= input(31);
output(6, 79) <= input(36);
output(6, 80) <= input(1);
output(6, 81) <= input(2);
output(6, 82) <= input(3);
output(6, 83) <= input(4);
output(6, 84) <= input(5);
output(6, 85) <= input(6);
output(6, 86) <= input(7);
output(6, 87) <= input(8);
output(6, 88) <= input(9);
output(6, 89) <= input(10);
output(6, 90) <= input(11);
output(6, 91) <= input(12);
output(6, 92) <= input(13);
output(6, 93) <= input(14);
output(6, 94) <= input(15);
output(6, 95) <= input(37);
output(6, 96) <= input(1);
output(6, 97) <= input(2);
output(6, 98) <= input(3);
output(6, 99) <= input(4);
output(6, 100) <= input(5);
output(6, 101) <= input(6);
output(6, 102) <= input(7);
output(6, 103) <= input(8);
output(6, 104) <= input(9);
output(6, 105) <= input(10);
output(6, 106) <= input(11);
output(6, 107) <= input(12);
output(6, 108) <= input(13);
output(6, 109) <= input(14);
output(6, 110) <= input(15);
output(6, 111) <= input(37);
output(6, 112) <= input(1);
output(6, 113) <= input(2);
output(6, 114) <= input(3);
output(6, 115) <= input(4);
output(6, 116) <= input(5);
output(6, 117) <= input(6);
output(6, 118) <= input(7);
output(6, 119) <= input(8);
output(6, 120) <= input(9);
output(6, 121) <= input(10);
output(6, 122) <= input(11);
output(6, 123) <= input(12);
output(6, 124) <= input(13);
output(6, 125) <= input(14);
output(6, 126) <= input(15);
output(6, 127) <= input(37);
output(6, 128) <= input(1);
output(6, 129) <= input(2);
output(6, 130) <= input(3);
output(6, 131) <= input(4);
output(6, 132) <= input(5);
output(6, 133) <= input(6);
output(6, 134) <= input(7);
output(6, 135) <= input(8);
output(6, 136) <= input(9);
output(6, 137) <= input(10);
output(6, 138) <= input(11);
output(6, 139) <= input(12);
output(6, 140) <= input(13);
output(6, 141) <= input(14);
output(6, 142) <= input(15);
output(6, 143) <= input(37);
output(6, 144) <= input(1);
output(6, 145) <= input(2);
output(6, 146) <= input(3);
output(6, 147) <= input(4);
output(6, 148) <= input(5);
output(6, 149) <= input(6);
output(6, 150) <= input(7);
output(6, 151) <= input(8);
output(6, 152) <= input(9);
output(6, 153) <= input(10);
output(6, 154) <= input(11);
output(6, 155) <= input(12);
output(6, 156) <= input(13);
output(6, 157) <= input(14);
output(6, 158) <= input(15);
output(6, 159) <= input(37);
output(6, 160) <= input(18);
output(6, 161) <= input(19);
output(6, 162) <= input(20);
output(6, 163) <= input(21);
output(6, 164) <= input(22);
output(6, 165) <= input(23);
output(6, 166) <= input(24);
output(6, 167) <= input(25);
output(6, 168) <= input(26);
output(6, 169) <= input(27);
output(6, 170) <= input(28);
output(6, 171) <= input(29);
output(6, 172) <= input(30);
output(6, 173) <= input(31);
output(6, 174) <= input(36);
output(6, 175) <= input(38);
output(6, 176) <= input(18);
output(6, 177) <= input(19);
output(6, 178) <= input(20);
output(6, 179) <= input(21);
output(6, 180) <= input(22);
output(6, 181) <= input(23);
output(6, 182) <= input(24);
output(6, 183) <= input(25);
output(6, 184) <= input(26);
output(6, 185) <= input(27);
output(6, 186) <= input(28);
output(6, 187) <= input(29);
output(6, 188) <= input(30);
output(6, 189) <= input(31);
output(6, 190) <= input(36);
output(6, 191) <= input(38);
output(6, 192) <= input(18);
output(6, 193) <= input(19);
output(6, 194) <= input(20);
output(6, 195) <= input(21);
output(6, 196) <= input(22);
output(6, 197) <= input(23);
output(6, 198) <= input(24);
output(6, 199) <= input(25);
output(6, 200) <= input(26);
output(6, 201) <= input(27);
output(6, 202) <= input(28);
output(6, 203) <= input(29);
output(6, 204) <= input(30);
output(6, 205) <= input(31);
output(6, 206) <= input(36);
output(6, 207) <= input(38);
output(6, 208) <= input(18);
output(6, 209) <= input(19);
output(6, 210) <= input(20);
output(6, 211) <= input(21);
output(6, 212) <= input(22);
output(6, 213) <= input(23);
output(6, 214) <= input(24);
output(6, 215) <= input(25);
output(6, 216) <= input(26);
output(6, 217) <= input(27);
output(6, 218) <= input(28);
output(6, 219) <= input(29);
output(6, 220) <= input(30);
output(6, 221) <= input(31);
output(6, 222) <= input(36);
output(6, 223) <= input(38);
output(6, 224) <= input(18);
output(6, 225) <= input(19);
output(6, 226) <= input(20);
output(6, 227) <= input(21);
output(6, 228) <= input(22);
output(6, 229) <= input(23);
output(6, 230) <= input(24);
output(6, 231) <= input(25);
output(6, 232) <= input(26);
output(6, 233) <= input(27);
output(6, 234) <= input(28);
output(6, 235) <= input(29);
output(6, 236) <= input(30);
output(6, 237) <= input(31);
output(6, 238) <= input(36);
output(6, 239) <= input(38);
output(6, 240) <= input(2);
output(6, 241) <= input(3);
output(6, 242) <= input(4);
output(6, 243) <= input(5);
output(6, 244) <= input(6);
output(6, 245) <= input(7);
output(6, 246) <= input(8);
output(6, 247) <= input(9);
output(6, 248) <= input(10);
output(6, 249) <= input(11);
output(6, 250) <= input(12);
output(6, 251) <= input(13);
output(6, 252) <= input(14);
output(6, 253) <= input(15);
output(6, 254) <= input(37);
output(6, 255) <= input(39);
output(7, 0) <= input(17);
output(7, 1) <= input(18);
output(7, 2) <= input(19);
output(7, 3) <= input(20);
output(7, 4) <= input(21);
output(7, 5) <= input(22);
output(7, 6) <= input(23);
output(7, 7) <= input(24);
output(7, 8) <= input(25);
output(7, 9) <= input(26);
output(7, 10) <= input(27);
output(7, 11) <= input(28);
output(7, 12) <= input(29);
output(7, 13) <= input(30);
output(7, 14) <= input(31);
output(7, 15) <= input(36);
output(7, 16) <= input(17);
output(7, 17) <= input(18);
output(7, 18) <= input(19);
output(7, 19) <= input(20);
output(7, 20) <= input(21);
output(7, 21) <= input(22);
output(7, 22) <= input(23);
output(7, 23) <= input(24);
output(7, 24) <= input(25);
output(7, 25) <= input(26);
output(7, 26) <= input(27);
output(7, 27) <= input(28);
output(7, 28) <= input(29);
output(7, 29) <= input(30);
output(7, 30) <= input(31);
output(7, 31) <= input(36);
output(7, 32) <= input(17);
output(7, 33) <= input(18);
output(7, 34) <= input(19);
output(7, 35) <= input(20);
output(7, 36) <= input(21);
output(7, 37) <= input(22);
output(7, 38) <= input(23);
output(7, 39) <= input(24);
output(7, 40) <= input(25);
output(7, 41) <= input(26);
output(7, 42) <= input(27);
output(7, 43) <= input(28);
output(7, 44) <= input(29);
output(7, 45) <= input(30);
output(7, 46) <= input(31);
output(7, 47) <= input(36);
output(7, 48) <= input(1);
output(7, 49) <= input(2);
output(7, 50) <= input(3);
output(7, 51) <= input(4);
output(7, 52) <= input(5);
output(7, 53) <= input(6);
output(7, 54) <= input(7);
output(7, 55) <= input(8);
output(7, 56) <= input(9);
output(7, 57) <= input(10);
output(7, 58) <= input(11);
output(7, 59) <= input(12);
output(7, 60) <= input(13);
output(7, 61) <= input(14);
output(7, 62) <= input(15);
output(7, 63) <= input(37);
output(7, 64) <= input(1);
output(7, 65) <= input(2);
output(7, 66) <= input(3);
output(7, 67) <= input(4);
output(7, 68) <= input(5);
output(7, 69) <= input(6);
output(7, 70) <= input(7);
output(7, 71) <= input(8);
output(7, 72) <= input(9);
output(7, 73) <= input(10);
output(7, 74) <= input(11);
output(7, 75) <= input(12);
output(7, 76) <= input(13);
output(7, 77) <= input(14);
output(7, 78) <= input(15);
output(7, 79) <= input(37);
output(7, 80) <= input(1);
output(7, 81) <= input(2);
output(7, 82) <= input(3);
output(7, 83) <= input(4);
output(7, 84) <= input(5);
output(7, 85) <= input(6);
output(7, 86) <= input(7);
output(7, 87) <= input(8);
output(7, 88) <= input(9);
output(7, 89) <= input(10);
output(7, 90) <= input(11);
output(7, 91) <= input(12);
output(7, 92) <= input(13);
output(7, 93) <= input(14);
output(7, 94) <= input(15);
output(7, 95) <= input(37);
output(7, 96) <= input(1);
output(7, 97) <= input(2);
output(7, 98) <= input(3);
output(7, 99) <= input(4);
output(7, 100) <= input(5);
output(7, 101) <= input(6);
output(7, 102) <= input(7);
output(7, 103) <= input(8);
output(7, 104) <= input(9);
output(7, 105) <= input(10);
output(7, 106) <= input(11);
output(7, 107) <= input(12);
output(7, 108) <= input(13);
output(7, 109) <= input(14);
output(7, 110) <= input(15);
output(7, 111) <= input(37);
output(7, 112) <= input(18);
output(7, 113) <= input(19);
output(7, 114) <= input(20);
output(7, 115) <= input(21);
output(7, 116) <= input(22);
output(7, 117) <= input(23);
output(7, 118) <= input(24);
output(7, 119) <= input(25);
output(7, 120) <= input(26);
output(7, 121) <= input(27);
output(7, 122) <= input(28);
output(7, 123) <= input(29);
output(7, 124) <= input(30);
output(7, 125) <= input(31);
output(7, 126) <= input(36);
output(7, 127) <= input(38);
output(7, 128) <= input(18);
output(7, 129) <= input(19);
output(7, 130) <= input(20);
output(7, 131) <= input(21);
output(7, 132) <= input(22);
output(7, 133) <= input(23);
output(7, 134) <= input(24);
output(7, 135) <= input(25);
output(7, 136) <= input(26);
output(7, 137) <= input(27);
output(7, 138) <= input(28);
output(7, 139) <= input(29);
output(7, 140) <= input(30);
output(7, 141) <= input(31);
output(7, 142) <= input(36);
output(7, 143) <= input(38);
output(7, 144) <= input(18);
output(7, 145) <= input(19);
output(7, 146) <= input(20);
output(7, 147) <= input(21);
output(7, 148) <= input(22);
output(7, 149) <= input(23);
output(7, 150) <= input(24);
output(7, 151) <= input(25);
output(7, 152) <= input(26);
output(7, 153) <= input(27);
output(7, 154) <= input(28);
output(7, 155) <= input(29);
output(7, 156) <= input(30);
output(7, 157) <= input(31);
output(7, 158) <= input(36);
output(7, 159) <= input(38);
output(7, 160) <= input(18);
output(7, 161) <= input(19);
output(7, 162) <= input(20);
output(7, 163) <= input(21);
output(7, 164) <= input(22);
output(7, 165) <= input(23);
output(7, 166) <= input(24);
output(7, 167) <= input(25);
output(7, 168) <= input(26);
output(7, 169) <= input(27);
output(7, 170) <= input(28);
output(7, 171) <= input(29);
output(7, 172) <= input(30);
output(7, 173) <= input(31);
output(7, 174) <= input(36);
output(7, 175) <= input(38);
output(7, 176) <= input(2);
output(7, 177) <= input(3);
output(7, 178) <= input(4);
output(7, 179) <= input(5);
output(7, 180) <= input(6);
output(7, 181) <= input(7);
output(7, 182) <= input(8);
output(7, 183) <= input(9);
output(7, 184) <= input(10);
output(7, 185) <= input(11);
output(7, 186) <= input(12);
output(7, 187) <= input(13);
output(7, 188) <= input(14);
output(7, 189) <= input(15);
output(7, 190) <= input(37);
output(7, 191) <= input(39);
output(7, 192) <= input(2);
output(7, 193) <= input(3);
output(7, 194) <= input(4);
output(7, 195) <= input(5);
output(7, 196) <= input(6);
output(7, 197) <= input(7);
output(7, 198) <= input(8);
output(7, 199) <= input(9);
output(7, 200) <= input(10);
output(7, 201) <= input(11);
output(7, 202) <= input(12);
output(7, 203) <= input(13);
output(7, 204) <= input(14);
output(7, 205) <= input(15);
output(7, 206) <= input(37);
output(7, 207) <= input(39);
output(7, 208) <= input(2);
output(7, 209) <= input(3);
output(7, 210) <= input(4);
output(7, 211) <= input(5);
output(7, 212) <= input(6);
output(7, 213) <= input(7);
output(7, 214) <= input(8);
output(7, 215) <= input(9);
output(7, 216) <= input(10);
output(7, 217) <= input(11);
output(7, 218) <= input(12);
output(7, 219) <= input(13);
output(7, 220) <= input(14);
output(7, 221) <= input(15);
output(7, 222) <= input(37);
output(7, 223) <= input(39);
output(7, 224) <= input(2);
output(7, 225) <= input(3);
output(7, 226) <= input(4);
output(7, 227) <= input(5);
output(7, 228) <= input(6);
output(7, 229) <= input(7);
output(7, 230) <= input(8);
output(7, 231) <= input(9);
output(7, 232) <= input(10);
output(7, 233) <= input(11);
output(7, 234) <= input(12);
output(7, 235) <= input(13);
output(7, 236) <= input(14);
output(7, 237) <= input(15);
output(7, 238) <= input(37);
output(7, 239) <= input(39);
output(7, 240) <= input(19);
output(7, 241) <= input(20);
output(7, 242) <= input(21);
output(7, 243) <= input(22);
output(7, 244) <= input(23);
output(7, 245) <= input(24);
output(7, 246) <= input(25);
output(7, 247) <= input(26);
output(7, 248) <= input(27);
output(7, 249) <= input(28);
output(7, 250) <= input(29);
output(7, 251) <= input(30);
output(7, 252) <= input(31);
output(7, 253) <= input(36);
output(7, 254) <= input(38);
output(7, 255) <= input(40);
when "1110" =>
output(0, 0) <= input(0);
output(0, 1) <= input(1);
output(0, 2) <= input(2);
output(0, 3) <= input(3);
output(0, 4) <= input(4);
output(0, 5) <= input(5);
output(0, 6) <= input(6);
output(0, 7) <= input(7);
output(0, 8) <= input(8);
output(0, 9) <= input(9);
output(0, 10) <= input(10);
output(0, 11) <= input(11);
output(0, 12) <= input(12);
output(0, 13) <= input(13);
output(0, 14) <= input(14);
output(0, 15) <= input(15);
output(0, 16) <= input(0);
output(0, 17) <= input(1);
output(0, 18) <= input(2);
output(0, 19) <= input(3);
output(0, 20) <= input(4);
output(0, 21) <= input(5);
output(0, 22) <= input(6);
output(0, 23) <= input(7);
output(0, 24) <= input(8);
output(0, 25) <= input(9);
output(0, 26) <= input(10);
output(0, 27) <= input(11);
output(0, 28) <= input(12);
output(0, 29) <= input(13);
output(0, 30) <= input(14);
output(0, 31) <= input(15);
output(0, 32) <= input(16);
output(0, 33) <= input(17);
output(0, 34) <= input(18);
output(0, 35) <= input(19);
output(0, 36) <= input(20);
output(0, 37) <= input(21);
output(0, 38) <= input(22);
output(0, 39) <= input(23);
output(0, 40) <= input(24);
output(0, 41) <= input(25);
output(0, 42) <= input(26);
output(0, 43) <= input(27);
output(0, 44) <= input(28);
output(0, 45) <= input(29);
output(0, 46) <= input(30);
output(0, 47) <= input(31);
output(0, 48) <= input(16);
output(0, 49) <= input(17);
output(0, 50) <= input(18);
output(0, 51) <= input(19);
output(0, 52) <= input(20);
output(0, 53) <= input(21);
output(0, 54) <= input(22);
output(0, 55) <= input(23);
output(0, 56) <= input(24);
output(0, 57) <= input(25);
output(0, 58) <= input(26);
output(0, 59) <= input(27);
output(0, 60) <= input(28);
output(0, 61) <= input(29);
output(0, 62) <= input(30);
output(0, 63) <= input(31);
output(0, 64) <= input(16);
output(0, 65) <= input(17);
output(0, 66) <= input(18);
output(0, 67) <= input(19);
output(0, 68) <= input(20);
output(0, 69) <= input(21);
output(0, 70) <= input(22);
output(0, 71) <= input(23);
output(0, 72) <= input(24);
output(0, 73) <= input(25);
output(0, 74) <= input(26);
output(0, 75) <= input(27);
output(0, 76) <= input(28);
output(0, 77) <= input(29);
output(0, 78) <= input(30);
output(0, 79) <= input(31);
output(0, 80) <= input(1);
output(0, 81) <= input(2);
output(0, 82) <= input(3);
output(0, 83) <= input(4);
output(0, 84) <= input(5);
output(0, 85) <= input(6);
output(0, 86) <= input(7);
output(0, 87) <= input(8);
output(0, 88) <= input(9);
output(0, 89) <= input(10);
output(0, 90) <= input(11);
output(0, 91) <= input(12);
output(0, 92) <= input(13);
output(0, 93) <= input(14);
output(0, 94) <= input(15);
output(0, 95) <= input(32);
output(0, 96) <= input(1);
output(0, 97) <= input(2);
output(0, 98) <= input(3);
output(0, 99) <= input(4);
output(0, 100) <= input(5);
output(0, 101) <= input(6);
output(0, 102) <= input(7);
output(0, 103) <= input(8);
output(0, 104) <= input(9);
output(0, 105) <= input(10);
output(0, 106) <= input(11);
output(0, 107) <= input(12);
output(0, 108) <= input(13);
output(0, 109) <= input(14);
output(0, 110) <= input(15);
output(0, 111) <= input(32);
output(0, 112) <= input(17);
output(0, 113) <= input(18);
output(0, 114) <= input(19);
output(0, 115) <= input(20);
output(0, 116) <= input(21);
output(0, 117) <= input(22);
output(0, 118) <= input(23);
output(0, 119) <= input(24);
output(0, 120) <= input(25);
output(0, 121) <= input(26);
output(0, 122) <= input(27);
output(0, 123) <= input(28);
output(0, 124) <= input(29);
output(0, 125) <= input(30);
output(0, 126) <= input(31);
output(0, 127) <= input(33);
output(0, 128) <= input(17);
output(0, 129) <= input(18);
output(0, 130) <= input(19);
output(0, 131) <= input(20);
output(0, 132) <= input(21);
output(0, 133) <= input(22);
output(0, 134) <= input(23);
output(0, 135) <= input(24);
output(0, 136) <= input(25);
output(0, 137) <= input(26);
output(0, 138) <= input(27);
output(0, 139) <= input(28);
output(0, 140) <= input(29);
output(0, 141) <= input(30);
output(0, 142) <= input(31);
output(0, 143) <= input(33);
output(0, 144) <= input(17);
output(0, 145) <= input(18);
output(0, 146) <= input(19);
output(0, 147) <= input(20);
output(0, 148) <= input(21);
output(0, 149) <= input(22);
output(0, 150) <= input(23);
output(0, 151) <= input(24);
output(0, 152) <= input(25);
output(0, 153) <= input(26);
output(0, 154) <= input(27);
output(0, 155) <= input(28);
output(0, 156) <= input(29);
output(0, 157) <= input(30);
output(0, 158) <= input(31);
output(0, 159) <= input(33);
output(0, 160) <= input(2);
output(0, 161) <= input(3);
output(0, 162) <= input(4);
output(0, 163) <= input(5);
output(0, 164) <= input(6);
output(0, 165) <= input(7);
output(0, 166) <= input(8);
output(0, 167) <= input(9);
output(0, 168) <= input(10);
output(0, 169) <= input(11);
output(0, 170) <= input(12);
output(0, 171) <= input(13);
output(0, 172) <= input(14);
output(0, 173) <= input(15);
output(0, 174) <= input(32);
output(0, 175) <= input(34);
output(0, 176) <= input(2);
output(0, 177) <= input(3);
output(0, 178) <= input(4);
output(0, 179) <= input(5);
output(0, 180) <= input(6);
output(0, 181) <= input(7);
output(0, 182) <= input(8);
output(0, 183) <= input(9);
output(0, 184) <= input(10);
output(0, 185) <= input(11);
output(0, 186) <= input(12);
output(0, 187) <= input(13);
output(0, 188) <= input(14);
output(0, 189) <= input(15);
output(0, 190) <= input(32);
output(0, 191) <= input(34);
output(0, 192) <= input(2);
output(0, 193) <= input(3);
output(0, 194) <= input(4);
output(0, 195) <= input(5);
output(0, 196) <= input(6);
output(0, 197) <= input(7);
output(0, 198) <= input(8);
output(0, 199) <= input(9);
output(0, 200) <= input(10);
output(0, 201) <= input(11);
output(0, 202) <= input(12);
output(0, 203) <= input(13);
output(0, 204) <= input(14);
output(0, 205) <= input(15);
output(0, 206) <= input(32);
output(0, 207) <= input(34);
output(0, 208) <= input(18);
output(0, 209) <= input(19);
output(0, 210) <= input(20);
output(0, 211) <= input(21);
output(0, 212) <= input(22);
output(0, 213) <= input(23);
output(0, 214) <= input(24);
output(0, 215) <= input(25);
output(0, 216) <= input(26);
output(0, 217) <= input(27);
output(0, 218) <= input(28);
output(0, 219) <= input(29);
output(0, 220) <= input(30);
output(0, 221) <= input(31);
output(0, 222) <= input(33);
output(0, 223) <= input(35);
output(0, 224) <= input(18);
output(0, 225) <= input(19);
output(0, 226) <= input(20);
output(0, 227) <= input(21);
output(0, 228) <= input(22);
output(0, 229) <= input(23);
output(0, 230) <= input(24);
output(0, 231) <= input(25);
output(0, 232) <= input(26);
output(0, 233) <= input(27);
output(0, 234) <= input(28);
output(0, 235) <= input(29);
output(0, 236) <= input(30);
output(0, 237) <= input(31);
output(0, 238) <= input(33);
output(0, 239) <= input(35);
output(0, 240) <= input(3);
output(0, 241) <= input(4);
output(0, 242) <= input(5);
output(0, 243) <= input(6);
output(0, 244) <= input(7);
output(0, 245) <= input(8);
output(0, 246) <= input(9);
output(0, 247) <= input(10);
output(0, 248) <= input(11);
output(0, 249) <= input(12);
output(0, 250) <= input(13);
output(0, 251) <= input(14);
output(0, 252) <= input(15);
output(0, 253) <= input(32);
output(0, 254) <= input(34);
output(0, 255) <= input(36);
output(1, 0) <= input(0);
output(1, 1) <= input(1);
output(1, 2) <= input(2);
output(1, 3) <= input(3);
output(1, 4) <= input(4);
output(1, 5) <= input(5);
output(1, 6) <= input(6);
output(1, 7) <= input(7);
output(1, 8) <= input(8);
output(1, 9) <= input(9);
output(1, 10) <= input(10);
output(1, 11) <= input(11);
output(1, 12) <= input(12);
output(1, 13) <= input(13);
output(1, 14) <= input(14);
output(1, 15) <= input(15);
output(1, 16) <= input(16);
output(1, 17) <= input(17);
output(1, 18) <= input(18);
output(1, 19) <= input(19);
output(1, 20) <= input(20);
output(1, 21) <= input(21);
output(1, 22) <= input(22);
output(1, 23) <= input(23);
output(1, 24) <= input(24);
output(1, 25) <= input(25);
output(1, 26) <= input(26);
output(1, 27) <= input(27);
output(1, 28) <= input(28);
output(1, 29) <= input(29);
output(1, 30) <= input(30);
output(1, 31) <= input(31);
output(1, 32) <= input(16);
output(1, 33) <= input(17);
output(1, 34) <= input(18);
output(1, 35) <= input(19);
output(1, 36) <= input(20);
output(1, 37) <= input(21);
output(1, 38) <= input(22);
output(1, 39) <= input(23);
output(1, 40) <= input(24);
output(1, 41) <= input(25);
output(1, 42) <= input(26);
output(1, 43) <= input(27);
output(1, 44) <= input(28);
output(1, 45) <= input(29);
output(1, 46) <= input(30);
output(1, 47) <= input(31);
output(1, 48) <= input(1);
output(1, 49) <= input(2);
output(1, 50) <= input(3);
output(1, 51) <= input(4);
output(1, 52) <= input(5);
output(1, 53) <= input(6);
output(1, 54) <= input(7);
output(1, 55) <= input(8);
output(1, 56) <= input(9);
output(1, 57) <= input(10);
output(1, 58) <= input(11);
output(1, 59) <= input(12);
output(1, 60) <= input(13);
output(1, 61) <= input(14);
output(1, 62) <= input(15);
output(1, 63) <= input(32);
output(1, 64) <= input(1);
output(1, 65) <= input(2);
output(1, 66) <= input(3);
output(1, 67) <= input(4);
output(1, 68) <= input(5);
output(1, 69) <= input(6);
output(1, 70) <= input(7);
output(1, 71) <= input(8);
output(1, 72) <= input(9);
output(1, 73) <= input(10);
output(1, 74) <= input(11);
output(1, 75) <= input(12);
output(1, 76) <= input(13);
output(1, 77) <= input(14);
output(1, 78) <= input(15);
output(1, 79) <= input(32);
output(1, 80) <= input(17);
output(1, 81) <= input(18);
output(1, 82) <= input(19);
output(1, 83) <= input(20);
output(1, 84) <= input(21);
output(1, 85) <= input(22);
output(1, 86) <= input(23);
output(1, 87) <= input(24);
output(1, 88) <= input(25);
output(1, 89) <= input(26);
output(1, 90) <= input(27);
output(1, 91) <= input(28);
output(1, 92) <= input(29);
output(1, 93) <= input(30);
output(1, 94) <= input(31);
output(1, 95) <= input(33);
output(1, 96) <= input(17);
output(1, 97) <= input(18);
output(1, 98) <= input(19);
output(1, 99) <= input(20);
output(1, 100) <= input(21);
output(1, 101) <= input(22);
output(1, 102) <= input(23);
output(1, 103) <= input(24);
output(1, 104) <= input(25);
output(1, 105) <= input(26);
output(1, 106) <= input(27);
output(1, 107) <= input(28);
output(1, 108) <= input(29);
output(1, 109) <= input(30);
output(1, 110) <= input(31);
output(1, 111) <= input(33);
output(1, 112) <= input(2);
output(1, 113) <= input(3);
output(1, 114) <= input(4);
output(1, 115) <= input(5);
output(1, 116) <= input(6);
output(1, 117) <= input(7);
output(1, 118) <= input(8);
output(1, 119) <= input(9);
output(1, 120) <= input(10);
output(1, 121) <= input(11);
output(1, 122) <= input(12);
output(1, 123) <= input(13);
output(1, 124) <= input(14);
output(1, 125) <= input(15);
output(1, 126) <= input(32);
output(1, 127) <= input(34);
output(1, 128) <= input(2);
output(1, 129) <= input(3);
output(1, 130) <= input(4);
output(1, 131) <= input(5);
output(1, 132) <= input(6);
output(1, 133) <= input(7);
output(1, 134) <= input(8);
output(1, 135) <= input(9);
output(1, 136) <= input(10);
output(1, 137) <= input(11);
output(1, 138) <= input(12);
output(1, 139) <= input(13);
output(1, 140) <= input(14);
output(1, 141) <= input(15);
output(1, 142) <= input(32);
output(1, 143) <= input(34);
output(1, 144) <= input(18);
output(1, 145) <= input(19);
output(1, 146) <= input(20);
output(1, 147) <= input(21);
output(1, 148) <= input(22);
output(1, 149) <= input(23);
output(1, 150) <= input(24);
output(1, 151) <= input(25);
output(1, 152) <= input(26);
output(1, 153) <= input(27);
output(1, 154) <= input(28);
output(1, 155) <= input(29);
output(1, 156) <= input(30);
output(1, 157) <= input(31);
output(1, 158) <= input(33);
output(1, 159) <= input(35);
output(1, 160) <= input(18);
output(1, 161) <= input(19);
output(1, 162) <= input(20);
output(1, 163) <= input(21);
output(1, 164) <= input(22);
output(1, 165) <= input(23);
output(1, 166) <= input(24);
output(1, 167) <= input(25);
output(1, 168) <= input(26);
output(1, 169) <= input(27);
output(1, 170) <= input(28);
output(1, 171) <= input(29);
output(1, 172) <= input(30);
output(1, 173) <= input(31);
output(1, 174) <= input(33);
output(1, 175) <= input(35);
output(1, 176) <= input(3);
output(1, 177) <= input(4);
output(1, 178) <= input(5);
output(1, 179) <= input(6);
output(1, 180) <= input(7);
output(1, 181) <= input(8);
output(1, 182) <= input(9);
output(1, 183) <= input(10);
output(1, 184) <= input(11);
output(1, 185) <= input(12);
output(1, 186) <= input(13);
output(1, 187) <= input(14);
output(1, 188) <= input(15);
output(1, 189) <= input(32);
output(1, 190) <= input(34);
output(1, 191) <= input(36);
output(1, 192) <= input(3);
output(1, 193) <= input(4);
output(1, 194) <= input(5);
output(1, 195) <= input(6);
output(1, 196) <= input(7);
output(1, 197) <= input(8);
output(1, 198) <= input(9);
output(1, 199) <= input(10);
output(1, 200) <= input(11);
output(1, 201) <= input(12);
output(1, 202) <= input(13);
output(1, 203) <= input(14);
output(1, 204) <= input(15);
output(1, 205) <= input(32);
output(1, 206) <= input(34);
output(1, 207) <= input(36);
output(1, 208) <= input(19);
output(1, 209) <= input(20);
output(1, 210) <= input(21);
output(1, 211) <= input(22);
output(1, 212) <= input(23);
output(1, 213) <= input(24);
output(1, 214) <= input(25);
output(1, 215) <= input(26);
output(1, 216) <= input(27);
output(1, 217) <= input(28);
output(1, 218) <= input(29);
output(1, 219) <= input(30);
output(1, 220) <= input(31);
output(1, 221) <= input(33);
output(1, 222) <= input(35);
output(1, 223) <= input(37);
output(1, 224) <= input(19);
output(1, 225) <= input(20);
output(1, 226) <= input(21);
output(1, 227) <= input(22);
output(1, 228) <= input(23);
output(1, 229) <= input(24);
output(1, 230) <= input(25);
output(1, 231) <= input(26);
output(1, 232) <= input(27);
output(1, 233) <= input(28);
output(1, 234) <= input(29);
output(1, 235) <= input(30);
output(1, 236) <= input(31);
output(1, 237) <= input(33);
output(1, 238) <= input(35);
output(1, 239) <= input(37);
output(1, 240) <= input(4);
output(1, 241) <= input(5);
output(1, 242) <= input(6);
output(1, 243) <= input(7);
output(1, 244) <= input(8);
output(1, 245) <= input(9);
output(1, 246) <= input(10);
output(1, 247) <= input(11);
output(1, 248) <= input(12);
output(1, 249) <= input(13);
output(1, 250) <= input(14);
output(1, 251) <= input(15);
output(1, 252) <= input(32);
output(1, 253) <= input(34);
output(1, 254) <= input(36);
output(1, 255) <= input(38);
output(2, 0) <= input(0);
output(2, 1) <= input(1);
output(2, 2) <= input(2);
output(2, 3) <= input(3);
output(2, 4) <= input(4);
output(2, 5) <= input(5);
output(2, 6) <= input(6);
output(2, 7) <= input(7);
output(2, 8) <= input(8);
output(2, 9) <= input(9);
output(2, 10) <= input(10);
output(2, 11) <= input(11);
output(2, 12) <= input(12);
output(2, 13) <= input(13);
output(2, 14) <= input(14);
output(2, 15) <= input(15);
output(2, 16) <= input(16);
output(2, 17) <= input(17);
output(2, 18) <= input(18);
output(2, 19) <= input(19);
output(2, 20) <= input(20);
output(2, 21) <= input(21);
output(2, 22) <= input(22);
output(2, 23) <= input(23);
output(2, 24) <= input(24);
output(2, 25) <= input(25);
output(2, 26) <= input(26);
output(2, 27) <= input(27);
output(2, 28) <= input(28);
output(2, 29) <= input(29);
output(2, 30) <= input(30);
output(2, 31) <= input(31);
output(2, 32) <= input(16);
output(2, 33) <= input(17);
output(2, 34) <= input(18);
output(2, 35) <= input(19);
output(2, 36) <= input(20);
output(2, 37) <= input(21);
output(2, 38) <= input(22);
output(2, 39) <= input(23);
output(2, 40) <= input(24);
output(2, 41) <= input(25);
output(2, 42) <= input(26);
output(2, 43) <= input(27);
output(2, 44) <= input(28);
output(2, 45) <= input(29);
output(2, 46) <= input(30);
output(2, 47) <= input(31);
output(2, 48) <= input(1);
output(2, 49) <= input(2);
output(2, 50) <= input(3);
output(2, 51) <= input(4);
output(2, 52) <= input(5);
output(2, 53) <= input(6);
output(2, 54) <= input(7);
output(2, 55) <= input(8);
output(2, 56) <= input(9);
output(2, 57) <= input(10);
output(2, 58) <= input(11);
output(2, 59) <= input(12);
output(2, 60) <= input(13);
output(2, 61) <= input(14);
output(2, 62) <= input(15);
output(2, 63) <= input(32);
output(2, 64) <= input(17);
output(2, 65) <= input(18);
output(2, 66) <= input(19);
output(2, 67) <= input(20);
output(2, 68) <= input(21);
output(2, 69) <= input(22);
output(2, 70) <= input(23);
output(2, 71) <= input(24);
output(2, 72) <= input(25);
output(2, 73) <= input(26);
output(2, 74) <= input(27);
output(2, 75) <= input(28);
output(2, 76) <= input(29);
output(2, 77) <= input(30);
output(2, 78) <= input(31);
output(2, 79) <= input(33);
output(2, 80) <= input(17);
output(2, 81) <= input(18);
output(2, 82) <= input(19);
output(2, 83) <= input(20);
output(2, 84) <= input(21);
output(2, 85) <= input(22);
output(2, 86) <= input(23);
output(2, 87) <= input(24);
output(2, 88) <= input(25);
output(2, 89) <= input(26);
output(2, 90) <= input(27);
output(2, 91) <= input(28);
output(2, 92) <= input(29);
output(2, 93) <= input(30);
output(2, 94) <= input(31);
output(2, 95) <= input(33);
output(2, 96) <= input(2);
output(2, 97) <= input(3);
output(2, 98) <= input(4);
output(2, 99) <= input(5);
output(2, 100) <= input(6);
output(2, 101) <= input(7);
output(2, 102) <= input(8);
output(2, 103) <= input(9);
output(2, 104) <= input(10);
output(2, 105) <= input(11);
output(2, 106) <= input(12);
output(2, 107) <= input(13);
output(2, 108) <= input(14);
output(2, 109) <= input(15);
output(2, 110) <= input(32);
output(2, 111) <= input(34);
output(2, 112) <= input(18);
output(2, 113) <= input(19);
output(2, 114) <= input(20);
output(2, 115) <= input(21);
output(2, 116) <= input(22);
output(2, 117) <= input(23);
output(2, 118) <= input(24);
output(2, 119) <= input(25);
output(2, 120) <= input(26);
output(2, 121) <= input(27);
output(2, 122) <= input(28);
output(2, 123) <= input(29);
output(2, 124) <= input(30);
output(2, 125) <= input(31);
output(2, 126) <= input(33);
output(2, 127) <= input(35);
output(2, 128) <= input(18);
output(2, 129) <= input(19);
output(2, 130) <= input(20);
output(2, 131) <= input(21);
output(2, 132) <= input(22);
output(2, 133) <= input(23);
output(2, 134) <= input(24);
output(2, 135) <= input(25);
output(2, 136) <= input(26);
output(2, 137) <= input(27);
output(2, 138) <= input(28);
output(2, 139) <= input(29);
output(2, 140) <= input(30);
output(2, 141) <= input(31);
output(2, 142) <= input(33);
output(2, 143) <= input(35);
output(2, 144) <= input(3);
output(2, 145) <= input(4);
output(2, 146) <= input(5);
output(2, 147) <= input(6);
output(2, 148) <= input(7);
output(2, 149) <= input(8);
output(2, 150) <= input(9);
output(2, 151) <= input(10);
output(2, 152) <= input(11);
output(2, 153) <= input(12);
output(2, 154) <= input(13);
output(2, 155) <= input(14);
output(2, 156) <= input(15);
output(2, 157) <= input(32);
output(2, 158) <= input(34);
output(2, 159) <= input(36);
output(2, 160) <= input(3);
output(2, 161) <= input(4);
output(2, 162) <= input(5);
output(2, 163) <= input(6);
output(2, 164) <= input(7);
output(2, 165) <= input(8);
output(2, 166) <= input(9);
output(2, 167) <= input(10);
output(2, 168) <= input(11);
output(2, 169) <= input(12);
output(2, 170) <= input(13);
output(2, 171) <= input(14);
output(2, 172) <= input(15);
output(2, 173) <= input(32);
output(2, 174) <= input(34);
output(2, 175) <= input(36);
output(2, 176) <= input(19);
output(2, 177) <= input(20);
output(2, 178) <= input(21);
output(2, 179) <= input(22);
output(2, 180) <= input(23);
output(2, 181) <= input(24);
output(2, 182) <= input(25);
output(2, 183) <= input(26);
output(2, 184) <= input(27);
output(2, 185) <= input(28);
output(2, 186) <= input(29);
output(2, 187) <= input(30);
output(2, 188) <= input(31);
output(2, 189) <= input(33);
output(2, 190) <= input(35);
output(2, 191) <= input(37);
output(2, 192) <= input(4);
output(2, 193) <= input(5);
output(2, 194) <= input(6);
output(2, 195) <= input(7);
output(2, 196) <= input(8);
output(2, 197) <= input(9);
output(2, 198) <= input(10);
output(2, 199) <= input(11);
output(2, 200) <= input(12);
output(2, 201) <= input(13);
output(2, 202) <= input(14);
output(2, 203) <= input(15);
output(2, 204) <= input(32);
output(2, 205) <= input(34);
output(2, 206) <= input(36);
output(2, 207) <= input(38);
output(2, 208) <= input(4);
output(2, 209) <= input(5);
output(2, 210) <= input(6);
output(2, 211) <= input(7);
output(2, 212) <= input(8);
output(2, 213) <= input(9);
output(2, 214) <= input(10);
output(2, 215) <= input(11);
output(2, 216) <= input(12);
output(2, 217) <= input(13);
output(2, 218) <= input(14);
output(2, 219) <= input(15);
output(2, 220) <= input(32);
output(2, 221) <= input(34);
output(2, 222) <= input(36);
output(2, 223) <= input(38);
output(2, 224) <= input(20);
output(2, 225) <= input(21);
output(2, 226) <= input(22);
output(2, 227) <= input(23);
output(2, 228) <= input(24);
output(2, 229) <= input(25);
output(2, 230) <= input(26);
output(2, 231) <= input(27);
output(2, 232) <= input(28);
output(2, 233) <= input(29);
output(2, 234) <= input(30);
output(2, 235) <= input(31);
output(2, 236) <= input(33);
output(2, 237) <= input(35);
output(2, 238) <= input(37);
output(2, 239) <= input(39);
output(2, 240) <= input(5);
output(2, 241) <= input(6);
output(2, 242) <= input(7);
output(2, 243) <= input(8);
output(2, 244) <= input(9);
output(2, 245) <= input(10);
output(2, 246) <= input(11);
output(2, 247) <= input(12);
output(2, 248) <= input(13);
output(2, 249) <= input(14);
output(2, 250) <= input(15);
output(2, 251) <= input(32);
output(2, 252) <= input(34);
output(2, 253) <= input(36);
output(2, 254) <= input(38);
output(2, 255) <= input(40);
output(3, 0) <= input(0);
output(3, 1) <= input(1);
output(3, 2) <= input(2);
output(3, 3) <= input(3);
output(3, 4) <= input(4);
output(3, 5) <= input(5);
output(3, 6) <= input(6);
output(3, 7) <= input(7);
output(3, 8) <= input(8);
output(3, 9) <= input(9);
output(3, 10) <= input(10);
output(3, 11) <= input(11);
output(3, 12) <= input(12);
output(3, 13) <= input(13);
output(3, 14) <= input(14);
output(3, 15) <= input(15);
output(3, 16) <= input(16);
output(3, 17) <= input(17);
output(3, 18) <= input(18);
output(3, 19) <= input(19);
output(3, 20) <= input(20);
output(3, 21) <= input(21);
output(3, 22) <= input(22);
output(3, 23) <= input(23);
output(3, 24) <= input(24);
output(3, 25) <= input(25);
output(3, 26) <= input(26);
output(3, 27) <= input(27);
output(3, 28) <= input(28);
output(3, 29) <= input(29);
output(3, 30) <= input(30);
output(3, 31) <= input(31);
output(3, 32) <= input(1);
output(3, 33) <= input(2);
output(3, 34) <= input(3);
output(3, 35) <= input(4);
output(3, 36) <= input(5);
output(3, 37) <= input(6);
output(3, 38) <= input(7);
output(3, 39) <= input(8);
output(3, 40) <= input(9);
output(3, 41) <= input(10);
output(3, 42) <= input(11);
output(3, 43) <= input(12);
output(3, 44) <= input(13);
output(3, 45) <= input(14);
output(3, 46) <= input(15);
output(3, 47) <= input(32);
output(3, 48) <= input(17);
output(3, 49) <= input(18);
output(3, 50) <= input(19);
output(3, 51) <= input(20);
output(3, 52) <= input(21);
output(3, 53) <= input(22);
output(3, 54) <= input(23);
output(3, 55) <= input(24);
output(3, 56) <= input(25);
output(3, 57) <= input(26);
output(3, 58) <= input(27);
output(3, 59) <= input(28);
output(3, 60) <= input(29);
output(3, 61) <= input(30);
output(3, 62) <= input(31);
output(3, 63) <= input(33);
output(3, 64) <= input(17);
output(3, 65) <= input(18);
output(3, 66) <= input(19);
output(3, 67) <= input(20);
output(3, 68) <= input(21);
output(3, 69) <= input(22);
output(3, 70) <= input(23);
output(3, 71) <= input(24);
output(3, 72) <= input(25);
output(3, 73) <= input(26);
output(3, 74) <= input(27);
output(3, 75) <= input(28);
output(3, 76) <= input(29);
output(3, 77) <= input(30);
output(3, 78) <= input(31);
output(3, 79) <= input(33);
output(3, 80) <= input(2);
output(3, 81) <= input(3);
output(3, 82) <= input(4);
output(3, 83) <= input(5);
output(3, 84) <= input(6);
output(3, 85) <= input(7);
output(3, 86) <= input(8);
output(3, 87) <= input(9);
output(3, 88) <= input(10);
output(3, 89) <= input(11);
output(3, 90) <= input(12);
output(3, 91) <= input(13);
output(3, 92) <= input(14);
output(3, 93) <= input(15);
output(3, 94) <= input(32);
output(3, 95) <= input(34);
output(3, 96) <= input(18);
output(3, 97) <= input(19);
output(3, 98) <= input(20);
output(3, 99) <= input(21);
output(3, 100) <= input(22);
output(3, 101) <= input(23);
output(3, 102) <= input(24);
output(3, 103) <= input(25);
output(3, 104) <= input(26);
output(3, 105) <= input(27);
output(3, 106) <= input(28);
output(3, 107) <= input(29);
output(3, 108) <= input(30);
output(3, 109) <= input(31);
output(3, 110) <= input(33);
output(3, 111) <= input(35);
output(3, 112) <= input(3);
output(3, 113) <= input(4);
output(3, 114) <= input(5);
output(3, 115) <= input(6);
output(3, 116) <= input(7);
output(3, 117) <= input(8);
output(3, 118) <= input(9);
output(3, 119) <= input(10);
output(3, 120) <= input(11);
output(3, 121) <= input(12);
output(3, 122) <= input(13);
output(3, 123) <= input(14);
output(3, 124) <= input(15);
output(3, 125) <= input(32);
output(3, 126) <= input(34);
output(3, 127) <= input(36);
output(3, 128) <= input(3);
output(3, 129) <= input(4);
output(3, 130) <= input(5);
output(3, 131) <= input(6);
output(3, 132) <= input(7);
output(3, 133) <= input(8);
output(3, 134) <= input(9);
output(3, 135) <= input(10);
output(3, 136) <= input(11);
output(3, 137) <= input(12);
output(3, 138) <= input(13);
output(3, 139) <= input(14);
output(3, 140) <= input(15);
output(3, 141) <= input(32);
output(3, 142) <= input(34);
output(3, 143) <= input(36);
output(3, 144) <= input(19);
output(3, 145) <= input(20);
output(3, 146) <= input(21);
output(3, 147) <= input(22);
output(3, 148) <= input(23);
output(3, 149) <= input(24);
output(3, 150) <= input(25);
output(3, 151) <= input(26);
output(3, 152) <= input(27);
output(3, 153) <= input(28);
output(3, 154) <= input(29);
output(3, 155) <= input(30);
output(3, 156) <= input(31);
output(3, 157) <= input(33);
output(3, 158) <= input(35);
output(3, 159) <= input(37);
output(3, 160) <= input(4);
output(3, 161) <= input(5);
output(3, 162) <= input(6);
output(3, 163) <= input(7);
output(3, 164) <= input(8);
output(3, 165) <= input(9);
output(3, 166) <= input(10);
output(3, 167) <= input(11);
output(3, 168) <= input(12);
output(3, 169) <= input(13);
output(3, 170) <= input(14);
output(3, 171) <= input(15);
output(3, 172) <= input(32);
output(3, 173) <= input(34);
output(3, 174) <= input(36);
output(3, 175) <= input(38);
output(3, 176) <= input(20);
output(3, 177) <= input(21);
output(3, 178) <= input(22);
output(3, 179) <= input(23);
output(3, 180) <= input(24);
output(3, 181) <= input(25);
output(3, 182) <= input(26);
output(3, 183) <= input(27);
output(3, 184) <= input(28);
output(3, 185) <= input(29);
output(3, 186) <= input(30);
output(3, 187) <= input(31);
output(3, 188) <= input(33);
output(3, 189) <= input(35);
output(3, 190) <= input(37);
output(3, 191) <= input(39);
output(3, 192) <= input(20);
output(3, 193) <= input(21);
output(3, 194) <= input(22);
output(3, 195) <= input(23);
output(3, 196) <= input(24);
output(3, 197) <= input(25);
output(3, 198) <= input(26);
output(3, 199) <= input(27);
output(3, 200) <= input(28);
output(3, 201) <= input(29);
output(3, 202) <= input(30);
output(3, 203) <= input(31);
output(3, 204) <= input(33);
output(3, 205) <= input(35);
output(3, 206) <= input(37);
output(3, 207) <= input(39);
output(3, 208) <= input(5);
output(3, 209) <= input(6);
output(3, 210) <= input(7);
output(3, 211) <= input(8);
output(3, 212) <= input(9);
output(3, 213) <= input(10);
output(3, 214) <= input(11);
output(3, 215) <= input(12);
output(3, 216) <= input(13);
output(3, 217) <= input(14);
output(3, 218) <= input(15);
output(3, 219) <= input(32);
output(3, 220) <= input(34);
output(3, 221) <= input(36);
output(3, 222) <= input(38);
output(3, 223) <= input(40);
output(3, 224) <= input(21);
output(3, 225) <= input(22);
output(3, 226) <= input(23);
output(3, 227) <= input(24);
output(3, 228) <= input(25);
output(3, 229) <= input(26);
output(3, 230) <= input(27);
output(3, 231) <= input(28);
output(3, 232) <= input(29);
output(3, 233) <= input(30);
output(3, 234) <= input(31);
output(3, 235) <= input(33);
output(3, 236) <= input(35);
output(3, 237) <= input(37);
output(3, 238) <= input(39);
output(3, 239) <= input(41);
output(3, 240) <= input(6);
output(3, 241) <= input(7);
output(3, 242) <= input(8);
output(3, 243) <= input(9);
output(3, 244) <= input(10);
output(3, 245) <= input(11);
output(3, 246) <= input(12);
output(3, 247) <= input(13);
output(3, 248) <= input(14);
output(3, 249) <= input(15);
output(3, 250) <= input(32);
output(3, 251) <= input(34);
output(3, 252) <= input(36);
output(3, 253) <= input(38);
output(3, 254) <= input(40);
output(3, 255) <= input(42);
output(4, 0) <= input(0);
output(4, 1) <= input(1);
output(4, 2) <= input(2);
output(4, 3) <= input(3);
output(4, 4) <= input(4);
output(4, 5) <= input(5);
output(4, 6) <= input(6);
output(4, 7) <= input(7);
output(4, 8) <= input(8);
output(4, 9) <= input(9);
output(4, 10) <= input(10);
output(4, 11) <= input(11);
output(4, 12) <= input(12);
output(4, 13) <= input(13);
output(4, 14) <= input(14);
output(4, 15) <= input(15);
output(4, 16) <= input(16);
output(4, 17) <= input(17);
output(4, 18) <= input(18);
output(4, 19) <= input(19);
output(4, 20) <= input(20);
output(4, 21) <= input(21);
output(4, 22) <= input(22);
output(4, 23) <= input(23);
output(4, 24) <= input(24);
output(4, 25) <= input(25);
output(4, 26) <= input(26);
output(4, 27) <= input(27);
output(4, 28) <= input(28);
output(4, 29) <= input(29);
output(4, 30) <= input(30);
output(4, 31) <= input(31);
output(4, 32) <= input(1);
output(4, 33) <= input(2);
output(4, 34) <= input(3);
output(4, 35) <= input(4);
output(4, 36) <= input(5);
output(4, 37) <= input(6);
output(4, 38) <= input(7);
output(4, 39) <= input(8);
output(4, 40) <= input(9);
output(4, 41) <= input(10);
output(4, 42) <= input(11);
output(4, 43) <= input(12);
output(4, 44) <= input(13);
output(4, 45) <= input(14);
output(4, 46) <= input(15);
output(4, 47) <= input(32);
output(4, 48) <= input(17);
output(4, 49) <= input(18);
output(4, 50) <= input(19);
output(4, 51) <= input(20);
output(4, 52) <= input(21);
output(4, 53) <= input(22);
output(4, 54) <= input(23);
output(4, 55) <= input(24);
output(4, 56) <= input(25);
output(4, 57) <= input(26);
output(4, 58) <= input(27);
output(4, 59) <= input(28);
output(4, 60) <= input(29);
output(4, 61) <= input(30);
output(4, 62) <= input(31);
output(4, 63) <= input(33);
output(4, 64) <= input(2);
output(4, 65) <= input(3);
output(4, 66) <= input(4);
output(4, 67) <= input(5);
output(4, 68) <= input(6);
output(4, 69) <= input(7);
output(4, 70) <= input(8);
output(4, 71) <= input(9);
output(4, 72) <= input(10);
output(4, 73) <= input(11);
output(4, 74) <= input(12);
output(4, 75) <= input(13);
output(4, 76) <= input(14);
output(4, 77) <= input(15);
output(4, 78) <= input(32);
output(4, 79) <= input(34);
output(4, 80) <= input(18);
output(4, 81) <= input(19);
output(4, 82) <= input(20);
output(4, 83) <= input(21);
output(4, 84) <= input(22);
output(4, 85) <= input(23);
output(4, 86) <= input(24);
output(4, 87) <= input(25);
output(4, 88) <= input(26);
output(4, 89) <= input(27);
output(4, 90) <= input(28);
output(4, 91) <= input(29);
output(4, 92) <= input(30);
output(4, 93) <= input(31);
output(4, 94) <= input(33);
output(4, 95) <= input(35);
output(4, 96) <= input(3);
output(4, 97) <= input(4);
output(4, 98) <= input(5);
output(4, 99) <= input(6);
output(4, 100) <= input(7);
output(4, 101) <= input(8);
output(4, 102) <= input(9);
output(4, 103) <= input(10);
output(4, 104) <= input(11);
output(4, 105) <= input(12);
output(4, 106) <= input(13);
output(4, 107) <= input(14);
output(4, 108) <= input(15);
output(4, 109) <= input(32);
output(4, 110) <= input(34);
output(4, 111) <= input(36);
output(4, 112) <= input(19);
output(4, 113) <= input(20);
output(4, 114) <= input(21);
output(4, 115) <= input(22);
output(4, 116) <= input(23);
output(4, 117) <= input(24);
output(4, 118) <= input(25);
output(4, 119) <= input(26);
output(4, 120) <= input(27);
output(4, 121) <= input(28);
output(4, 122) <= input(29);
output(4, 123) <= input(30);
output(4, 124) <= input(31);
output(4, 125) <= input(33);
output(4, 126) <= input(35);
output(4, 127) <= input(37);
output(4, 128) <= input(19);
output(4, 129) <= input(20);
output(4, 130) <= input(21);
output(4, 131) <= input(22);
output(4, 132) <= input(23);
output(4, 133) <= input(24);
output(4, 134) <= input(25);
output(4, 135) <= input(26);
output(4, 136) <= input(27);
output(4, 137) <= input(28);
output(4, 138) <= input(29);
output(4, 139) <= input(30);
output(4, 140) <= input(31);
output(4, 141) <= input(33);
output(4, 142) <= input(35);
output(4, 143) <= input(37);
output(4, 144) <= input(4);
output(4, 145) <= input(5);
output(4, 146) <= input(6);
output(4, 147) <= input(7);
output(4, 148) <= input(8);
output(4, 149) <= input(9);
output(4, 150) <= input(10);
output(4, 151) <= input(11);
output(4, 152) <= input(12);
output(4, 153) <= input(13);
output(4, 154) <= input(14);
output(4, 155) <= input(15);
output(4, 156) <= input(32);
output(4, 157) <= input(34);
output(4, 158) <= input(36);
output(4, 159) <= input(38);
output(4, 160) <= input(20);
output(4, 161) <= input(21);
output(4, 162) <= input(22);
output(4, 163) <= input(23);
output(4, 164) <= input(24);
output(4, 165) <= input(25);
output(4, 166) <= input(26);
output(4, 167) <= input(27);
output(4, 168) <= input(28);
output(4, 169) <= input(29);
output(4, 170) <= input(30);
output(4, 171) <= input(31);
output(4, 172) <= input(33);
output(4, 173) <= input(35);
output(4, 174) <= input(37);
output(4, 175) <= input(39);
output(4, 176) <= input(5);
output(4, 177) <= input(6);
output(4, 178) <= input(7);
output(4, 179) <= input(8);
output(4, 180) <= input(9);
output(4, 181) <= input(10);
output(4, 182) <= input(11);
output(4, 183) <= input(12);
output(4, 184) <= input(13);
output(4, 185) <= input(14);
output(4, 186) <= input(15);
output(4, 187) <= input(32);
output(4, 188) <= input(34);
output(4, 189) <= input(36);
output(4, 190) <= input(38);
output(4, 191) <= input(40);
output(4, 192) <= input(21);
output(4, 193) <= input(22);
output(4, 194) <= input(23);
output(4, 195) <= input(24);
output(4, 196) <= input(25);
output(4, 197) <= input(26);
output(4, 198) <= input(27);
output(4, 199) <= input(28);
output(4, 200) <= input(29);
output(4, 201) <= input(30);
output(4, 202) <= input(31);
output(4, 203) <= input(33);
output(4, 204) <= input(35);
output(4, 205) <= input(37);
output(4, 206) <= input(39);
output(4, 207) <= input(41);
output(4, 208) <= input(6);
output(4, 209) <= input(7);
output(4, 210) <= input(8);
output(4, 211) <= input(9);
output(4, 212) <= input(10);
output(4, 213) <= input(11);
output(4, 214) <= input(12);
output(4, 215) <= input(13);
output(4, 216) <= input(14);
output(4, 217) <= input(15);
output(4, 218) <= input(32);
output(4, 219) <= input(34);
output(4, 220) <= input(36);
output(4, 221) <= input(38);
output(4, 222) <= input(40);
output(4, 223) <= input(42);
output(4, 224) <= input(22);
output(4, 225) <= input(23);
output(4, 226) <= input(24);
output(4, 227) <= input(25);
output(4, 228) <= input(26);
output(4, 229) <= input(27);
output(4, 230) <= input(28);
output(4, 231) <= input(29);
output(4, 232) <= input(30);
output(4, 233) <= input(31);
output(4, 234) <= input(33);
output(4, 235) <= input(35);
output(4, 236) <= input(37);
output(4, 237) <= input(39);
output(4, 238) <= input(41);
output(4, 239) <= input(43);
output(4, 240) <= input(7);
output(4, 241) <= input(8);
output(4, 242) <= input(9);
output(4, 243) <= input(10);
output(4, 244) <= input(11);
output(4, 245) <= input(12);
output(4, 246) <= input(13);
output(4, 247) <= input(14);
output(4, 248) <= input(15);
output(4, 249) <= input(32);
output(4, 250) <= input(34);
output(4, 251) <= input(36);
output(4, 252) <= input(38);
output(4, 253) <= input(40);
output(4, 254) <= input(42);
output(4, 255) <= input(44);
output(5, 0) <= input(16);
output(5, 1) <= input(17);
output(5, 2) <= input(18);
output(5, 3) <= input(19);
output(5, 4) <= input(20);
output(5, 5) <= input(21);
output(5, 6) <= input(22);
output(5, 7) <= input(23);
output(5, 8) <= input(24);
output(5, 9) <= input(25);
output(5, 10) <= input(26);
output(5, 11) <= input(27);
output(5, 12) <= input(28);
output(5, 13) <= input(29);
output(5, 14) <= input(30);
output(5, 15) <= input(31);
output(5, 16) <= input(1);
output(5, 17) <= input(2);
output(5, 18) <= input(3);
output(5, 19) <= input(4);
output(5, 20) <= input(5);
output(5, 21) <= input(6);
output(5, 22) <= input(7);
output(5, 23) <= input(8);
output(5, 24) <= input(9);
output(5, 25) <= input(10);
output(5, 26) <= input(11);
output(5, 27) <= input(12);
output(5, 28) <= input(13);
output(5, 29) <= input(14);
output(5, 30) <= input(15);
output(5, 31) <= input(32);
output(5, 32) <= input(17);
output(5, 33) <= input(18);
output(5, 34) <= input(19);
output(5, 35) <= input(20);
output(5, 36) <= input(21);
output(5, 37) <= input(22);
output(5, 38) <= input(23);
output(5, 39) <= input(24);
output(5, 40) <= input(25);
output(5, 41) <= input(26);
output(5, 42) <= input(27);
output(5, 43) <= input(28);
output(5, 44) <= input(29);
output(5, 45) <= input(30);
output(5, 46) <= input(31);
output(5, 47) <= input(33);
output(5, 48) <= input(2);
output(5, 49) <= input(3);
output(5, 50) <= input(4);
output(5, 51) <= input(5);
output(5, 52) <= input(6);
output(5, 53) <= input(7);
output(5, 54) <= input(8);
output(5, 55) <= input(9);
output(5, 56) <= input(10);
output(5, 57) <= input(11);
output(5, 58) <= input(12);
output(5, 59) <= input(13);
output(5, 60) <= input(14);
output(5, 61) <= input(15);
output(5, 62) <= input(32);
output(5, 63) <= input(34);
output(5, 64) <= input(18);
output(5, 65) <= input(19);
output(5, 66) <= input(20);
output(5, 67) <= input(21);
output(5, 68) <= input(22);
output(5, 69) <= input(23);
output(5, 70) <= input(24);
output(5, 71) <= input(25);
output(5, 72) <= input(26);
output(5, 73) <= input(27);
output(5, 74) <= input(28);
output(5, 75) <= input(29);
output(5, 76) <= input(30);
output(5, 77) <= input(31);
output(5, 78) <= input(33);
output(5, 79) <= input(35);
output(5, 80) <= input(3);
output(5, 81) <= input(4);
output(5, 82) <= input(5);
output(5, 83) <= input(6);
output(5, 84) <= input(7);
output(5, 85) <= input(8);
output(5, 86) <= input(9);
output(5, 87) <= input(10);
output(5, 88) <= input(11);
output(5, 89) <= input(12);
output(5, 90) <= input(13);
output(5, 91) <= input(14);
output(5, 92) <= input(15);
output(5, 93) <= input(32);
output(5, 94) <= input(34);
output(5, 95) <= input(36);
output(5, 96) <= input(19);
output(5, 97) <= input(20);
output(5, 98) <= input(21);
output(5, 99) <= input(22);
output(5, 100) <= input(23);
output(5, 101) <= input(24);
output(5, 102) <= input(25);
output(5, 103) <= input(26);
output(5, 104) <= input(27);
output(5, 105) <= input(28);
output(5, 106) <= input(29);
output(5, 107) <= input(30);
output(5, 108) <= input(31);
output(5, 109) <= input(33);
output(5, 110) <= input(35);
output(5, 111) <= input(37);
output(5, 112) <= input(4);
output(5, 113) <= input(5);
output(5, 114) <= input(6);
output(5, 115) <= input(7);
output(5, 116) <= input(8);
output(5, 117) <= input(9);
output(5, 118) <= input(10);
output(5, 119) <= input(11);
output(5, 120) <= input(12);
output(5, 121) <= input(13);
output(5, 122) <= input(14);
output(5, 123) <= input(15);
output(5, 124) <= input(32);
output(5, 125) <= input(34);
output(5, 126) <= input(36);
output(5, 127) <= input(38);
output(5, 128) <= input(20);
output(5, 129) <= input(21);
output(5, 130) <= input(22);
output(5, 131) <= input(23);
output(5, 132) <= input(24);
output(5, 133) <= input(25);
output(5, 134) <= input(26);
output(5, 135) <= input(27);
output(5, 136) <= input(28);
output(5, 137) <= input(29);
output(5, 138) <= input(30);
output(5, 139) <= input(31);
output(5, 140) <= input(33);
output(5, 141) <= input(35);
output(5, 142) <= input(37);
output(5, 143) <= input(39);
output(5, 144) <= input(5);
output(5, 145) <= input(6);
output(5, 146) <= input(7);
output(5, 147) <= input(8);
output(5, 148) <= input(9);
output(5, 149) <= input(10);
output(5, 150) <= input(11);
output(5, 151) <= input(12);
output(5, 152) <= input(13);
output(5, 153) <= input(14);
output(5, 154) <= input(15);
output(5, 155) <= input(32);
output(5, 156) <= input(34);
output(5, 157) <= input(36);
output(5, 158) <= input(38);
output(5, 159) <= input(40);
output(5, 160) <= input(21);
output(5, 161) <= input(22);
output(5, 162) <= input(23);
output(5, 163) <= input(24);
output(5, 164) <= input(25);
output(5, 165) <= input(26);
output(5, 166) <= input(27);
output(5, 167) <= input(28);
output(5, 168) <= input(29);
output(5, 169) <= input(30);
output(5, 170) <= input(31);
output(5, 171) <= input(33);
output(5, 172) <= input(35);
output(5, 173) <= input(37);
output(5, 174) <= input(39);
output(5, 175) <= input(41);
output(5, 176) <= input(6);
output(5, 177) <= input(7);
output(5, 178) <= input(8);
output(5, 179) <= input(9);
output(5, 180) <= input(10);
output(5, 181) <= input(11);
output(5, 182) <= input(12);
output(5, 183) <= input(13);
output(5, 184) <= input(14);
output(5, 185) <= input(15);
output(5, 186) <= input(32);
output(5, 187) <= input(34);
output(5, 188) <= input(36);
output(5, 189) <= input(38);
output(5, 190) <= input(40);
output(5, 191) <= input(42);
output(5, 192) <= input(22);
output(5, 193) <= input(23);
output(5, 194) <= input(24);
output(5, 195) <= input(25);
output(5, 196) <= input(26);
output(5, 197) <= input(27);
output(5, 198) <= input(28);
output(5, 199) <= input(29);
output(5, 200) <= input(30);
output(5, 201) <= input(31);
output(5, 202) <= input(33);
output(5, 203) <= input(35);
output(5, 204) <= input(37);
output(5, 205) <= input(39);
output(5, 206) <= input(41);
output(5, 207) <= input(43);
output(5, 208) <= input(7);
output(5, 209) <= input(8);
output(5, 210) <= input(9);
output(5, 211) <= input(10);
output(5, 212) <= input(11);
output(5, 213) <= input(12);
output(5, 214) <= input(13);
output(5, 215) <= input(14);
output(5, 216) <= input(15);
output(5, 217) <= input(32);
output(5, 218) <= input(34);
output(5, 219) <= input(36);
output(5, 220) <= input(38);
output(5, 221) <= input(40);
output(5, 222) <= input(42);
output(5, 223) <= input(44);
output(5, 224) <= input(23);
output(5, 225) <= input(24);
output(5, 226) <= input(25);
output(5, 227) <= input(26);
output(5, 228) <= input(27);
output(5, 229) <= input(28);
output(5, 230) <= input(29);
output(5, 231) <= input(30);
output(5, 232) <= input(31);
output(5, 233) <= input(33);
output(5, 234) <= input(35);
output(5, 235) <= input(37);
output(5, 236) <= input(39);
output(5, 237) <= input(41);
output(5, 238) <= input(43);
output(5, 239) <= input(45);
output(5, 240) <= input(8);
output(5, 241) <= input(9);
output(5, 242) <= input(10);
output(5, 243) <= input(11);
output(5, 244) <= input(12);
output(5, 245) <= input(13);
output(5, 246) <= input(14);
output(5, 247) <= input(15);
output(5, 248) <= input(32);
output(5, 249) <= input(34);
output(5, 250) <= input(36);
output(5, 251) <= input(38);
output(5, 252) <= input(40);
output(5, 253) <= input(42);
output(5, 254) <= input(44);
output(5, 255) <= input(46);
when "1111" =>
output(0, 0) <= input(0);
output(0, 1) <= input(1);
output(0, 2) <= input(2);
output(0, 3) <= input(3);
output(0, 4) <= input(4);
output(0, 5) <= input(5);
output(0, 6) <= input(6);
output(0, 7) <= input(7);
output(0, 8) <= input(8);
output(0, 9) <= input(9);
output(0, 10) <= input(10);
output(0, 11) <= input(11);
output(0, 12) <= input(12);
output(0, 13) <= input(13);
output(0, 14) <= input(14);
output(0, 15) <= input(15);
output(0, 16) <= input(16);
output(0, 17) <= input(17);
output(0, 18) <= input(18);
output(0, 19) <= input(19);
output(0, 20) <= input(20);
output(0, 21) <= input(21);
output(0, 22) <= input(22);
output(0, 23) <= input(23);
output(0, 24) <= input(24);
output(0, 25) <= input(25);
output(0, 26) <= input(26);
output(0, 27) <= input(27);
output(0, 28) <= input(28);
output(0, 29) <= input(29);
output(0, 30) <= input(30);
output(0, 31) <= input(31);
output(0, 32) <= input(1);
output(0, 33) <= input(2);
output(0, 34) <= input(3);
output(0, 35) <= input(4);
output(0, 36) <= input(5);
output(0, 37) <= input(6);
output(0, 38) <= input(7);
output(0, 39) <= input(8);
output(0, 40) <= input(9);
output(0, 41) <= input(10);
output(0, 42) <= input(11);
output(0, 43) <= input(12);
output(0, 44) <= input(13);
output(0, 45) <= input(14);
output(0, 46) <= input(15);
output(0, 47) <= input(32);
output(0, 48) <= input(17);
output(0, 49) <= input(18);
output(0, 50) <= input(19);
output(0, 51) <= input(20);
output(0, 52) <= input(21);
output(0, 53) <= input(22);
output(0, 54) <= input(23);
output(0, 55) <= input(24);
output(0, 56) <= input(25);
output(0, 57) <= input(26);
output(0, 58) <= input(27);
output(0, 59) <= input(28);
output(0, 60) <= input(29);
output(0, 61) <= input(30);
output(0, 62) <= input(31);
output(0, 63) <= input(33);
output(0, 64) <= input(2);
output(0, 65) <= input(3);
output(0, 66) <= input(4);
output(0, 67) <= input(5);
output(0, 68) <= input(6);
output(0, 69) <= input(7);
output(0, 70) <= input(8);
output(0, 71) <= input(9);
output(0, 72) <= input(10);
output(0, 73) <= input(11);
output(0, 74) <= input(12);
output(0, 75) <= input(13);
output(0, 76) <= input(14);
output(0, 77) <= input(15);
output(0, 78) <= input(32);
output(0, 79) <= input(34);
output(0, 80) <= input(18);
output(0, 81) <= input(19);
output(0, 82) <= input(20);
output(0, 83) <= input(21);
output(0, 84) <= input(22);
output(0, 85) <= input(23);
output(0, 86) <= input(24);
output(0, 87) <= input(25);
output(0, 88) <= input(26);
output(0, 89) <= input(27);
output(0, 90) <= input(28);
output(0, 91) <= input(29);
output(0, 92) <= input(30);
output(0, 93) <= input(31);
output(0, 94) <= input(33);
output(0, 95) <= input(35);
output(0, 96) <= input(3);
output(0, 97) <= input(4);
output(0, 98) <= input(5);
output(0, 99) <= input(6);
output(0, 100) <= input(7);
output(0, 101) <= input(8);
output(0, 102) <= input(9);
output(0, 103) <= input(10);
output(0, 104) <= input(11);
output(0, 105) <= input(12);
output(0, 106) <= input(13);
output(0, 107) <= input(14);
output(0, 108) <= input(15);
output(0, 109) <= input(32);
output(0, 110) <= input(34);
output(0, 111) <= input(36);
output(0, 112) <= input(4);
output(0, 113) <= input(5);
output(0, 114) <= input(6);
output(0, 115) <= input(7);
output(0, 116) <= input(8);
output(0, 117) <= input(9);
output(0, 118) <= input(10);
output(0, 119) <= input(11);
output(0, 120) <= input(12);
output(0, 121) <= input(13);
output(0, 122) <= input(14);
output(0, 123) <= input(15);
output(0, 124) <= input(32);
output(0, 125) <= input(34);
output(0, 126) <= input(36);
output(0, 127) <= input(37);
output(0, 128) <= input(20);
output(0, 129) <= input(21);
output(0, 130) <= input(22);
output(0, 131) <= input(23);
output(0, 132) <= input(24);
output(0, 133) <= input(25);
output(0, 134) <= input(26);
output(0, 135) <= input(27);
output(0, 136) <= input(28);
output(0, 137) <= input(29);
output(0, 138) <= input(30);
output(0, 139) <= input(31);
output(0, 140) <= input(33);
output(0, 141) <= input(35);
output(0, 142) <= input(38);
output(0, 143) <= input(39);
output(0, 144) <= input(5);
output(0, 145) <= input(6);
output(0, 146) <= input(7);
output(0, 147) <= input(8);
output(0, 148) <= input(9);
output(0, 149) <= input(10);
output(0, 150) <= input(11);
output(0, 151) <= input(12);
output(0, 152) <= input(13);
output(0, 153) <= input(14);
output(0, 154) <= input(15);
output(0, 155) <= input(32);
output(0, 156) <= input(34);
output(0, 157) <= input(36);
output(0, 158) <= input(37);
output(0, 159) <= input(40);
output(0, 160) <= input(21);
output(0, 161) <= input(22);
output(0, 162) <= input(23);
output(0, 163) <= input(24);
output(0, 164) <= input(25);
output(0, 165) <= input(26);
output(0, 166) <= input(27);
output(0, 167) <= input(28);
output(0, 168) <= input(29);
output(0, 169) <= input(30);
output(0, 170) <= input(31);
output(0, 171) <= input(33);
output(0, 172) <= input(35);
output(0, 173) <= input(38);
output(0, 174) <= input(39);
output(0, 175) <= input(41);
output(0, 176) <= input(6);
output(0, 177) <= input(7);
output(0, 178) <= input(8);
output(0, 179) <= input(9);
output(0, 180) <= input(10);
output(0, 181) <= input(11);
output(0, 182) <= input(12);
output(0, 183) <= input(13);
output(0, 184) <= input(14);
output(0, 185) <= input(15);
output(0, 186) <= input(32);
output(0, 187) <= input(34);
output(0, 188) <= input(36);
output(0, 189) <= input(37);
output(0, 190) <= input(40);
output(0, 191) <= input(42);
output(0, 192) <= input(22);
output(0, 193) <= input(23);
output(0, 194) <= input(24);
output(0, 195) <= input(25);
output(0, 196) <= input(26);
output(0, 197) <= input(27);
output(0, 198) <= input(28);
output(0, 199) <= input(29);
output(0, 200) <= input(30);
output(0, 201) <= input(31);
output(0, 202) <= input(33);
output(0, 203) <= input(35);
output(0, 204) <= input(38);
output(0, 205) <= input(39);
output(0, 206) <= input(41);
output(0, 207) <= input(43);
output(0, 208) <= input(7);
output(0, 209) <= input(8);
output(0, 210) <= input(9);
output(0, 211) <= input(10);
output(0, 212) <= input(11);
output(0, 213) <= input(12);
output(0, 214) <= input(13);
output(0, 215) <= input(14);
output(0, 216) <= input(15);
output(0, 217) <= input(32);
output(0, 218) <= input(34);
output(0, 219) <= input(36);
output(0, 220) <= input(37);
output(0, 221) <= input(40);
output(0, 222) <= input(42);
output(0, 223) <= input(44);
output(0, 224) <= input(23);
output(0, 225) <= input(24);
output(0, 226) <= input(25);
output(0, 227) <= input(26);
output(0, 228) <= input(27);
output(0, 229) <= input(28);
output(0, 230) <= input(29);
output(0, 231) <= input(30);
output(0, 232) <= input(31);
output(0, 233) <= input(33);
output(0, 234) <= input(35);
output(0, 235) <= input(38);
output(0, 236) <= input(39);
output(0, 237) <= input(41);
output(0, 238) <= input(43);
output(0, 239) <= input(45);
output(0, 240) <= input(24);
output(0, 241) <= input(25);
output(0, 242) <= input(26);
output(0, 243) <= input(27);
output(0, 244) <= input(28);
output(0, 245) <= input(29);
output(0, 246) <= input(30);
output(0, 247) <= input(31);
output(0, 248) <= input(33);
output(0, 249) <= input(35);
output(0, 250) <= input(38);
output(0, 251) <= input(39);
output(0, 252) <= input(41);
output(0, 253) <= input(43);
output(0, 254) <= input(45);
output(0, 255) <= input(46);
output(1, 0) <= input(0);
output(1, 1) <= input(1);
output(1, 2) <= input(2);
output(1, 3) <= input(3);
output(1, 4) <= input(4);
output(1, 5) <= input(5);
output(1, 6) <= input(6);
output(1, 7) <= input(7);
output(1, 8) <= input(8);
output(1, 9) <= input(9);
output(1, 10) <= input(10);
output(1, 11) <= input(11);
output(1, 12) <= input(12);
output(1, 13) <= input(13);
output(1, 14) <= input(14);
output(1, 15) <= input(15);
output(1, 16) <= input(16);
output(1, 17) <= input(17);
output(1, 18) <= input(18);
output(1, 19) <= input(19);
output(1, 20) <= input(20);
output(1, 21) <= input(21);
output(1, 22) <= input(22);
output(1, 23) <= input(23);
output(1, 24) <= input(24);
output(1, 25) <= input(25);
output(1, 26) <= input(26);
output(1, 27) <= input(27);
output(1, 28) <= input(28);
output(1, 29) <= input(29);
output(1, 30) <= input(30);
output(1, 31) <= input(31);
output(1, 32) <= input(1);
output(1, 33) <= input(2);
output(1, 34) <= input(3);
output(1, 35) <= input(4);
output(1, 36) <= input(5);
output(1, 37) <= input(6);
output(1, 38) <= input(7);
output(1, 39) <= input(8);
output(1, 40) <= input(9);
output(1, 41) <= input(10);
output(1, 42) <= input(11);
output(1, 43) <= input(12);
output(1, 44) <= input(13);
output(1, 45) <= input(14);
output(1, 46) <= input(15);
output(1, 47) <= input(32);
output(1, 48) <= input(2);
output(1, 49) <= input(3);
output(1, 50) <= input(4);
output(1, 51) <= input(5);
output(1, 52) <= input(6);
output(1, 53) <= input(7);
output(1, 54) <= input(8);
output(1, 55) <= input(9);
output(1, 56) <= input(10);
output(1, 57) <= input(11);
output(1, 58) <= input(12);
output(1, 59) <= input(13);
output(1, 60) <= input(14);
output(1, 61) <= input(15);
output(1, 62) <= input(32);
output(1, 63) <= input(34);
output(1, 64) <= input(18);
output(1, 65) <= input(19);
output(1, 66) <= input(20);
output(1, 67) <= input(21);
output(1, 68) <= input(22);
output(1, 69) <= input(23);
output(1, 70) <= input(24);
output(1, 71) <= input(25);
output(1, 72) <= input(26);
output(1, 73) <= input(27);
output(1, 74) <= input(28);
output(1, 75) <= input(29);
output(1, 76) <= input(30);
output(1, 77) <= input(31);
output(1, 78) <= input(33);
output(1, 79) <= input(35);
output(1, 80) <= input(3);
output(1, 81) <= input(4);
output(1, 82) <= input(5);
output(1, 83) <= input(6);
output(1, 84) <= input(7);
output(1, 85) <= input(8);
output(1, 86) <= input(9);
output(1, 87) <= input(10);
output(1, 88) <= input(11);
output(1, 89) <= input(12);
output(1, 90) <= input(13);
output(1, 91) <= input(14);
output(1, 92) <= input(15);
output(1, 93) <= input(32);
output(1, 94) <= input(34);
output(1, 95) <= input(36);
output(1, 96) <= input(19);
output(1, 97) <= input(20);
output(1, 98) <= input(21);
output(1, 99) <= input(22);
output(1, 100) <= input(23);
output(1, 101) <= input(24);
output(1, 102) <= input(25);
output(1, 103) <= input(26);
output(1, 104) <= input(27);
output(1, 105) <= input(28);
output(1, 106) <= input(29);
output(1, 107) <= input(30);
output(1, 108) <= input(31);
output(1, 109) <= input(33);
output(1, 110) <= input(35);
output(1, 111) <= input(38);
output(1, 112) <= input(20);
output(1, 113) <= input(21);
output(1, 114) <= input(22);
output(1, 115) <= input(23);
output(1, 116) <= input(24);
output(1, 117) <= input(25);
output(1, 118) <= input(26);
output(1, 119) <= input(27);
output(1, 120) <= input(28);
output(1, 121) <= input(29);
output(1, 122) <= input(30);
output(1, 123) <= input(31);
output(1, 124) <= input(33);
output(1, 125) <= input(35);
output(1, 126) <= input(38);
output(1, 127) <= input(39);
output(1, 128) <= input(5);
output(1, 129) <= input(6);
output(1, 130) <= input(7);
output(1, 131) <= input(8);
output(1, 132) <= input(9);
output(1, 133) <= input(10);
output(1, 134) <= input(11);
output(1, 135) <= input(12);
output(1, 136) <= input(13);
output(1, 137) <= input(14);
output(1, 138) <= input(15);
output(1, 139) <= input(32);
output(1, 140) <= input(34);
output(1, 141) <= input(36);
output(1, 142) <= input(37);
output(1, 143) <= input(40);
output(1, 144) <= input(21);
output(1, 145) <= input(22);
output(1, 146) <= input(23);
output(1, 147) <= input(24);
output(1, 148) <= input(25);
output(1, 149) <= input(26);
output(1, 150) <= input(27);
output(1, 151) <= input(28);
output(1, 152) <= input(29);
output(1, 153) <= input(30);
output(1, 154) <= input(31);
output(1, 155) <= input(33);
output(1, 156) <= input(35);
output(1, 157) <= input(38);
output(1, 158) <= input(39);
output(1, 159) <= input(41);
output(1, 160) <= input(6);
output(1, 161) <= input(7);
output(1, 162) <= input(8);
output(1, 163) <= input(9);
output(1, 164) <= input(10);
output(1, 165) <= input(11);
output(1, 166) <= input(12);
output(1, 167) <= input(13);
output(1, 168) <= input(14);
output(1, 169) <= input(15);
output(1, 170) <= input(32);
output(1, 171) <= input(34);
output(1, 172) <= input(36);
output(1, 173) <= input(37);
output(1, 174) <= input(40);
output(1, 175) <= input(42);
output(1, 176) <= input(7);
output(1, 177) <= input(8);
output(1, 178) <= input(9);
output(1, 179) <= input(10);
output(1, 180) <= input(11);
output(1, 181) <= input(12);
output(1, 182) <= input(13);
output(1, 183) <= input(14);
output(1, 184) <= input(15);
output(1, 185) <= input(32);
output(1, 186) <= input(34);
output(1, 187) <= input(36);
output(1, 188) <= input(37);
output(1, 189) <= input(40);
output(1, 190) <= input(42);
output(1, 191) <= input(44);
output(1, 192) <= input(23);
output(1, 193) <= input(24);
output(1, 194) <= input(25);
output(1, 195) <= input(26);
output(1, 196) <= input(27);
output(1, 197) <= input(28);
output(1, 198) <= input(29);
output(1, 199) <= input(30);
output(1, 200) <= input(31);
output(1, 201) <= input(33);
output(1, 202) <= input(35);
output(1, 203) <= input(38);
output(1, 204) <= input(39);
output(1, 205) <= input(41);
output(1, 206) <= input(43);
output(1, 207) <= input(45);
output(1, 208) <= input(8);
output(1, 209) <= input(9);
output(1, 210) <= input(10);
output(1, 211) <= input(11);
output(1, 212) <= input(12);
output(1, 213) <= input(13);
output(1, 214) <= input(14);
output(1, 215) <= input(15);
output(1, 216) <= input(32);
output(1, 217) <= input(34);
output(1, 218) <= input(36);
output(1, 219) <= input(37);
output(1, 220) <= input(40);
output(1, 221) <= input(42);
output(1, 222) <= input(44);
output(1, 223) <= input(47);
output(1, 224) <= input(24);
output(1, 225) <= input(25);
output(1, 226) <= input(26);
output(1, 227) <= input(27);
output(1, 228) <= input(28);
output(1, 229) <= input(29);
output(1, 230) <= input(30);
output(1, 231) <= input(31);
output(1, 232) <= input(33);
output(1, 233) <= input(35);
output(1, 234) <= input(38);
output(1, 235) <= input(39);
output(1, 236) <= input(41);
output(1, 237) <= input(43);
output(1, 238) <= input(45);
output(1, 239) <= input(46);
output(1, 240) <= input(25);
output(1, 241) <= input(26);
output(1, 242) <= input(27);
output(1, 243) <= input(28);
output(1, 244) <= input(29);
output(1, 245) <= input(30);
output(1, 246) <= input(31);
output(1, 247) <= input(33);
output(1, 248) <= input(35);
output(1, 249) <= input(38);
output(1, 250) <= input(39);
output(1, 251) <= input(41);
output(1, 252) <= input(43);
output(1, 253) <= input(45);
output(1, 254) <= input(46);
output(1, 255) <= input(48);
output(2, 0) <= input(0);
output(2, 1) <= input(1);
output(2, 2) <= input(2);
output(2, 3) <= input(3);
output(2, 4) <= input(4);
output(2, 5) <= input(5);
output(2, 6) <= input(6);
output(2, 7) <= input(7);
output(2, 8) <= input(8);
output(2, 9) <= input(9);
output(2, 10) <= input(10);
output(2, 11) <= input(11);
output(2, 12) <= input(12);
output(2, 13) <= input(13);
output(2, 14) <= input(14);
output(2, 15) <= input(15);
output(2, 16) <= input(16);
output(2, 17) <= input(17);
output(2, 18) <= input(18);
output(2, 19) <= input(19);
output(2, 20) <= input(20);
output(2, 21) <= input(21);
output(2, 22) <= input(22);
output(2, 23) <= input(23);
output(2, 24) <= input(24);
output(2, 25) <= input(25);
output(2, 26) <= input(26);
output(2, 27) <= input(27);
output(2, 28) <= input(28);
output(2, 29) <= input(29);
output(2, 30) <= input(30);
output(2, 31) <= input(31);
output(2, 32) <= input(17);
output(2, 33) <= input(18);
output(2, 34) <= input(19);
output(2, 35) <= input(20);
output(2, 36) <= input(21);
output(2, 37) <= input(22);
output(2, 38) <= input(23);
output(2, 39) <= input(24);
output(2, 40) <= input(25);
output(2, 41) <= input(26);
output(2, 42) <= input(27);
output(2, 43) <= input(28);
output(2, 44) <= input(29);
output(2, 45) <= input(30);
output(2, 46) <= input(31);
output(2, 47) <= input(33);
output(2, 48) <= input(2);
output(2, 49) <= input(3);
output(2, 50) <= input(4);
output(2, 51) <= input(5);
output(2, 52) <= input(6);
output(2, 53) <= input(7);
output(2, 54) <= input(8);
output(2, 55) <= input(9);
output(2, 56) <= input(10);
output(2, 57) <= input(11);
output(2, 58) <= input(12);
output(2, 59) <= input(13);
output(2, 60) <= input(14);
output(2, 61) <= input(15);
output(2, 62) <= input(32);
output(2, 63) <= input(34);
output(2, 64) <= input(3);
output(2, 65) <= input(4);
output(2, 66) <= input(5);
output(2, 67) <= input(6);
output(2, 68) <= input(7);
output(2, 69) <= input(8);
output(2, 70) <= input(9);
output(2, 71) <= input(10);
output(2, 72) <= input(11);
output(2, 73) <= input(12);
output(2, 74) <= input(13);
output(2, 75) <= input(14);
output(2, 76) <= input(15);
output(2, 77) <= input(32);
output(2, 78) <= input(34);
output(2, 79) <= input(36);
output(2, 80) <= input(19);
output(2, 81) <= input(20);
output(2, 82) <= input(21);
output(2, 83) <= input(22);
output(2, 84) <= input(23);
output(2, 85) <= input(24);
output(2, 86) <= input(25);
output(2, 87) <= input(26);
output(2, 88) <= input(27);
output(2, 89) <= input(28);
output(2, 90) <= input(29);
output(2, 91) <= input(30);
output(2, 92) <= input(31);
output(2, 93) <= input(33);
output(2, 94) <= input(35);
output(2, 95) <= input(38);
output(2, 96) <= input(20);
output(2, 97) <= input(21);
output(2, 98) <= input(22);
output(2, 99) <= input(23);
output(2, 100) <= input(24);
output(2, 101) <= input(25);
output(2, 102) <= input(26);
output(2, 103) <= input(27);
output(2, 104) <= input(28);
output(2, 105) <= input(29);
output(2, 106) <= input(30);
output(2, 107) <= input(31);
output(2, 108) <= input(33);
output(2, 109) <= input(35);
output(2, 110) <= input(38);
output(2, 111) <= input(39);
output(2, 112) <= input(5);
output(2, 113) <= input(6);
output(2, 114) <= input(7);
output(2, 115) <= input(8);
output(2, 116) <= input(9);
output(2, 117) <= input(10);
output(2, 118) <= input(11);
output(2, 119) <= input(12);
output(2, 120) <= input(13);
output(2, 121) <= input(14);
output(2, 122) <= input(15);
output(2, 123) <= input(32);
output(2, 124) <= input(34);
output(2, 125) <= input(36);
output(2, 126) <= input(37);
output(2, 127) <= input(40);
output(2, 128) <= input(21);
output(2, 129) <= input(22);
output(2, 130) <= input(23);
output(2, 131) <= input(24);
output(2, 132) <= input(25);
output(2, 133) <= input(26);
output(2, 134) <= input(27);
output(2, 135) <= input(28);
output(2, 136) <= input(29);
output(2, 137) <= input(30);
output(2, 138) <= input(31);
output(2, 139) <= input(33);
output(2, 140) <= input(35);
output(2, 141) <= input(38);
output(2, 142) <= input(39);
output(2, 143) <= input(41);
output(2, 144) <= input(22);
output(2, 145) <= input(23);
output(2, 146) <= input(24);
output(2, 147) <= input(25);
output(2, 148) <= input(26);
output(2, 149) <= input(27);
output(2, 150) <= input(28);
output(2, 151) <= input(29);
output(2, 152) <= input(30);
output(2, 153) <= input(31);
output(2, 154) <= input(33);
output(2, 155) <= input(35);
output(2, 156) <= input(38);
output(2, 157) <= input(39);
output(2, 158) <= input(41);
output(2, 159) <= input(43);
output(2, 160) <= input(7);
output(2, 161) <= input(8);
output(2, 162) <= input(9);
output(2, 163) <= input(10);
output(2, 164) <= input(11);
output(2, 165) <= input(12);
output(2, 166) <= input(13);
output(2, 167) <= input(14);
output(2, 168) <= input(15);
output(2, 169) <= input(32);
output(2, 170) <= input(34);
output(2, 171) <= input(36);
output(2, 172) <= input(37);
output(2, 173) <= input(40);
output(2, 174) <= input(42);
output(2, 175) <= input(44);
output(2, 176) <= input(8);
output(2, 177) <= input(9);
output(2, 178) <= input(10);
output(2, 179) <= input(11);
output(2, 180) <= input(12);
output(2, 181) <= input(13);
output(2, 182) <= input(14);
output(2, 183) <= input(15);
output(2, 184) <= input(32);
output(2, 185) <= input(34);
output(2, 186) <= input(36);
output(2, 187) <= input(37);
output(2, 188) <= input(40);
output(2, 189) <= input(42);
output(2, 190) <= input(44);
output(2, 191) <= input(47);
output(2, 192) <= input(24);
output(2, 193) <= input(25);
output(2, 194) <= input(26);
output(2, 195) <= input(27);
output(2, 196) <= input(28);
output(2, 197) <= input(29);
output(2, 198) <= input(30);
output(2, 199) <= input(31);
output(2, 200) <= input(33);
output(2, 201) <= input(35);
output(2, 202) <= input(38);
output(2, 203) <= input(39);
output(2, 204) <= input(41);
output(2, 205) <= input(43);
output(2, 206) <= input(45);
output(2, 207) <= input(46);
output(2, 208) <= input(25);
output(2, 209) <= input(26);
output(2, 210) <= input(27);
output(2, 211) <= input(28);
output(2, 212) <= input(29);
output(2, 213) <= input(30);
output(2, 214) <= input(31);
output(2, 215) <= input(33);
output(2, 216) <= input(35);
output(2, 217) <= input(38);
output(2, 218) <= input(39);
output(2, 219) <= input(41);
output(2, 220) <= input(43);
output(2, 221) <= input(45);
output(2, 222) <= input(46);
output(2, 223) <= input(48);
output(2, 224) <= input(10);
output(2, 225) <= input(11);
output(2, 226) <= input(12);
output(2, 227) <= input(13);
output(2, 228) <= input(14);
output(2, 229) <= input(15);
output(2, 230) <= input(32);
output(2, 231) <= input(34);
output(2, 232) <= input(36);
output(2, 233) <= input(37);
output(2, 234) <= input(40);
output(2, 235) <= input(42);
output(2, 236) <= input(44);
output(2, 237) <= input(47);
output(2, 238) <= input(49);
output(2, 239) <= input(50);
output(2, 240) <= input(11);
output(2, 241) <= input(12);
output(2, 242) <= input(13);
output(2, 243) <= input(14);
output(2, 244) <= input(15);
output(2, 245) <= input(32);
output(2, 246) <= input(34);
output(2, 247) <= input(36);
output(2, 248) <= input(37);
output(2, 249) <= input(40);
output(2, 250) <= input(42);
output(2, 251) <= input(44);
output(2, 252) <= input(47);
output(2, 253) <= input(49);
output(2, 254) <= input(50);
output(2, 255) <= input(51);
output(3, 0) <= input(0);
output(3, 1) <= input(1);
output(3, 2) <= input(2);
output(3, 3) <= input(3);
output(3, 4) <= input(4);
output(3, 5) <= input(5);
output(3, 6) <= input(6);
output(3, 7) <= input(7);
output(3, 8) <= input(8);
output(3, 9) <= input(9);
output(3, 10) <= input(10);
output(3, 11) <= input(11);
output(3, 12) <= input(12);
output(3, 13) <= input(13);
output(3, 14) <= input(14);
output(3, 15) <= input(15);
output(3, 16) <= input(1);
output(3, 17) <= input(2);
output(3, 18) <= input(3);
output(3, 19) <= input(4);
output(3, 20) <= input(5);
output(3, 21) <= input(6);
output(3, 22) <= input(7);
output(3, 23) <= input(8);
output(3, 24) <= input(9);
output(3, 25) <= input(10);
output(3, 26) <= input(11);
output(3, 27) <= input(12);
output(3, 28) <= input(13);
output(3, 29) <= input(14);
output(3, 30) <= input(15);
output(3, 31) <= input(32);
output(3, 32) <= input(17);
output(3, 33) <= input(18);
output(3, 34) <= input(19);
output(3, 35) <= input(20);
output(3, 36) <= input(21);
output(3, 37) <= input(22);
output(3, 38) <= input(23);
output(3, 39) <= input(24);
output(3, 40) <= input(25);
output(3, 41) <= input(26);
output(3, 42) <= input(27);
output(3, 43) <= input(28);
output(3, 44) <= input(29);
output(3, 45) <= input(30);
output(3, 46) <= input(31);
output(3, 47) <= input(33);
output(3, 48) <= input(18);
output(3, 49) <= input(19);
output(3, 50) <= input(20);
output(3, 51) <= input(21);
output(3, 52) <= input(22);
output(3, 53) <= input(23);
output(3, 54) <= input(24);
output(3, 55) <= input(25);
output(3, 56) <= input(26);
output(3, 57) <= input(27);
output(3, 58) <= input(28);
output(3, 59) <= input(29);
output(3, 60) <= input(30);
output(3, 61) <= input(31);
output(3, 62) <= input(33);
output(3, 63) <= input(35);
output(3, 64) <= input(19);
output(3, 65) <= input(20);
output(3, 66) <= input(21);
output(3, 67) <= input(22);
output(3, 68) <= input(23);
output(3, 69) <= input(24);
output(3, 70) <= input(25);
output(3, 71) <= input(26);
output(3, 72) <= input(27);
output(3, 73) <= input(28);
output(3, 74) <= input(29);
output(3, 75) <= input(30);
output(3, 76) <= input(31);
output(3, 77) <= input(33);
output(3, 78) <= input(35);
output(3, 79) <= input(38);
output(3, 80) <= input(4);
output(3, 81) <= input(5);
output(3, 82) <= input(6);
output(3, 83) <= input(7);
output(3, 84) <= input(8);
output(3, 85) <= input(9);
output(3, 86) <= input(10);
output(3, 87) <= input(11);
output(3, 88) <= input(12);
output(3, 89) <= input(13);
output(3, 90) <= input(14);
output(3, 91) <= input(15);
output(3, 92) <= input(32);
output(3, 93) <= input(34);
output(3, 94) <= input(36);
output(3, 95) <= input(37);
output(3, 96) <= input(5);
output(3, 97) <= input(6);
output(3, 98) <= input(7);
output(3, 99) <= input(8);
output(3, 100) <= input(9);
output(3, 101) <= input(10);
output(3, 102) <= input(11);
output(3, 103) <= input(12);
output(3, 104) <= input(13);
output(3, 105) <= input(14);
output(3, 106) <= input(15);
output(3, 107) <= input(32);
output(3, 108) <= input(34);
output(3, 109) <= input(36);
output(3, 110) <= input(37);
output(3, 111) <= input(40);
output(3, 112) <= input(6);
output(3, 113) <= input(7);
output(3, 114) <= input(8);
output(3, 115) <= input(9);
output(3, 116) <= input(10);
output(3, 117) <= input(11);
output(3, 118) <= input(12);
output(3, 119) <= input(13);
output(3, 120) <= input(14);
output(3, 121) <= input(15);
output(3, 122) <= input(32);
output(3, 123) <= input(34);
output(3, 124) <= input(36);
output(3, 125) <= input(37);
output(3, 126) <= input(40);
output(3, 127) <= input(42);
output(3, 128) <= input(22);
output(3, 129) <= input(23);
output(3, 130) <= input(24);
output(3, 131) <= input(25);
output(3, 132) <= input(26);
output(3, 133) <= input(27);
output(3, 134) <= input(28);
output(3, 135) <= input(29);
output(3, 136) <= input(30);
output(3, 137) <= input(31);
output(3, 138) <= input(33);
output(3, 139) <= input(35);
output(3, 140) <= input(38);
output(3, 141) <= input(39);
output(3, 142) <= input(41);
output(3, 143) <= input(43);
output(3, 144) <= input(23);
output(3, 145) <= input(24);
output(3, 146) <= input(25);
output(3, 147) <= input(26);
output(3, 148) <= input(27);
output(3, 149) <= input(28);
output(3, 150) <= input(29);
output(3, 151) <= input(30);
output(3, 152) <= input(31);
output(3, 153) <= input(33);
output(3, 154) <= input(35);
output(3, 155) <= input(38);
output(3, 156) <= input(39);
output(3, 157) <= input(41);
output(3, 158) <= input(43);
output(3, 159) <= input(45);
output(3, 160) <= input(8);
output(3, 161) <= input(9);
output(3, 162) <= input(10);
output(3, 163) <= input(11);
output(3, 164) <= input(12);
output(3, 165) <= input(13);
output(3, 166) <= input(14);
output(3, 167) <= input(15);
output(3, 168) <= input(32);
output(3, 169) <= input(34);
output(3, 170) <= input(36);
output(3, 171) <= input(37);
output(3, 172) <= input(40);
output(3, 173) <= input(42);
output(3, 174) <= input(44);
output(3, 175) <= input(47);
output(3, 176) <= input(9);
output(3, 177) <= input(10);
output(3, 178) <= input(11);
output(3, 179) <= input(12);
output(3, 180) <= input(13);
output(3, 181) <= input(14);
output(3, 182) <= input(15);
output(3, 183) <= input(32);
output(3, 184) <= input(34);
output(3, 185) <= input(36);
output(3, 186) <= input(37);
output(3, 187) <= input(40);
output(3, 188) <= input(42);
output(3, 189) <= input(44);
output(3, 190) <= input(47);
output(3, 191) <= input(49);
output(3, 192) <= input(10);
output(3, 193) <= input(11);
output(3, 194) <= input(12);
output(3, 195) <= input(13);
output(3, 196) <= input(14);
output(3, 197) <= input(15);
output(3, 198) <= input(32);
output(3, 199) <= input(34);
output(3, 200) <= input(36);
output(3, 201) <= input(37);
output(3, 202) <= input(40);
output(3, 203) <= input(42);
output(3, 204) <= input(44);
output(3, 205) <= input(47);
output(3, 206) <= input(49);
output(3, 207) <= input(50);
output(3, 208) <= input(26);
output(3, 209) <= input(27);
output(3, 210) <= input(28);
output(3, 211) <= input(29);
output(3, 212) <= input(30);
output(3, 213) <= input(31);
output(3, 214) <= input(33);
output(3, 215) <= input(35);
output(3, 216) <= input(38);
output(3, 217) <= input(39);
output(3, 218) <= input(41);
output(3, 219) <= input(43);
output(3, 220) <= input(45);
output(3, 221) <= input(46);
output(3, 222) <= input(48);
output(3, 223) <= input(52);
output(3, 224) <= input(27);
output(3, 225) <= input(28);
output(3, 226) <= input(29);
output(3, 227) <= input(30);
output(3, 228) <= input(31);
output(3, 229) <= input(33);
output(3, 230) <= input(35);
output(3, 231) <= input(38);
output(3, 232) <= input(39);
output(3, 233) <= input(41);
output(3, 234) <= input(43);
output(3, 235) <= input(45);
output(3, 236) <= input(46);
output(3, 237) <= input(48);
output(3, 238) <= input(52);
output(3, 239) <= input(53);
output(3, 240) <= input(28);
output(3, 241) <= input(29);
output(3, 242) <= input(30);
output(3, 243) <= input(31);
output(3, 244) <= input(33);
output(3, 245) <= input(35);
output(3, 246) <= input(38);
output(3, 247) <= input(39);
output(3, 248) <= input(41);
output(3, 249) <= input(43);
output(3, 250) <= input(45);
output(3, 251) <= input(46);
output(3, 252) <= input(48);
output(3, 253) <= input(52);
output(3, 254) <= input(53);
output(3, 255) <= input(54);
output(4, 0) <= input(0);
output(4, 1) <= input(1);
output(4, 2) <= input(2);
output(4, 3) <= input(3);
output(4, 4) <= input(4);
output(4, 5) <= input(5);
output(4, 6) <= input(6);
output(4, 7) <= input(7);
output(4, 8) <= input(8);
output(4, 9) <= input(9);
output(4, 10) <= input(10);
output(4, 11) <= input(11);
output(4, 12) <= input(12);
output(4, 13) <= input(13);
output(4, 14) <= input(14);
output(4, 15) <= input(15);
output(4, 16) <= input(1);
output(4, 17) <= input(2);
output(4, 18) <= input(3);
output(4, 19) <= input(4);
output(4, 20) <= input(5);
output(4, 21) <= input(6);
output(4, 22) <= input(7);
output(4, 23) <= input(8);
output(4, 24) <= input(9);
output(4, 25) <= input(10);
output(4, 26) <= input(11);
output(4, 27) <= input(12);
output(4, 28) <= input(13);
output(4, 29) <= input(14);
output(4, 30) <= input(15);
output(4, 31) <= input(32);
output(4, 32) <= input(2);
output(4, 33) <= input(3);
output(4, 34) <= input(4);
output(4, 35) <= input(5);
output(4, 36) <= input(6);
output(4, 37) <= input(7);
output(4, 38) <= input(8);
output(4, 39) <= input(9);
output(4, 40) <= input(10);
output(4, 41) <= input(11);
output(4, 42) <= input(12);
output(4, 43) <= input(13);
output(4, 44) <= input(14);
output(4, 45) <= input(15);
output(4, 46) <= input(32);
output(4, 47) <= input(34);
output(4, 48) <= input(3);
output(4, 49) <= input(4);
output(4, 50) <= input(5);
output(4, 51) <= input(6);
output(4, 52) <= input(7);
output(4, 53) <= input(8);
output(4, 54) <= input(9);
output(4, 55) <= input(10);
output(4, 56) <= input(11);
output(4, 57) <= input(12);
output(4, 58) <= input(13);
output(4, 59) <= input(14);
output(4, 60) <= input(15);
output(4, 61) <= input(32);
output(4, 62) <= input(34);
output(4, 63) <= input(36);
output(4, 64) <= input(4);
output(4, 65) <= input(5);
output(4, 66) <= input(6);
output(4, 67) <= input(7);
output(4, 68) <= input(8);
output(4, 69) <= input(9);
output(4, 70) <= input(10);
output(4, 71) <= input(11);
output(4, 72) <= input(12);
output(4, 73) <= input(13);
output(4, 74) <= input(14);
output(4, 75) <= input(15);
output(4, 76) <= input(32);
output(4, 77) <= input(34);
output(4, 78) <= input(36);
output(4, 79) <= input(37);
output(4, 80) <= input(20);
output(4, 81) <= input(21);
output(4, 82) <= input(22);
output(4, 83) <= input(23);
output(4, 84) <= input(24);
output(4, 85) <= input(25);
output(4, 86) <= input(26);
output(4, 87) <= input(27);
output(4, 88) <= input(28);
output(4, 89) <= input(29);
output(4, 90) <= input(30);
output(4, 91) <= input(31);
output(4, 92) <= input(33);
output(4, 93) <= input(35);
output(4, 94) <= input(38);
output(4, 95) <= input(39);
output(4, 96) <= input(21);
output(4, 97) <= input(22);
output(4, 98) <= input(23);
output(4, 99) <= input(24);
output(4, 100) <= input(25);
output(4, 101) <= input(26);
output(4, 102) <= input(27);
output(4, 103) <= input(28);
output(4, 104) <= input(29);
output(4, 105) <= input(30);
output(4, 106) <= input(31);
output(4, 107) <= input(33);
output(4, 108) <= input(35);
output(4, 109) <= input(38);
output(4, 110) <= input(39);
output(4, 111) <= input(41);
output(4, 112) <= input(22);
output(4, 113) <= input(23);
output(4, 114) <= input(24);
output(4, 115) <= input(25);
output(4, 116) <= input(26);
output(4, 117) <= input(27);
output(4, 118) <= input(28);
output(4, 119) <= input(29);
output(4, 120) <= input(30);
output(4, 121) <= input(31);
output(4, 122) <= input(33);
output(4, 123) <= input(35);
output(4, 124) <= input(38);
output(4, 125) <= input(39);
output(4, 126) <= input(41);
output(4, 127) <= input(43);
output(4, 128) <= input(23);
output(4, 129) <= input(24);
output(4, 130) <= input(25);
output(4, 131) <= input(26);
output(4, 132) <= input(27);
output(4, 133) <= input(28);
output(4, 134) <= input(29);
output(4, 135) <= input(30);
output(4, 136) <= input(31);
output(4, 137) <= input(33);
output(4, 138) <= input(35);
output(4, 139) <= input(38);
output(4, 140) <= input(39);
output(4, 141) <= input(41);
output(4, 142) <= input(43);
output(4, 143) <= input(45);
output(4, 144) <= input(24);
output(4, 145) <= input(25);
output(4, 146) <= input(26);
output(4, 147) <= input(27);
output(4, 148) <= input(28);
output(4, 149) <= input(29);
output(4, 150) <= input(30);
output(4, 151) <= input(31);
output(4, 152) <= input(33);
output(4, 153) <= input(35);
output(4, 154) <= input(38);
output(4, 155) <= input(39);
output(4, 156) <= input(41);
output(4, 157) <= input(43);
output(4, 158) <= input(45);
output(4, 159) <= input(46);
output(4, 160) <= input(9);
output(4, 161) <= input(10);
output(4, 162) <= input(11);
output(4, 163) <= input(12);
output(4, 164) <= input(13);
output(4, 165) <= input(14);
output(4, 166) <= input(15);
output(4, 167) <= input(32);
output(4, 168) <= input(34);
output(4, 169) <= input(36);
output(4, 170) <= input(37);
output(4, 171) <= input(40);
output(4, 172) <= input(42);
output(4, 173) <= input(44);
output(4, 174) <= input(47);
output(4, 175) <= input(49);
output(4, 176) <= input(10);
output(4, 177) <= input(11);
output(4, 178) <= input(12);
output(4, 179) <= input(13);
output(4, 180) <= input(14);
output(4, 181) <= input(15);
output(4, 182) <= input(32);
output(4, 183) <= input(34);
output(4, 184) <= input(36);
output(4, 185) <= input(37);
output(4, 186) <= input(40);
output(4, 187) <= input(42);
output(4, 188) <= input(44);
output(4, 189) <= input(47);
output(4, 190) <= input(49);
output(4, 191) <= input(50);
output(4, 192) <= input(11);
output(4, 193) <= input(12);
output(4, 194) <= input(13);
output(4, 195) <= input(14);
output(4, 196) <= input(15);
output(4, 197) <= input(32);
output(4, 198) <= input(34);
output(4, 199) <= input(36);
output(4, 200) <= input(37);
output(4, 201) <= input(40);
output(4, 202) <= input(42);
output(4, 203) <= input(44);
output(4, 204) <= input(47);
output(4, 205) <= input(49);
output(4, 206) <= input(50);
output(4, 207) <= input(51);
output(4, 208) <= input(12);
output(4, 209) <= input(13);
output(4, 210) <= input(14);
output(4, 211) <= input(15);
output(4, 212) <= input(32);
output(4, 213) <= input(34);
output(4, 214) <= input(36);
output(4, 215) <= input(37);
output(4, 216) <= input(40);
output(4, 217) <= input(42);
output(4, 218) <= input(44);
output(4, 219) <= input(47);
output(4, 220) <= input(49);
output(4, 221) <= input(50);
output(4, 222) <= input(51);
output(4, 223) <= input(55);
output(4, 224) <= input(13);
output(4, 225) <= input(14);
output(4, 226) <= input(15);
output(4, 227) <= input(32);
output(4, 228) <= input(34);
output(4, 229) <= input(36);
output(4, 230) <= input(37);
output(4, 231) <= input(40);
output(4, 232) <= input(42);
output(4, 233) <= input(44);
output(4, 234) <= input(47);
output(4, 235) <= input(49);
output(4, 236) <= input(50);
output(4, 237) <= input(51);
output(4, 238) <= input(55);
output(4, 239) <= input(56);
output(4, 240) <= input(14);
output(4, 241) <= input(15);
output(4, 242) <= input(32);
output(4, 243) <= input(34);
output(4, 244) <= input(36);
output(4, 245) <= input(37);
output(4, 246) <= input(40);
output(4, 247) <= input(42);
output(4, 248) <= input(44);
output(4, 249) <= input(47);
output(4, 250) <= input(49);
output(4, 251) <= input(50);
output(4, 252) <= input(51);
output(4, 253) <= input(55);
output(4, 254) <= input(56);
output(4, 255) <= input(57);
output(5, 0) <= input(16);
output(5, 1) <= input(17);
output(5, 2) <= input(18);
output(5, 3) <= input(19);
output(5, 4) <= input(20);
output(5, 5) <= input(21);
output(5, 6) <= input(22);
output(5, 7) <= input(23);
output(5, 8) <= input(24);
output(5, 9) <= input(25);
output(5, 10) <= input(26);
output(5, 11) <= input(27);
output(5, 12) <= input(28);
output(5, 13) <= input(29);
output(5, 14) <= input(30);
output(5, 15) <= input(31);
output(5, 16) <= input(17);
output(5, 17) <= input(18);
output(5, 18) <= input(19);
output(5, 19) <= input(20);
output(5, 20) <= input(21);
output(5, 21) <= input(22);
output(5, 22) <= input(23);
output(5, 23) <= input(24);
output(5, 24) <= input(25);
output(5, 25) <= input(26);
output(5, 26) <= input(27);
output(5, 27) <= input(28);
output(5, 28) <= input(29);
output(5, 29) <= input(30);
output(5, 30) <= input(31);
output(5, 31) <= input(33);
output(5, 32) <= input(18);
output(5, 33) <= input(19);
output(5, 34) <= input(20);
output(5, 35) <= input(21);
output(5, 36) <= input(22);
output(5, 37) <= input(23);
output(5, 38) <= input(24);
output(5, 39) <= input(25);
output(5, 40) <= input(26);
output(5, 41) <= input(27);
output(5, 42) <= input(28);
output(5, 43) <= input(29);
output(5, 44) <= input(30);
output(5, 45) <= input(31);
output(5, 46) <= input(33);
output(5, 47) <= input(35);
output(5, 48) <= input(19);
output(5, 49) <= input(20);
output(5, 50) <= input(21);
output(5, 51) <= input(22);
output(5, 52) <= input(23);
output(5, 53) <= input(24);
output(5, 54) <= input(25);
output(5, 55) <= input(26);
output(5, 56) <= input(27);
output(5, 57) <= input(28);
output(5, 58) <= input(29);
output(5, 59) <= input(30);
output(5, 60) <= input(31);
output(5, 61) <= input(33);
output(5, 62) <= input(35);
output(5, 63) <= input(38);
output(5, 64) <= input(20);
output(5, 65) <= input(21);
output(5, 66) <= input(22);
output(5, 67) <= input(23);
output(5, 68) <= input(24);
output(5, 69) <= input(25);
output(5, 70) <= input(26);
output(5, 71) <= input(27);
output(5, 72) <= input(28);
output(5, 73) <= input(29);
output(5, 74) <= input(30);
output(5, 75) <= input(31);
output(5, 76) <= input(33);
output(5, 77) <= input(35);
output(5, 78) <= input(38);
output(5, 79) <= input(39);
output(5, 80) <= input(21);
output(5, 81) <= input(22);
output(5, 82) <= input(23);
output(5, 83) <= input(24);
output(5, 84) <= input(25);
output(5, 85) <= input(26);
output(5, 86) <= input(27);
output(5, 87) <= input(28);
output(5, 88) <= input(29);
output(5, 89) <= input(30);
output(5, 90) <= input(31);
output(5, 91) <= input(33);
output(5, 92) <= input(35);
output(5, 93) <= input(38);
output(5, 94) <= input(39);
output(5, 95) <= input(41);
output(5, 96) <= input(22);
output(5, 97) <= input(23);
output(5, 98) <= input(24);
output(5, 99) <= input(25);
output(5, 100) <= input(26);
output(5, 101) <= input(27);
output(5, 102) <= input(28);
output(5, 103) <= input(29);
output(5, 104) <= input(30);
output(5, 105) <= input(31);
output(5, 106) <= input(33);
output(5, 107) <= input(35);
output(5, 108) <= input(38);
output(5, 109) <= input(39);
output(5, 110) <= input(41);
output(5, 111) <= input(43);
output(5, 112) <= input(23);
output(5, 113) <= input(24);
output(5, 114) <= input(25);
output(5, 115) <= input(26);
output(5, 116) <= input(27);
output(5, 117) <= input(28);
output(5, 118) <= input(29);
output(5, 119) <= input(30);
output(5, 120) <= input(31);
output(5, 121) <= input(33);
output(5, 122) <= input(35);
output(5, 123) <= input(38);
output(5, 124) <= input(39);
output(5, 125) <= input(41);
output(5, 126) <= input(43);
output(5, 127) <= input(45);
output(5, 128) <= input(24);
output(5, 129) <= input(25);
output(5, 130) <= input(26);
output(5, 131) <= input(27);
output(5, 132) <= input(28);
output(5, 133) <= input(29);
output(5, 134) <= input(30);
output(5, 135) <= input(31);
output(5, 136) <= input(33);
output(5, 137) <= input(35);
output(5, 138) <= input(38);
output(5, 139) <= input(39);
output(5, 140) <= input(41);
output(5, 141) <= input(43);
output(5, 142) <= input(45);
output(5, 143) <= input(46);
output(5, 144) <= input(25);
output(5, 145) <= input(26);
output(5, 146) <= input(27);
output(5, 147) <= input(28);
output(5, 148) <= input(29);
output(5, 149) <= input(30);
output(5, 150) <= input(31);
output(5, 151) <= input(33);
output(5, 152) <= input(35);
output(5, 153) <= input(38);
output(5, 154) <= input(39);
output(5, 155) <= input(41);
output(5, 156) <= input(43);
output(5, 157) <= input(45);
output(5, 158) <= input(46);
output(5, 159) <= input(48);
output(5, 160) <= input(26);
output(5, 161) <= input(27);
output(5, 162) <= input(28);
output(5, 163) <= input(29);
output(5, 164) <= input(30);
output(5, 165) <= input(31);
output(5, 166) <= input(33);
output(5, 167) <= input(35);
output(5, 168) <= input(38);
output(5, 169) <= input(39);
output(5, 170) <= input(41);
output(5, 171) <= input(43);
output(5, 172) <= input(45);
output(5, 173) <= input(46);
output(5, 174) <= input(48);
output(5, 175) <= input(52);
output(5, 176) <= input(27);
output(5, 177) <= input(28);
output(5, 178) <= input(29);
output(5, 179) <= input(30);
output(5, 180) <= input(31);
output(5, 181) <= input(33);
output(5, 182) <= input(35);
output(5, 183) <= input(38);
output(5, 184) <= input(39);
output(5, 185) <= input(41);
output(5, 186) <= input(43);
output(5, 187) <= input(45);
output(5, 188) <= input(46);
output(5, 189) <= input(48);
output(5, 190) <= input(52);
output(5, 191) <= input(53);
output(5, 192) <= input(28);
output(5, 193) <= input(29);
output(5, 194) <= input(30);
output(5, 195) <= input(31);
output(5, 196) <= input(33);
output(5, 197) <= input(35);
output(5, 198) <= input(38);
output(5, 199) <= input(39);
output(5, 200) <= input(41);
output(5, 201) <= input(43);
output(5, 202) <= input(45);
output(5, 203) <= input(46);
output(5, 204) <= input(48);
output(5, 205) <= input(52);
output(5, 206) <= input(53);
output(5, 207) <= input(54);
output(5, 208) <= input(29);
output(5, 209) <= input(30);
output(5, 210) <= input(31);
output(5, 211) <= input(33);
output(5, 212) <= input(35);
output(5, 213) <= input(38);
output(5, 214) <= input(39);
output(5, 215) <= input(41);
output(5, 216) <= input(43);
output(5, 217) <= input(45);
output(5, 218) <= input(46);
output(5, 219) <= input(48);
output(5, 220) <= input(52);
output(5, 221) <= input(53);
output(5, 222) <= input(54);
output(5, 223) <= input(58);
output(5, 224) <= input(30);
output(5, 225) <= input(31);
output(5, 226) <= input(33);
output(5, 227) <= input(35);
output(5, 228) <= input(38);
output(5, 229) <= input(39);
output(5, 230) <= input(41);
output(5, 231) <= input(43);
output(5, 232) <= input(45);
output(5, 233) <= input(46);
output(5, 234) <= input(48);
output(5, 235) <= input(52);
output(5, 236) <= input(53);
output(5, 237) <= input(54);
output(5, 238) <= input(58);
output(5, 239) <= input(59);
output(5, 240) <= input(31);
output(5, 241) <= input(33);
output(5, 242) <= input(35);
output(5, 243) <= input(38);
output(5, 244) <= input(39);
output(5, 245) <= input(41);
output(5, 246) <= input(43);
output(5, 247) <= input(45);
output(5, 248) <= input(46);
output(5, 249) <= input(48);
output(5, 250) <= input(52);
output(5, 251) <= input(53);
output(5, 252) <= input(54);
output(5, 253) <= input(58);
output(5, 254) <= input(59);
output(5, 255) <= input(60);
when others => for i in 0 to 7 loop for j in 0 to 255 loop output(i,j) <= "00000000"; end loop; end loop;
end case;
elsif control = "001" then 
case iteration_control is
when "0000" =>
output(0, 0) <= input(0);
output(0, 1) <= input(1);
output(0, 2) <= input(2);
output(0, 3) <= input(3);
output(0, 4) <= input(4);
output(0, 5) <= input(5);
output(0, 6) <= input(6);
output(0, 7) <= input(7);
output(0, 8) <= input(8);
output(0, 9) <= input(9);
output(0, 10) <= input(10);
output(0, 11) <= input(11);
output(0, 12) <= input(12);
output(0, 13) <= input(13);
output(0, 14) <= input(14);
output(0, 15) <= input(15);
output(0, 16) <= input(1);
output(0, 17) <= input(2);
output(0, 18) <= input(3);
output(0, 19) <= input(4);
output(0, 20) <= input(5);
output(0, 21) <= input(6);
output(0, 22) <= input(7);
output(0, 23) <= input(8);
output(0, 24) <= input(9);
output(0, 25) <= input(10);
output(0, 26) <= input(11);
output(0, 27) <= input(12);
output(0, 28) <= input(13);
output(0, 29) <= input(14);
output(0, 30) <= input(15);
output(0, 31) <= input(16);
output(0, 32) <= input(2);
output(0, 33) <= input(3);
output(0, 34) <= input(4);
output(0, 35) <= input(5);
output(0, 36) <= input(6);
output(0, 37) <= input(7);
output(0, 38) <= input(8);
output(0, 39) <= input(9);
output(0, 40) <= input(10);
output(0, 41) <= input(11);
output(0, 42) <= input(12);
output(0, 43) <= input(13);
output(0, 44) <= input(14);
output(0, 45) <= input(15);
output(0, 46) <= input(16);
output(0, 47) <= input(17);
output(0, 48) <= input(3);
output(0, 49) <= input(4);
output(0, 50) <= input(5);
output(0, 51) <= input(6);
output(0, 52) <= input(7);
output(0, 53) <= input(8);
output(0, 54) <= input(9);
output(0, 55) <= input(10);
output(0, 56) <= input(11);
output(0, 57) <= input(12);
output(0, 58) <= input(13);
output(0, 59) <= input(14);
output(0, 60) <= input(15);
output(0, 61) <= input(16);
output(0, 62) <= input(17);
output(0, 63) <= input(18);
output(0, 64) <= input(4);
output(0, 65) <= input(5);
output(0, 66) <= input(6);
output(0, 67) <= input(7);
output(0, 68) <= input(8);
output(0, 69) <= input(9);
output(0, 70) <= input(10);
output(0, 71) <= input(11);
output(0, 72) <= input(12);
output(0, 73) <= input(13);
output(0, 74) <= input(14);
output(0, 75) <= input(15);
output(0, 76) <= input(16);
output(0, 77) <= input(17);
output(0, 78) <= input(18);
output(0, 79) <= input(19);
output(0, 80) <= input(5);
output(0, 81) <= input(6);
output(0, 82) <= input(7);
output(0, 83) <= input(8);
output(0, 84) <= input(9);
output(0, 85) <= input(10);
output(0, 86) <= input(11);
output(0, 87) <= input(12);
output(0, 88) <= input(13);
output(0, 89) <= input(14);
output(0, 90) <= input(15);
output(0, 91) <= input(16);
output(0, 92) <= input(17);
output(0, 93) <= input(18);
output(0, 94) <= input(19);
output(0, 95) <= input(20);
output(0, 96) <= input(6);
output(0, 97) <= input(7);
output(0, 98) <= input(8);
output(0, 99) <= input(9);
output(0, 100) <= input(10);
output(0, 101) <= input(11);
output(0, 102) <= input(12);
output(0, 103) <= input(13);
output(0, 104) <= input(14);
output(0, 105) <= input(15);
output(0, 106) <= input(16);
output(0, 107) <= input(17);
output(0, 108) <= input(18);
output(0, 109) <= input(19);
output(0, 110) <= input(20);
output(0, 111) <= input(21);
output(0, 112) <= input(7);
output(0, 113) <= input(8);
output(0, 114) <= input(9);
output(0, 115) <= input(10);
output(0, 116) <= input(11);
output(0, 117) <= input(12);
output(0, 118) <= input(13);
output(0, 119) <= input(14);
output(0, 120) <= input(15);
output(0, 121) <= input(16);
output(0, 122) <= input(17);
output(0, 123) <= input(18);
output(0, 124) <= input(19);
output(0, 125) <= input(20);
output(0, 126) <= input(21);
output(0, 127) <= input(22);
output(0, 128) <= input(8);
output(0, 129) <= input(9);
output(0, 130) <= input(10);
output(0, 131) <= input(11);
output(0, 132) <= input(12);
output(0, 133) <= input(13);
output(0, 134) <= input(14);
output(0, 135) <= input(15);
output(0, 136) <= input(16);
output(0, 137) <= input(17);
output(0, 138) <= input(18);
output(0, 139) <= input(19);
output(0, 140) <= input(20);
output(0, 141) <= input(21);
output(0, 142) <= input(22);
output(0, 143) <= input(23);
output(0, 144) <= input(9);
output(0, 145) <= input(10);
output(0, 146) <= input(11);
output(0, 147) <= input(12);
output(0, 148) <= input(13);
output(0, 149) <= input(14);
output(0, 150) <= input(15);
output(0, 151) <= input(16);
output(0, 152) <= input(17);
output(0, 153) <= input(18);
output(0, 154) <= input(19);
output(0, 155) <= input(20);
output(0, 156) <= input(21);
output(0, 157) <= input(22);
output(0, 158) <= input(23);
output(0, 159) <= input(24);
output(0, 160) <= input(10);
output(0, 161) <= input(11);
output(0, 162) <= input(12);
output(0, 163) <= input(13);
output(0, 164) <= input(14);
output(0, 165) <= input(15);
output(0, 166) <= input(16);
output(0, 167) <= input(17);
output(0, 168) <= input(18);
output(0, 169) <= input(19);
output(0, 170) <= input(20);
output(0, 171) <= input(21);
output(0, 172) <= input(22);
output(0, 173) <= input(23);
output(0, 174) <= input(24);
output(0, 175) <= input(25);
output(0, 176) <= input(11);
output(0, 177) <= input(12);
output(0, 178) <= input(13);
output(0, 179) <= input(14);
output(0, 180) <= input(15);
output(0, 181) <= input(16);
output(0, 182) <= input(17);
output(0, 183) <= input(18);
output(0, 184) <= input(19);
output(0, 185) <= input(20);
output(0, 186) <= input(21);
output(0, 187) <= input(22);
output(0, 188) <= input(23);
output(0, 189) <= input(24);
output(0, 190) <= input(25);
output(0, 191) <= input(26);
output(0, 192) <= input(12);
output(0, 193) <= input(13);
output(0, 194) <= input(14);
output(0, 195) <= input(15);
output(0, 196) <= input(16);
output(0, 197) <= input(17);
output(0, 198) <= input(18);
output(0, 199) <= input(19);
output(0, 200) <= input(20);
output(0, 201) <= input(21);
output(0, 202) <= input(22);
output(0, 203) <= input(23);
output(0, 204) <= input(24);
output(0, 205) <= input(25);
output(0, 206) <= input(26);
output(0, 207) <= input(27);
output(0, 208) <= input(13);
output(0, 209) <= input(14);
output(0, 210) <= input(15);
output(0, 211) <= input(16);
output(0, 212) <= input(17);
output(0, 213) <= input(18);
output(0, 214) <= input(19);
output(0, 215) <= input(20);
output(0, 216) <= input(21);
output(0, 217) <= input(22);
output(0, 218) <= input(23);
output(0, 219) <= input(24);
output(0, 220) <= input(25);
output(0, 221) <= input(26);
output(0, 222) <= input(27);
output(0, 223) <= input(28);
output(0, 224) <= input(14);
output(0, 225) <= input(15);
output(0, 226) <= input(16);
output(0, 227) <= input(17);
output(0, 228) <= input(18);
output(0, 229) <= input(19);
output(0, 230) <= input(20);
output(0, 231) <= input(21);
output(0, 232) <= input(22);
output(0, 233) <= input(23);
output(0, 234) <= input(24);
output(0, 235) <= input(25);
output(0, 236) <= input(26);
output(0, 237) <= input(27);
output(0, 238) <= input(28);
output(0, 239) <= input(29);
output(0, 240) <= input(15);
output(0, 241) <= input(16);
output(0, 242) <= input(17);
output(0, 243) <= input(18);
output(0, 244) <= input(19);
output(0, 245) <= input(20);
output(0, 246) <= input(21);
output(0, 247) <= input(22);
output(0, 248) <= input(23);
output(0, 249) <= input(24);
output(0, 250) <= input(25);
output(0, 251) <= input(26);
output(0, 252) <= input(27);
output(0, 253) <= input(28);
output(0, 254) <= input(29);
output(0, 255) <= input(30);
output(1, 0) <= input(31);
output(1, 1) <= input(32);
output(1, 2) <= input(33);
output(1, 3) <= input(34);
output(1, 4) <= input(35);
output(1, 5) <= input(36);
output(1, 6) <= input(37);
output(1, 7) <= input(38);
output(1, 8) <= input(39);
output(1, 9) <= input(40);
output(1, 10) <= input(41);
output(1, 11) <= input(42);
output(1, 12) <= input(43);
output(1, 13) <= input(44);
output(1, 14) <= input(45);
output(1, 15) <= input(46);
output(1, 16) <= input(32);
output(1, 17) <= input(33);
output(1, 18) <= input(34);
output(1, 19) <= input(35);
output(1, 20) <= input(36);
output(1, 21) <= input(37);
output(1, 22) <= input(38);
output(1, 23) <= input(39);
output(1, 24) <= input(40);
output(1, 25) <= input(41);
output(1, 26) <= input(42);
output(1, 27) <= input(43);
output(1, 28) <= input(44);
output(1, 29) <= input(45);
output(1, 30) <= input(46);
output(1, 31) <= input(47);
output(1, 32) <= input(33);
output(1, 33) <= input(34);
output(1, 34) <= input(35);
output(1, 35) <= input(36);
output(1, 36) <= input(37);
output(1, 37) <= input(38);
output(1, 38) <= input(39);
output(1, 39) <= input(40);
output(1, 40) <= input(41);
output(1, 41) <= input(42);
output(1, 42) <= input(43);
output(1, 43) <= input(44);
output(1, 44) <= input(45);
output(1, 45) <= input(46);
output(1, 46) <= input(47);
output(1, 47) <= input(48);
output(1, 48) <= input(34);
output(1, 49) <= input(35);
output(1, 50) <= input(36);
output(1, 51) <= input(37);
output(1, 52) <= input(38);
output(1, 53) <= input(39);
output(1, 54) <= input(40);
output(1, 55) <= input(41);
output(1, 56) <= input(42);
output(1, 57) <= input(43);
output(1, 58) <= input(44);
output(1, 59) <= input(45);
output(1, 60) <= input(46);
output(1, 61) <= input(47);
output(1, 62) <= input(48);
output(1, 63) <= input(49);
output(1, 64) <= input(35);
output(1, 65) <= input(36);
output(1, 66) <= input(37);
output(1, 67) <= input(38);
output(1, 68) <= input(39);
output(1, 69) <= input(40);
output(1, 70) <= input(41);
output(1, 71) <= input(42);
output(1, 72) <= input(43);
output(1, 73) <= input(44);
output(1, 74) <= input(45);
output(1, 75) <= input(46);
output(1, 76) <= input(47);
output(1, 77) <= input(48);
output(1, 78) <= input(49);
output(1, 79) <= input(50);
output(1, 80) <= input(4);
output(1, 81) <= input(5);
output(1, 82) <= input(6);
output(1, 83) <= input(7);
output(1, 84) <= input(8);
output(1, 85) <= input(9);
output(1, 86) <= input(10);
output(1, 87) <= input(11);
output(1, 88) <= input(12);
output(1, 89) <= input(13);
output(1, 90) <= input(14);
output(1, 91) <= input(15);
output(1, 92) <= input(16);
output(1, 93) <= input(17);
output(1, 94) <= input(18);
output(1, 95) <= input(19);
output(1, 96) <= input(5);
output(1, 97) <= input(6);
output(1, 98) <= input(7);
output(1, 99) <= input(8);
output(1, 100) <= input(9);
output(1, 101) <= input(10);
output(1, 102) <= input(11);
output(1, 103) <= input(12);
output(1, 104) <= input(13);
output(1, 105) <= input(14);
output(1, 106) <= input(15);
output(1, 107) <= input(16);
output(1, 108) <= input(17);
output(1, 109) <= input(18);
output(1, 110) <= input(19);
output(1, 111) <= input(20);
output(1, 112) <= input(6);
output(1, 113) <= input(7);
output(1, 114) <= input(8);
output(1, 115) <= input(9);
output(1, 116) <= input(10);
output(1, 117) <= input(11);
output(1, 118) <= input(12);
output(1, 119) <= input(13);
output(1, 120) <= input(14);
output(1, 121) <= input(15);
output(1, 122) <= input(16);
output(1, 123) <= input(17);
output(1, 124) <= input(18);
output(1, 125) <= input(19);
output(1, 126) <= input(20);
output(1, 127) <= input(21);
output(1, 128) <= input(7);
output(1, 129) <= input(8);
output(1, 130) <= input(9);
output(1, 131) <= input(10);
output(1, 132) <= input(11);
output(1, 133) <= input(12);
output(1, 134) <= input(13);
output(1, 135) <= input(14);
output(1, 136) <= input(15);
output(1, 137) <= input(16);
output(1, 138) <= input(17);
output(1, 139) <= input(18);
output(1, 140) <= input(19);
output(1, 141) <= input(20);
output(1, 142) <= input(21);
output(1, 143) <= input(22);
output(1, 144) <= input(8);
output(1, 145) <= input(9);
output(1, 146) <= input(10);
output(1, 147) <= input(11);
output(1, 148) <= input(12);
output(1, 149) <= input(13);
output(1, 150) <= input(14);
output(1, 151) <= input(15);
output(1, 152) <= input(16);
output(1, 153) <= input(17);
output(1, 154) <= input(18);
output(1, 155) <= input(19);
output(1, 156) <= input(20);
output(1, 157) <= input(21);
output(1, 158) <= input(22);
output(1, 159) <= input(23);
output(1, 160) <= input(40);
output(1, 161) <= input(41);
output(1, 162) <= input(42);
output(1, 163) <= input(43);
output(1, 164) <= input(44);
output(1, 165) <= input(45);
output(1, 166) <= input(46);
output(1, 167) <= input(47);
output(1, 168) <= input(48);
output(1, 169) <= input(49);
output(1, 170) <= input(50);
output(1, 171) <= input(51);
output(1, 172) <= input(52);
output(1, 173) <= input(53);
output(1, 174) <= input(54);
output(1, 175) <= input(55);
output(1, 176) <= input(41);
output(1, 177) <= input(42);
output(1, 178) <= input(43);
output(1, 179) <= input(44);
output(1, 180) <= input(45);
output(1, 181) <= input(46);
output(1, 182) <= input(47);
output(1, 183) <= input(48);
output(1, 184) <= input(49);
output(1, 185) <= input(50);
output(1, 186) <= input(51);
output(1, 187) <= input(52);
output(1, 188) <= input(53);
output(1, 189) <= input(54);
output(1, 190) <= input(55);
output(1, 191) <= input(56);
output(1, 192) <= input(42);
output(1, 193) <= input(43);
output(1, 194) <= input(44);
output(1, 195) <= input(45);
output(1, 196) <= input(46);
output(1, 197) <= input(47);
output(1, 198) <= input(48);
output(1, 199) <= input(49);
output(1, 200) <= input(50);
output(1, 201) <= input(51);
output(1, 202) <= input(52);
output(1, 203) <= input(53);
output(1, 204) <= input(54);
output(1, 205) <= input(55);
output(1, 206) <= input(56);
output(1, 207) <= input(57);
output(1, 208) <= input(43);
output(1, 209) <= input(44);
output(1, 210) <= input(45);
output(1, 211) <= input(46);
output(1, 212) <= input(47);
output(1, 213) <= input(48);
output(1, 214) <= input(49);
output(1, 215) <= input(50);
output(1, 216) <= input(51);
output(1, 217) <= input(52);
output(1, 218) <= input(53);
output(1, 219) <= input(54);
output(1, 220) <= input(55);
output(1, 221) <= input(56);
output(1, 222) <= input(57);
output(1, 223) <= input(58);
output(1, 224) <= input(44);
output(1, 225) <= input(45);
output(1, 226) <= input(46);
output(1, 227) <= input(47);
output(1, 228) <= input(48);
output(1, 229) <= input(49);
output(1, 230) <= input(50);
output(1, 231) <= input(51);
output(1, 232) <= input(52);
output(1, 233) <= input(53);
output(1, 234) <= input(54);
output(1, 235) <= input(55);
output(1, 236) <= input(56);
output(1, 237) <= input(57);
output(1, 238) <= input(58);
output(1, 239) <= input(59);
output(1, 240) <= input(45);
output(1, 241) <= input(46);
output(1, 242) <= input(47);
output(1, 243) <= input(48);
output(1, 244) <= input(49);
output(1, 245) <= input(50);
output(1, 246) <= input(51);
output(1, 247) <= input(52);
output(1, 248) <= input(53);
output(1, 249) <= input(54);
output(1, 250) <= input(55);
output(1, 251) <= input(56);
output(1, 252) <= input(57);
output(1, 253) <= input(58);
output(1, 254) <= input(59);
output(1, 255) <= input(60);
output(2, 0) <= input(31);
output(2, 1) <= input(32);
output(2, 2) <= input(33);
output(2, 3) <= input(34);
output(2, 4) <= input(35);
output(2, 5) <= input(36);
output(2, 6) <= input(37);
output(2, 7) <= input(38);
output(2, 8) <= input(39);
output(2, 9) <= input(40);
output(2, 10) <= input(41);
output(2, 11) <= input(42);
output(2, 12) <= input(43);
output(2, 13) <= input(44);
output(2, 14) <= input(45);
output(2, 15) <= input(46);
output(2, 16) <= input(32);
output(2, 17) <= input(33);
output(2, 18) <= input(34);
output(2, 19) <= input(35);
output(2, 20) <= input(36);
output(2, 21) <= input(37);
output(2, 22) <= input(38);
output(2, 23) <= input(39);
output(2, 24) <= input(40);
output(2, 25) <= input(41);
output(2, 26) <= input(42);
output(2, 27) <= input(43);
output(2, 28) <= input(44);
output(2, 29) <= input(45);
output(2, 30) <= input(46);
output(2, 31) <= input(47);
output(2, 32) <= input(1);
output(2, 33) <= input(2);
output(2, 34) <= input(3);
output(2, 35) <= input(4);
output(2, 36) <= input(5);
output(2, 37) <= input(6);
output(2, 38) <= input(7);
output(2, 39) <= input(8);
output(2, 40) <= input(9);
output(2, 41) <= input(10);
output(2, 42) <= input(11);
output(2, 43) <= input(12);
output(2, 44) <= input(13);
output(2, 45) <= input(14);
output(2, 46) <= input(15);
output(2, 47) <= input(16);
output(2, 48) <= input(2);
output(2, 49) <= input(3);
output(2, 50) <= input(4);
output(2, 51) <= input(5);
output(2, 52) <= input(6);
output(2, 53) <= input(7);
output(2, 54) <= input(8);
output(2, 55) <= input(9);
output(2, 56) <= input(10);
output(2, 57) <= input(11);
output(2, 58) <= input(12);
output(2, 59) <= input(13);
output(2, 60) <= input(14);
output(2, 61) <= input(15);
output(2, 62) <= input(16);
output(2, 63) <= input(17);
output(2, 64) <= input(3);
output(2, 65) <= input(4);
output(2, 66) <= input(5);
output(2, 67) <= input(6);
output(2, 68) <= input(7);
output(2, 69) <= input(8);
output(2, 70) <= input(9);
output(2, 71) <= input(10);
output(2, 72) <= input(11);
output(2, 73) <= input(12);
output(2, 74) <= input(13);
output(2, 75) <= input(14);
output(2, 76) <= input(15);
output(2, 77) <= input(16);
output(2, 78) <= input(17);
output(2, 79) <= input(18);
output(2, 80) <= input(35);
output(2, 81) <= input(36);
output(2, 82) <= input(37);
output(2, 83) <= input(38);
output(2, 84) <= input(39);
output(2, 85) <= input(40);
output(2, 86) <= input(41);
output(2, 87) <= input(42);
output(2, 88) <= input(43);
output(2, 89) <= input(44);
output(2, 90) <= input(45);
output(2, 91) <= input(46);
output(2, 92) <= input(47);
output(2, 93) <= input(48);
output(2, 94) <= input(49);
output(2, 95) <= input(50);
output(2, 96) <= input(36);
output(2, 97) <= input(37);
output(2, 98) <= input(38);
output(2, 99) <= input(39);
output(2, 100) <= input(40);
output(2, 101) <= input(41);
output(2, 102) <= input(42);
output(2, 103) <= input(43);
output(2, 104) <= input(44);
output(2, 105) <= input(45);
output(2, 106) <= input(46);
output(2, 107) <= input(47);
output(2, 108) <= input(48);
output(2, 109) <= input(49);
output(2, 110) <= input(50);
output(2, 111) <= input(51);
output(2, 112) <= input(37);
output(2, 113) <= input(38);
output(2, 114) <= input(39);
output(2, 115) <= input(40);
output(2, 116) <= input(41);
output(2, 117) <= input(42);
output(2, 118) <= input(43);
output(2, 119) <= input(44);
output(2, 120) <= input(45);
output(2, 121) <= input(46);
output(2, 122) <= input(47);
output(2, 123) <= input(48);
output(2, 124) <= input(49);
output(2, 125) <= input(50);
output(2, 126) <= input(51);
output(2, 127) <= input(52);
output(2, 128) <= input(6);
output(2, 129) <= input(7);
output(2, 130) <= input(8);
output(2, 131) <= input(9);
output(2, 132) <= input(10);
output(2, 133) <= input(11);
output(2, 134) <= input(12);
output(2, 135) <= input(13);
output(2, 136) <= input(14);
output(2, 137) <= input(15);
output(2, 138) <= input(16);
output(2, 139) <= input(17);
output(2, 140) <= input(18);
output(2, 141) <= input(19);
output(2, 142) <= input(20);
output(2, 143) <= input(21);
output(2, 144) <= input(7);
output(2, 145) <= input(8);
output(2, 146) <= input(9);
output(2, 147) <= input(10);
output(2, 148) <= input(11);
output(2, 149) <= input(12);
output(2, 150) <= input(13);
output(2, 151) <= input(14);
output(2, 152) <= input(15);
output(2, 153) <= input(16);
output(2, 154) <= input(17);
output(2, 155) <= input(18);
output(2, 156) <= input(19);
output(2, 157) <= input(20);
output(2, 158) <= input(21);
output(2, 159) <= input(22);
output(2, 160) <= input(39);
output(2, 161) <= input(40);
output(2, 162) <= input(41);
output(2, 163) <= input(42);
output(2, 164) <= input(43);
output(2, 165) <= input(44);
output(2, 166) <= input(45);
output(2, 167) <= input(46);
output(2, 168) <= input(47);
output(2, 169) <= input(48);
output(2, 170) <= input(49);
output(2, 171) <= input(50);
output(2, 172) <= input(51);
output(2, 173) <= input(52);
output(2, 174) <= input(53);
output(2, 175) <= input(54);
output(2, 176) <= input(40);
output(2, 177) <= input(41);
output(2, 178) <= input(42);
output(2, 179) <= input(43);
output(2, 180) <= input(44);
output(2, 181) <= input(45);
output(2, 182) <= input(46);
output(2, 183) <= input(47);
output(2, 184) <= input(48);
output(2, 185) <= input(49);
output(2, 186) <= input(50);
output(2, 187) <= input(51);
output(2, 188) <= input(52);
output(2, 189) <= input(53);
output(2, 190) <= input(54);
output(2, 191) <= input(55);
output(2, 192) <= input(41);
output(2, 193) <= input(42);
output(2, 194) <= input(43);
output(2, 195) <= input(44);
output(2, 196) <= input(45);
output(2, 197) <= input(46);
output(2, 198) <= input(47);
output(2, 199) <= input(48);
output(2, 200) <= input(49);
output(2, 201) <= input(50);
output(2, 202) <= input(51);
output(2, 203) <= input(52);
output(2, 204) <= input(53);
output(2, 205) <= input(54);
output(2, 206) <= input(55);
output(2, 207) <= input(56);
output(2, 208) <= input(10);
output(2, 209) <= input(11);
output(2, 210) <= input(12);
output(2, 211) <= input(13);
output(2, 212) <= input(14);
output(2, 213) <= input(15);
output(2, 214) <= input(16);
output(2, 215) <= input(17);
output(2, 216) <= input(18);
output(2, 217) <= input(19);
output(2, 218) <= input(20);
output(2, 219) <= input(21);
output(2, 220) <= input(22);
output(2, 221) <= input(23);
output(2, 222) <= input(24);
output(2, 223) <= input(25);
output(2, 224) <= input(11);
output(2, 225) <= input(12);
output(2, 226) <= input(13);
output(2, 227) <= input(14);
output(2, 228) <= input(15);
output(2, 229) <= input(16);
output(2, 230) <= input(17);
output(2, 231) <= input(18);
output(2, 232) <= input(19);
output(2, 233) <= input(20);
output(2, 234) <= input(21);
output(2, 235) <= input(22);
output(2, 236) <= input(23);
output(2, 237) <= input(24);
output(2, 238) <= input(25);
output(2, 239) <= input(26);
output(2, 240) <= input(12);
output(2, 241) <= input(13);
output(2, 242) <= input(14);
output(2, 243) <= input(15);
output(2, 244) <= input(16);
output(2, 245) <= input(17);
output(2, 246) <= input(18);
output(2, 247) <= input(19);
output(2, 248) <= input(20);
output(2, 249) <= input(21);
output(2, 250) <= input(22);
output(2, 251) <= input(23);
output(2, 252) <= input(24);
output(2, 253) <= input(25);
output(2, 254) <= input(26);
output(2, 255) <= input(27);
output(3, 0) <= input(31);
output(3, 1) <= input(32);
output(3, 2) <= input(33);
output(3, 3) <= input(34);
output(3, 4) <= input(35);
output(3, 5) <= input(36);
output(3, 6) <= input(37);
output(3, 7) <= input(38);
output(3, 8) <= input(39);
output(3, 9) <= input(40);
output(3, 10) <= input(41);
output(3, 11) <= input(42);
output(3, 12) <= input(43);
output(3, 13) <= input(44);
output(3, 14) <= input(45);
output(3, 15) <= input(46);
output(3, 16) <= input(0);
output(3, 17) <= input(1);
output(3, 18) <= input(2);
output(3, 19) <= input(3);
output(3, 20) <= input(4);
output(3, 21) <= input(5);
output(3, 22) <= input(6);
output(3, 23) <= input(7);
output(3, 24) <= input(8);
output(3, 25) <= input(9);
output(3, 26) <= input(10);
output(3, 27) <= input(11);
output(3, 28) <= input(12);
output(3, 29) <= input(13);
output(3, 30) <= input(14);
output(3, 31) <= input(15);
output(3, 32) <= input(1);
output(3, 33) <= input(2);
output(3, 34) <= input(3);
output(3, 35) <= input(4);
output(3, 36) <= input(5);
output(3, 37) <= input(6);
output(3, 38) <= input(7);
output(3, 39) <= input(8);
output(3, 40) <= input(9);
output(3, 41) <= input(10);
output(3, 42) <= input(11);
output(3, 43) <= input(12);
output(3, 44) <= input(13);
output(3, 45) <= input(14);
output(3, 46) <= input(15);
output(3, 47) <= input(16);
output(3, 48) <= input(33);
output(3, 49) <= input(34);
output(3, 50) <= input(35);
output(3, 51) <= input(36);
output(3, 52) <= input(37);
output(3, 53) <= input(38);
output(3, 54) <= input(39);
output(3, 55) <= input(40);
output(3, 56) <= input(41);
output(3, 57) <= input(42);
output(3, 58) <= input(43);
output(3, 59) <= input(44);
output(3, 60) <= input(45);
output(3, 61) <= input(46);
output(3, 62) <= input(47);
output(3, 63) <= input(48);
output(3, 64) <= input(34);
output(3, 65) <= input(35);
output(3, 66) <= input(36);
output(3, 67) <= input(37);
output(3, 68) <= input(38);
output(3, 69) <= input(39);
output(3, 70) <= input(40);
output(3, 71) <= input(41);
output(3, 72) <= input(42);
output(3, 73) <= input(43);
output(3, 74) <= input(44);
output(3, 75) <= input(45);
output(3, 76) <= input(46);
output(3, 77) <= input(47);
output(3, 78) <= input(48);
output(3, 79) <= input(49);
output(3, 80) <= input(3);
output(3, 81) <= input(4);
output(3, 82) <= input(5);
output(3, 83) <= input(6);
output(3, 84) <= input(7);
output(3, 85) <= input(8);
output(3, 86) <= input(9);
output(3, 87) <= input(10);
output(3, 88) <= input(11);
output(3, 89) <= input(12);
output(3, 90) <= input(13);
output(3, 91) <= input(14);
output(3, 92) <= input(15);
output(3, 93) <= input(16);
output(3, 94) <= input(17);
output(3, 95) <= input(18);
output(3, 96) <= input(4);
output(3, 97) <= input(5);
output(3, 98) <= input(6);
output(3, 99) <= input(7);
output(3, 100) <= input(8);
output(3, 101) <= input(9);
output(3, 102) <= input(10);
output(3, 103) <= input(11);
output(3, 104) <= input(12);
output(3, 105) <= input(13);
output(3, 106) <= input(14);
output(3, 107) <= input(15);
output(3, 108) <= input(16);
output(3, 109) <= input(17);
output(3, 110) <= input(18);
output(3, 111) <= input(19);
output(3, 112) <= input(36);
output(3, 113) <= input(37);
output(3, 114) <= input(38);
output(3, 115) <= input(39);
output(3, 116) <= input(40);
output(3, 117) <= input(41);
output(3, 118) <= input(42);
output(3, 119) <= input(43);
output(3, 120) <= input(44);
output(3, 121) <= input(45);
output(3, 122) <= input(46);
output(3, 123) <= input(47);
output(3, 124) <= input(48);
output(3, 125) <= input(49);
output(3, 126) <= input(50);
output(3, 127) <= input(51);
output(3, 128) <= input(5);
output(3, 129) <= input(6);
output(3, 130) <= input(7);
output(3, 131) <= input(8);
output(3, 132) <= input(9);
output(3, 133) <= input(10);
output(3, 134) <= input(11);
output(3, 135) <= input(12);
output(3, 136) <= input(13);
output(3, 137) <= input(14);
output(3, 138) <= input(15);
output(3, 139) <= input(16);
output(3, 140) <= input(17);
output(3, 141) <= input(18);
output(3, 142) <= input(19);
output(3, 143) <= input(20);
output(3, 144) <= input(6);
output(3, 145) <= input(7);
output(3, 146) <= input(8);
output(3, 147) <= input(9);
output(3, 148) <= input(10);
output(3, 149) <= input(11);
output(3, 150) <= input(12);
output(3, 151) <= input(13);
output(3, 152) <= input(14);
output(3, 153) <= input(15);
output(3, 154) <= input(16);
output(3, 155) <= input(17);
output(3, 156) <= input(18);
output(3, 157) <= input(19);
output(3, 158) <= input(20);
output(3, 159) <= input(21);
output(3, 160) <= input(38);
output(3, 161) <= input(39);
output(3, 162) <= input(40);
output(3, 163) <= input(41);
output(3, 164) <= input(42);
output(3, 165) <= input(43);
output(3, 166) <= input(44);
output(3, 167) <= input(45);
output(3, 168) <= input(46);
output(3, 169) <= input(47);
output(3, 170) <= input(48);
output(3, 171) <= input(49);
output(3, 172) <= input(50);
output(3, 173) <= input(51);
output(3, 174) <= input(52);
output(3, 175) <= input(53);
output(3, 176) <= input(39);
output(3, 177) <= input(40);
output(3, 178) <= input(41);
output(3, 179) <= input(42);
output(3, 180) <= input(43);
output(3, 181) <= input(44);
output(3, 182) <= input(45);
output(3, 183) <= input(46);
output(3, 184) <= input(47);
output(3, 185) <= input(48);
output(3, 186) <= input(49);
output(3, 187) <= input(50);
output(3, 188) <= input(51);
output(3, 189) <= input(52);
output(3, 190) <= input(53);
output(3, 191) <= input(54);
output(3, 192) <= input(8);
output(3, 193) <= input(9);
output(3, 194) <= input(10);
output(3, 195) <= input(11);
output(3, 196) <= input(12);
output(3, 197) <= input(13);
output(3, 198) <= input(14);
output(3, 199) <= input(15);
output(3, 200) <= input(16);
output(3, 201) <= input(17);
output(3, 202) <= input(18);
output(3, 203) <= input(19);
output(3, 204) <= input(20);
output(3, 205) <= input(21);
output(3, 206) <= input(22);
output(3, 207) <= input(23);
output(3, 208) <= input(9);
output(3, 209) <= input(10);
output(3, 210) <= input(11);
output(3, 211) <= input(12);
output(3, 212) <= input(13);
output(3, 213) <= input(14);
output(3, 214) <= input(15);
output(3, 215) <= input(16);
output(3, 216) <= input(17);
output(3, 217) <= input(18);
output(3, 218) <= input(19);
output(3, 219) <= input(20);
output(3, 220) <= input(21);
output(3, 221) <= input(22);
output(3, 222) <= input(23);
output(3, 223) <= input(24);
output(3, 224) <= input(41);
output(3, 225) <= input(42);
output(3, 226) <= input(43);
output(3, 227) <= input(44);
output(3, 228) <= input(45);
output(3, 229) <= input(46);
output(3, 230) <= input(47);
output(3, 231) <= input(48);
output(3, 232) <= input(49);
output(3, 233) <= input(50);
output(3, 234) <= input(51);
output(3, 235) <= input(52);
output(3, 236) <= input(53);
output(3, 237) <= input(54);
output(3, 238) <= input(55);
output(3, 239) <= input(56);
output(3, 240) <= input(42);
output(3, 241) <= input(43);
output(3, 242) <= input(44);
output(3, 243) <= input(45);
output(3, 244) <= input(46);
output(3, 245) <= input(47);
output(3, 246) <= input(48);
output(3, 247) <= input(49);
output(3, 248) <= input(50);
output(3, 249) <= input(51);
output(3, 250) <= input(52);
output(3, 251) <= input(53);
output(3, 252) <= input(54);
output(3, 253) <= input(55);
output(3, 254) <= input(56);
output(3, 255) <= input(57);
output(4, 0) <= input(31);
output(4, 1) <= input(32);
output(4, 2) <= input(33);
output(4, 3) <= input(34);
output(4, 4) <= input(35);
output(4, 5) <= input(36);
output(4, 6) <= input(37);
output(4, 7) <= input(38);
output(4, 8) <= input(39);
output(4, 9) <= input(40);
output(4, 10) <= input(41);
output(4, 11) <= input(42);
output(4, 12) <= input(43);
output(4, 13) <= input(44);
output(4, 14) <= input(45);
output(4, 15) <= input(46);
output(4, 16) <= input(0);
output(4, 17) <= input(1);
output(4, 18) <= input(2);
output(4, 19) <= input(3);
output(4, 20) <= input(4);
output(4, 21) <= input(5);
output(4, 22) <= input(6);
output(4, 23) <= input(7);
output(4, 24) <= input(8);
output(4, 25) <= input(9);
output(4, 26) <= input(10);
output(4, 27) <= input(11);
output(4, 28) <= input(12);
output(4, 29) <= input(13);
output(4, 30) <= input(14);
output(4, 31) <= input(15);
output(4, 32) <= input(32);
output(4, 33) <= input(33);
output(4, 34) <= input(34);
output(4, 35) <= input(35);
output(4, 36) <= input(36);
output(4, 37) <= input(37);
output(4, 38) <= input(38);
output(4, 39) <= input(39);
output(4, 40) <= input(40);
output(4, 41) <= input(41);
output(4, 42) <= input(42);
output(4, 43) <= input(43);
output(4, 44) <= input(44);
output(4, 45) <= input(45);
output(4, 46) <= input(46);
output(4, 47) <= input(47);
output(4, 48) <= input(33);
output(4, 49) <= input(34);
output(4, 50) <= input(35);
output(4, 51) <= input(36);
output(4, 52) <= input(37);
output(4, 53) <= input(38);
output(4, 54) <= input(39);
output(4, 55) <= input(40);
output(4, 56) <= input(41);
output(4, 57) <= input(42);
output(4, 58) <= input(43);
output(4, 59) <= input(44);
output(4, 60) <= input(45);
output(4, 61) <= input(46);
output(4, 62) <= input(47);
output(4, 63) <= input(48);
output(4, 64) <= input(2);
output(4, 65) <= input(3);
output(4, 66) <= input(4);
output(4, 67) <= input(5);
output(4, 68) <= input(6);
output(4, 69) <= input(7);
output(4, 70) <= input(8);
output(4, 71) <= input(9);
output(4, 72) <= input(10);
output(4, 73) <= input(11);
output(4, 74) <= input(12);
output(4, 75) <= input(13);
output(4, 76) <= input(14);
output(4, 77) <= input(15);
output(4, 78) <= input(16);
output(4, 79) <= input(17);
output(4, 80) <= input(34);
output(4, 81) <= input(35);
output(4, 82) <= input(36);
output(4, 83) <= input(37);
output(4, 84) <= input(38);
output(4, 85) <= input(39);
output(4, 86) <= input(40);
output(4, 87) <= input(41);
output(4, 88) <= input(42);
output(4, 89) <= input(43);
output(4, 90) <= input(44);
output(4, 91) <= input(45);
output(4, 92) <= input(46);
output(4, 93) <= input(47);
output(4, 94) <= input(48);
output(4, 95) <= input(49);
output(4, 96) <= input(3);
output(4, 97) <= input(4);
output(4, 98) <= input(5);
output(4, 99) <= input(6);
output(4, 100) <= input(7);
output(4, 101) <= input(8);
output(4, 102) <= input(9);
output(4, 103) <= input(10);
output(4, 104) <= input(11);
output(4, 105) <= input(12);
output(4, 106) <= input(13);
output(4, 107) <= input(14);
output(4, 108) <= input(15);
output(4, 109) <= input(16);
output(4, 110) <= input(17);
output(4, 111) <= input(18);
output(4, 112) <= input(4);
output(4, 113) <= input(5);
output(4, 114) <= input(6);
output(4, 115) <= input(7);
output(4, 116) <= input(8);
output(4, 117) <= input(9);
output(4, 118) <= input(10);
output(4, 119) <= input(11);
output(4, 120) <= input(12);
output(4, 121) <= input(13);
output(4, 122) <= input(14);
output(4, 123) <= input(15);
output(4, 124) <= input(16);
output(4, 125) <= input(17);
output(4, 126) <= input(18);
output(4, 127) <= input(19);
output(4, 128) <= input(36);
output(4, 129) <= input(37);
output(4, 130) <= input(38);
output(4, 131) <= input(39);
output(4, 132) <= input(40);
output(4, 133) <= input(41);
output(4, 134) <= input(42);
output(4, 135) <= input(43);
output(4, 136) <= input(44);
output(4, 137) <= input(45);
output(4, 138) <= input(46);
output(4, 139) <= input(47);
output(4, 140) <= input(48);
output(4, 141) <= input(49);
output(4, 142) <= input(50);
output(4, 143) <= input(51);
output(4, 144) <= input(5);
output(4, 145) <= input(6);
output(4, 146) <= input(7);
output(4, 147) <= input(8);
output(4, 148) <= input(9);
output(4, 149) <= input(10);
output(4, 150) <= input(11);
output(4, 151) <= input(12);
output(4, 152) <= input(13);
output(4, 153) <= input(14);
output(4, 154) <= input(15);
output(4, 155) <= input(16);
output(4, 156) <= input(17);
output(4, 157) <= input(18);
output(4, 158) <= input(19);
output(4, 159) <= input(20);
output(4, 160) <= input(37);
output(4, 161) <= input(38);
output(4, 162) <= input(39);
output(4, 163) <= input(40);
output(4, 164) <= input(41);
output(4, 165) <= input(42);
output(4, 166) <= input(43);
output(4, 167) <= input(44);
output(4, 168) <= input(45);
output(4, 169) <= input(46);
output(4, 170) <= input(47);
output(4, 171) <= input(48);
output(4, 172) <= input(49);
output(4, 173) <= input(50);
output(4, 174) <= input(51);
output(4, 175) <= input(52);
output(4, 176) <= input(38);
output(4, 177) <= input(39);
output(4, 178) <= input(40);
output(4, 179) <= input(41);
output(4, 180) <= input(42);
output(4, 181) <= input(43);
output(4, 182) <= input(44);
output(4, 183) <= input(45);
output(4, 184) <= input(46);
output(4, 185) <= input(47);
output(4, 186) <= input(48);
output(4, 187) <= input(49);
output(4, 188) <= input(50);
output(4, 189) <= input(51);
output(4, 190) <= input(52);
output(4, 191) <= input(53);
output(4, 192) <= input(7);
output(4, 193) <= input(8);
output(4, 194) <= input(9);
output(4, 195) <= input(10);
output(4, 196) <= input(11);
output(4, 197) <= input(12);
output(4, 198) <= input(13);
output(4, 199) <= input(14);
output(4, 200) <= input(15);
output(4, 201) <= input(16);
output(4, 202) <= input(17);
output(4, 203) <= input(18);
output(4, 204) <= input(19);
output(4, 205) <= input(20);
output(4, 206) <= input(21);
output(4, 207) <= input(22);
output(4, 208) <= input(39);
output(4, 209) <= input(40);
output(4, 210) <= input(41);
output(4, 211) <= input(42);
output(4, 212) <= input(43);
output(4, 213) <= input(44);
output(4, 214) <= input(45);
output(4, 215) <= input(46);
output(4, 216) <= input(47);
output(4, 217) <= input(48);
output(4, 218) <= input(49);
output(4, 219) <= input(50);
output(4, 220) <= input(51);
output(4, 221) <= input(52);
output(4, 222) <= input(53);
output(4, 223) <= input(54);
output(4, 224) <= input(8);
output(4, 225) <= input(9);
output(4, 226) <= input(10);
output(4, 227) <= input(11);
output(4, 228) <= input(12);
output(4, 229) <= input(13);
output(4, 230) <= input(14);
output(4, 231) <= input(15);
output(4, 232) <= input(16);
output(4, 233) <= input(17);
output(4, 234) <= input(18);
output(4, 235) <= input(19);
output(4, 236) <= input(20);
output(4, 237) <= input(21);
output(4, 238) <= input(22);
output(4, 239) <= input(23);
output(4, 240) <= input(9);
output(4, 241) <= input(10);
output(4, 242) <= input(11);
output(4, 243) <= input(12);
output(4, 244) <= input(13);
output(4, 245) <= input(14);
output(4, 246) <= input(15);
output(4, 247) <= input(16);
output(4, 248) <= input(17);
output(4, 249) <= input(18);
output(4, 250) <= input(19);
output(4, 251) <= input(20);
output(4, 252) <= input(21);
output(4, 253) <= input(22);
output(4, 254) <= input(23);
output(4, 255) <= input(24);
output(5, 0) <= input(31);
output(5, 1) <= input(32);
output(5, 2) <= input(33);
output(5, 3) <= input(34);
output(5, 4) <= input(35);
output(5, 5) <= input(36);
output(5, 6) <= input(37);
output(5, 7) <= input(38);
output(5, 8) <= input(39);
output(5, 9) <= input(40);
output(5, 10) <= input(41);
output(5, 11) <= input(42);
output(5, 12) <= input(43);
output(5, 13) <= input(44);
output(5, 14) <= input(45);
output(5, 15) <= input(46);
output(5, 16) <= input(0);
output(5, 17) <= input(1);
output(5, 18) <= input(2);
output(5, 19) <= input(3);
output(5, 20) <= input(4);
output(5, 21) <= input(5);
output(5, 22) <= input(6);
output(5, 23) <= input(7);
output(5, 24) <= input(8);
output(5, 25) <= input(9);
output(5, 26) <= input(10);
output(5, 27) <= input(11);
output(5, 28) <= input(12);
output(5, 29) <= input(13);
output(5, 30) <= input(14);
output(5, 31) <= input(15);
output(5, 32) <= input(32);
output(5, 33) <= input(33);
output(5, 34) <= input(34);
output(5, 35) <= input(35);
output(5, 36) <= input(36);
output(5, 37) <= input(37);
output(5, 38) <= input(38);
output(5, 39) <= input(39);
output(5, 40) <= input(40);
output(5, 41) <= input(41);
output(5, 42) <= input(42);
output(5, 43) <= input(43);
output(5, 44) <= input(44);
output(5, 45) <= input(45);
output(5, 46) <= input(46);
output(5, 47) <= input(47);
output(5, 48) <= input(1);
output(5, 49) <= input(2);
output(5, 50) <= input(3);
output(5, 51) <= input(4);
output(5, 52) <= input(5);
output(5, 53) <= input(6);
output(5, 54) <= input(7);
output(5, 55) <= input(8);
output(5, 56) <= input(9);
output(5, 57) <= input(10);
output(5, 58) <= input(11);
output(5, 59) <= input(12);
output(5, 60) <= input(13);
output(5, 61) <= input(14);
output(5, 62) <= input(15);
output(5, 63) <= input(16);
output(5, 64) <= input(33);
output(5, 65) <= input(34);
output(5, 66) <= input(35);
output(5, 67) <= input(36);
output(5, 68) <= input(37);
output(5, 69) <= input(38);
output(5, 70) <= input(39);
output(5, 71) <= input(40);
output(5, 72) <= input(41);
output(5, 73) <= input(42);
output(5, 74) <= input(43);
output(5, 75) <= input(44);
output(5, 76) <= input(45);
output(5, 77) <= input(46);
output(5, 78) <= input(47);
output(5, 79) <= input(48);
output(5, 80) <= input(2);
output(5, 81) <= input(3);
output(5, 82) <= input(4);
output(5, 83) <= input(5);
output(5, 84) <= input(6);
output(5, 85) <= input(7);
output(5, 86) <= input(8);
output(5, 87) <= input(9);
output(5, 88) <= input(10);
output(5, 89) <= input(11);
output(5, 90) <= input(12);
output(5, 91) <= input(13);
output(5, 92) <= input(14);
output(5, 93) <= input(15);
output(5, 94) <= input(16);
output(5, 95) <= input(17);
output(5, 96) <= input(34);
output(5, 97) <= input(35);
output(5, 98) <= input(36);
output(5, 99) <= input(37);
output(5, 100) <= input(38);
output(5, 101) <= input(39);
output(5, 102) <= input(40);
output(5, 103) <= input(41);
output(5, 104) <= input(42);
output(5, 105) <= input(43);
output(5, 106) <= input(44);
output(5, 107) <= input(45);
output(5, 108) <= input(46);
output(5, 109) <= input(47);
output(5, 110) <= input(48);
output(5, 111) <= input(49);
output(5, 112) <= input(35);
output(5, 113) <= input(36);
output(5, 114) <= input(37);
output(5, 115) <= input(38);
output(5, 116) <= input(39);
output(5, 117) <= input(40);
output(5, 118) <= input(41);
output(5, 119) <= input(42);
output(5, 120) <= input(43);
output(5, 121) <= input(44);
output(5, 122) <= input(45);
output(5, 123) <= input(46);
output(5, 124) <= input(47);
output(5, 125) <= input(48);
output(5, 126) <= input(49);
output(5, 127) <= input(50);
output(5, 128) <= input(4);
output(5, 129) <= input(5);
output(5, 130) <= input(6);
output(5, 131) <= input(7);
output(5, 132) <= input(8);
output(5, 133) <= input(9);
output(5, 134) <= input(10);
output(5, 135) <= input(11);
output(5, 136) <= input(12);
output(5, 137) <= input(13);
output(5, 138) <= input(14);
output(5, 139) <= input(15);
output(5, 140) <= input(16);
output(5, 141) <= input(17);
output(5, 142) <= input(18);
output(5, 143) <= input(19);
output(5, 144) <= input(36);
output(5, 145) <= input(37);
output(5, 146) <= input(38);
output(5, 147) <= input(39);
output(5, 148) <= input(40);
output(5, 149) <= input(41);
output(5, 150) <= input(42);
output(5, 151) <= input(43);
output(5, 152) <= input(44);
output(5, 153) <= input(45);
output(5, 154) <= input(46);
output(5, 155) <= input(47);
output(5, 156) <= input(48);
output(5, 157) <= input(49);
output(5, 158) <= input(50);
output(5, 159) <= input(51);
output(5, 160) <= input(5);
output(5, 161) <= input(6);
output(5, 162) <= input(7);
output(5, 163) <= input(8);
output(5, 164) <= input(9);
output(5, 165) <= input(10);
output(5, 166) <= input(11);
output(5, 167) <= input(12);
output(5, 168) <= input(13);
output(5, 169) <= input(14);
output(5, 170) <= input(15);
output(5, 171) <= input(16);
output(5, 172) <= input(17);
output(5, 173) <= input(18);
output(5, 174) <= input(19);
output(5, 175) <= input(20);
output(5, 176) <= input(37);
output(5, 177) <= input(38);
output(5, 178) <= input(39);
output(5, 179) <= input(40);
output(5, 180) <= input(41);
output(5, 181) <= input(42);
output(5, 182) <= input(43);
output(5, 183) <= input(44);
output(5, 184) <= input(45);
output(5, 185) <= input(46);
output(5, 186) <= input(47);
output(5, 187) <= input(48);
output(5, 188) <= input(49);
output(5, 189) <= input(50);
output(5, 190) <= input(51);
output(5, 191) <= input(52);
output(5, 192) <= input(6);
output(5, 193) <= input(7);
output(5, 194) <= input(8);
output(5, 195) <= input(9);
output(5, 196) <= input(10);
output(5, 197) <= input(11);
output(5, 198) <= input(12);
output(5, 199) <= input(13);
output(5, 200) <= input(14);
output(5, 201) <= input(15);
output(5, 202) <= input(16);
output(5, 203) <= input(17);
output(5, 204) <= input(18);
output(5, 205) <= input(19);
output(5, 206) <= input(20);
output(5, 207) <= input(21);
output(5, 208) <= input(38);
output(5, 209) <= input(39);
output(5, 210) <= input(40);
output(5, 211) <= input(41);
output(5, 212) <= input(42);
output(5, 213) <= input(43);
output(5, 214) <= input(44);
output(5, 215) <= input(45);
output(5, 216) <= input(46);
output(5, 217) <= input(47);
output(5, 218) <= input(48);
output(5, 219) <= input(49);
output(5, 220) <= input(50);
output(5, 221) <= input(51);
output(5, 222) <= input(52);
output(5, 223) <= input(53);
output(5, 224) <= input(7);
output(5, 225) <= input(8);
output(5, 226) <= input(9);
output(5, 227) <= input(10);
output(5, 228) <= input(11);
output(5, 229) <= input(12);
output(5, 230) <= input(13);
output(5, 231) <= input(14);
output(5, 232) <= input(15);
output(5, 233) <= input(16);
output(5, 234) <= input(17);
output(5, 235) <= input(18);
output(5, 236) <= input(19);
output(5, 237) <= input(20);
output(5, 238) <= input(21);
output(5, 239) <= input(22);
output(5, 240) <= input(8);
output(5, 241) <= input(9);
output(5, 242) <= input(10);
output(5, 243) <= input(11);
output(5, 244) <= input(12);
output(5, 245) <= input(13);
output(5, 246) <= input(14);
output(5, 247) <= input(15);
output(5, 248) <= input(16);
output(5, 249) <= input(17);
output(5, 250) <= input(18);
output(5, 251) <= input(19);
output(5, 252) <= input(20);
output(5, 253) <= input(21);
output(5, 254) <= input(22);
output(5, 255) <= input(23);
when "0001" =>
output(0, 0) <= input(0);
output(0, 1) <= input(1);
output(0, 2) <= input(2);
output(0, 3) <= input(3);
output(0, 4) <= input(4);
output(0, 5) <= input(5);
output(0, 6) <= input(6);
output(0, 7) <= input(7);
output(0, 8) <= input(8);
output(0, 9) <= input(9);
output(0, 10) <= input(10);
output(0, 11) <= input(11);
output(0, 12) <= input(12);
output(0, 13) <= input(13);
output(0, 14) <= input(14);
output(0, 15) <= input(15);
output(0, 16) <= input(16);
output(0, 17) <= input(17);
output(0, 18) <= input(18);
output(0, 19) <= input(19);
output(0, 20) <= input(20);
output(0, 21) <= input(21);
output(0, 22) <= input(22);
output(0, 23) <= input(23);
output(0, 24) <= input(24);
output(0, 25) <= input(25);
output(0, 26) <= input(26);
output(0, 27) <= input(27);
output(0, 28) <= input(28);
output(0, 29) <= input(29);
output(0, 30) <= input(30);
output(0, 31) <= input(31);
output(0, 32) <= input(1);
output(0, 33) <= input(2);
output(0, 34) <= input(3);
output(0, 35) <= input(4);
output(0, 36) <= input(5);
output(0, 37) <= input(6);
output(0, 38) <= input(7);
output(0, 39) <= input(8);
output(0, 40) <= input(9);
output(0, 41) <= input(10);
output(0, 42) <= input(11);
output(0, 43) <= input(12);
output(0, 44) <= input(13);
output(0, 45) <= input(14);
output(0, 46) <= input(15);
output(0, 47) <= input(32);
output(0, 48) <= input(17);
output(0, 49) <= input(18);
output(0, 50) <= input(19);
output(0, 51) <= input(20);
output(0, 52) <= input(21);
output(0, 53) <= input(22);
output(0, 54) <= input(23);
output(0, 55) <= input(24);
output(0, 56) <= input(25);
output(0, 57) <= input(26);
output(0, 58) <= input(27);
output(0, 59) <= input(28);
output(0, 60) <= input(29);
output(0, 61) <= input(30);
output(0, 62) <= input(31);
output(0, 63) <= input(33);
output(0, 64) <= input(2);
output(0, 65) <= input(3);
output(0, 66) <= input(4);
output(0, 67) <= input(5);
output(0, 68) <= input(6);
output(0, 69) <= input(7);
output(0, 70) <= input(8);
output(0, 71) <= input(9);
output(0, 72) <= input(10);
output(0, 73) <= input(11);
output(0, 74) <= input(12);
output(0, 75) <= input(13);
output(0, 76) <= input(14);
output(0, 77) <= input(15);
output(0, 78) <= input(32);
output(0, 79) <= input(34);
output(0, 80) <= input(18);
output(0, 81) <= input(19);
output(0, 82) <= input(20);
output(0, 83) <= input(21);
output(0, 84) <= input(22);
output(0, 85) <= input(23);
output(0, 86) <= input(24);
output(0, 87) <= input(25);
output(0, 88) <= input(26);
output(0, 89) <= input(27);
output(0, 90) <= input(28);
output(0, 91) <= input(29);
output(0, 92) <= input(30);
output(0, 93) <= input(31);
output(0, 94) <= input(33);
output(0, 95) <= input(35);
output(0, 96) <= input(3);
output(0, 97) <= input(4);
output(0, 98) <= input(5);
output(0, 99) <= input(6);
output(0, 100) <= input(7);
output(0, 101) <= input(8);
output(0, 102) <= input(9);
output(0, 103) <= input(10);
output(0, 104) <= input(11);
output(0, 105) <= input(12);
output(0, 106) <= input(13);
output(0, 107) <= input(14);
output(0, 108) <= input(15);
output(0, 109) <= input(32);
output(0, 110) <= input(34);
output(0, 111) <= input(36);
output(0, 112) <= input(19);
output(0, 113) <= input(20);
output(0, 114) <= input(21);
output(0, 115) <= input(22);
output(0, 116) <= input(23);
output(0, 117) <= input(24);
output(0, 118) <= input(25);
output(0, 119) <= input(26);
output(0, 120) <= input(27);
output(0, 121) <= input(28);
output(0, 122) <= input(29);
output(0, 123) <= input(30);
output(0, 124) <= input(31);
output(0, 125) <= input(33);
output(0, 126) <= input(35);
output(0, 127) <= input(37);
output(0, 128) <= input(4);
output(0, 129) <= input(5);
output(0, 130) <= input(6);
output(0, 131) <= input(7);
output(0, 132) <= input(8);
output(0, 133) <= input(9);
output(0, 134) <= input(10);
output(0, 135) <= input(11);
output(0, 136) <= input(12);
output(0, 137) <= input(13);
output(0, 138) <= input(14);
output(0, 139) <= input(15);
output(0, 140) <= input(32);
output(0, 141) <= input(34);
output(0, 142) <= input(36);
output(0, 143) <= input(38);
output(0, 144) <= input(20);
output(0, 145) <= input(21);
output(0, 146) <= input(22);
output(0, 147) <= input(23);
output(0, 148) <= input(24);
output(0, 149) <= input(25);
output(0, 150) <= input(26);
output(0, 151) <= input(27);
output(0, 152) <= input(28);
output(0, 153) <= input(29);
output(0, 154) <= input(30);
output(0, 155) <= input(31);
output(0, 156) <= input(33);
output(0, 157) <= input(35);
output(0, 158) <= input(37);
output(0, 159) <= input(39);
output(0, 160) <= input(5);
output(0, 161) <= input(6);
output(0, 162) <= input(7);
output(0, 163) <= input(8);
output(0, 164) <= input(9);
output(0, 165) <= input(10);
output(0, 166) <= input(11);
output(0, 167) <= input(12);
output(0, 168) <= input(13);
output(0, 169) <= input(14);
output(0, 170) <= input(15);
output(0, 171) <= input(32);
output(0, 172) <= input(34);
output(0, 173) <= input(36);
output(0, 174) <= input(38);
output(0, 175) <= input(40);
output(0, 176) <= input(21);
output(0, 177) <= input(22);
output(0, 178) <= input(23);
output(0, 179) <= input(24);
output(0, 180) <= input(25);
output(0, 181) <= input(26);
output(0, 182) <= input(27);
output(0, 183) <= input(28);
output(0, 184) <= input(29);
output(0, 185) <= input(30);
output(0, 186) <= input(31);
output(0, 187) <= input(33);
output(0, 188) <= input(35);
output(0, 189) <= input(37);
output(0, 190) <= input(39);
output(0, 191) <= input(41);
output(0, 192) <= input(6);
output(0, 193) <= input(7);
output(0, 194) <= input(8);
output(0, 195) <= input(9);
output(0, 196) <= input(10);
output(0, 197) <= input(11);
output(0, 198) <= input(12);
output(0, 199) <= input(13);
output(0, 200) <= input(14);
output(0, 201) <= input(15);
output(0, 202) <= input(32);
output(0, 203) <= input(34);
output(0, 204) <= input(36);
output(0, 205) <= input(38);
output(0, 206) <= input(40);
output(0, 207) <= input(42);
output(0, 208) <= input(22);
output(0, 209) <= input(23);
output(0, 210) <= input(24);
output(0, 211) <= input(25);
output(0, 212) <= input(26);
output(0, 213) <= input(27);
output(0, 214) <= input(28);
output(0, 215) <= input(29);
output(0, 216) <= input(30);
output(0, 217) <= input(31);
output(0, 218) <= input(33);
output(0, 219) <= input(35);
output(0, 220) <= input(37);
output(0, 221) <= input(39);
output(0, 222) <= input(41);
output(0, 223) <= input(43);
output(0, 224) <= input(7);
output(0, 225) <= input(8);
output(0, 226) <= input(9);
output(0, 227) <= input(10);
output(0, 228) <= input(11);
output(0, 229) <= input(12);
output(0, 230) <= input(13);
output(0, 231) <= input(14);
output(0, 232) <= input(15);
output(0, 233) <= input(32);
output(0, 234) <= input(34);
output(0, 235) <= input(36);
output(0, 236) <= input(38);
output(0, 237) <= input(40);
output(0, 238) <= input(42);
output(0, 239) <= input(44);
output(0, 240) <= input(23);
output(0, 241) <= input(24);
output(0, 242) <= input(25);
output(0, 243) <= input(26);
output(0, 244) <= input(27);
output(0, 245) <= input(28);
output(0, 246) <= input(29);
output(0, 247) <= input(30);
output(0, 248) <= input(31);
output(0, 249) <= input(33);
output(0, 250) <= input(35);
output(0, 251) <= input(37);
output(0, 252) <= input(39);
output(0, 253) <= input(41);
output(0, 254) <= input(43);
output(0, 255) <= input(45);
output(1, 0) <= input(46);
output(1, 1) <= input(16);
output(1, 2) <= input(17);
output(1, 3) <= input(18);
output(1, 4) <= input(19);
output(1, 5) <= input(20);
output(1, 6) <= input(21);
output(1, 7) <= input(22);
output(1, 8) <= input(23);
output(1, 9) <= input(24);
output(1, 10) <= input(25);
output(1, 11) <= input(26);
output(1, 12) <= input(27);
output(1, 13) <= input(28);
output(1, 14) <= input(29);
output(1, 15) <= input(30);
output(1, 16) <= input(0);
output(1, 17) <= input(1);
output(1, 18) <= input(2);
output(1, 19) <= input(3);
output(1, 20) <= input(4);
output(1, 21) <= input(5);
output(1, 22) <= input(6);
output(1, 23) <= input(7);
output(1, 24) <= input(8);
output(1, 25) <= input(9);
output(1, 26) <= input(10);
output(1, 27) <= input(11);
output(1, 28) <= input(12);
output(1, 29) <= input(13);
output(1, 30) <= input(14);
output(1, 31) <= input(15);
output(1, 32) <= input(16);
output(1, 33) <= input(17);
output(1, 34) <= input(18);
output(1, 35) <= input(19);
output(1, 36) <= input(20);
output(1, 37) <= input(21);
output(1, 38) <= input(22);
output(1, 39) <= input(23);
output(1, 40) <= input(24);
output(1, 41) <= input(25);
output(1, 42) <= input(26);
output(1, 43) <= input(27);
output(1, 44) <= input(28);
output(1, 45) <= input(29);
output(1, 46) <= input(30);
output(1, 47) <= input(31);
output(1, 48) <= input(1);
output(1, 49) <= input(2);
output(1, 50) <= input(3);
output(1, 51) <= input(4);
output(1, 52) <= input(5);
output(1, 53) <= input(6);
output(1, 54) <= input(7);
output(1, 55) <= input(8);
output(1, 56) <= input(9);
output(1, 57) <= input(10);
output(1, 58) <= input(11);
output(1, 59) <= input(12);
output(1, 60) <= input(13);
output(1, 61) <= input(14);
output(1, 62) <= input(15);
output(1, 63) <= input(32);
output(1, 64) <= input(17);
output(1, 65) <= input(18);
output(1, 66) <= input(19);
output(1, 67) <= input(20);
output(1, 68) <= input(21);
output(1, 69) <= input(22);
output(1, 70) <= input(23);
output(1, 71) <= input(24);
output(1, 72) <= input(25);
output(1, 73) <= input(26);
output(1, 74) <= input(27);
output(1, 75) <= input(28);
output(1, 76) <= input(29);
output(1, 77) <= input(30);
output(1, 78) <= input(31);
output(1, 79) <= input(33);
output(1, 80) <= input(2);
output(1, 81) <= input(3);
output(1, 82) <= input(4);
output(1, 83) <= input(5);
output(1, 84) <= input(6);
output(1, 85) <= input(7);
output(1, 86) <= input(8);
output(1, 87) <= input(9);
output(1, 88) <= input(10);
output(1, 89) <= input(11);
output(1, 90) <= input(12);
output(1, 91) <= input(13);
output(1, 92) <= input(14);
output(1, 93) <= input(15);
output(1, 94) <= input(32);
output(1, 95) <= input(34);
output(1, 96) <= input(18);
output(1, 97) <= input(19);
output(1, 98) <= input(20);
output(1, 99) <= input(21);
output(1, 100) <= input(22);
output(1, 101) <= input(23);
output(1, 102) <= input(24);
output(1, 103) <= input(25);
output(1, 104) <= input(26);
output(1, 105) <= input(27);
output(1, 106) <= input(28);
output(1, 107) <= input(29);
output(1, 108) <= input(30);
output(1, 109) <= input(31);
output(1, 110) <= input(33);
output(1, 111) <= input(35);
output(1, 112) <= input(3);
output(1, 113) <= input(4);
output(1, 114) <= input(5);
output(1, 115) <= input(6);
output(1, 116) <= input(7);
output(1, 117) <= input(8);
output(1, 118) <= input(9);
output(1, 119) <= input(10);
output(1, 120) <= input(11);
output(1, 121) <= input(12);
output(1, 122) <= input(13);
output(1, 123) <= input(14);
output(1, 124) <= input(15);
output(1, 125) <= input(32);
output(1, 126) <= input(34);
output(1, 127) <= input(36);
output(1, 128) <= input(3);
output(1, 129) <= input(4);
output(1, 130) <= input(5);
output(1, 131) <= input(6);
output(1, 132) <= input(7);
output(1, 133) <= input(8);
output(1, 134) <= input(9);
output(1, 135) <= input(10);
output(1, 136) <= input(11);
output(1, 137) <= input(12);
output(1, 138) <= input(13);
output(1, 139) <= input(14);
output(1, 140) <= input(15);
output(1, 141) <= input(32);
output(1, 142) <= input(34);
output(1, 143) <= input(36);
output(1, 144) <= input(19);
output(1, 145) <= input(20);
output(1, 146) <= input(21);
output(1, 147) <= input(22);
output(1, 148) <= input(23);
output(1, 149) <= input(24);
output(1, 150) <= input(25);
output(1, 151) <= input(26);
output(1, 152) <= input(27);
output(1, 153) <= input(28);
output(1, 154) <= input(29);
output(1, 155) <= input(30);
output(1, 156) <= input(31);
output(1, 157) <= input(33);
output(1, 158) <= input(35);
output(1, 159) <= input(37);
output(1, 160) <= input(4);
output(1, 161) <= input(5);
output(1, 162) <= input(6);
output(1, 163) <= input(7);
output(1, 164) <= input(8);
output(1, 165) <= input(9);
output(1, 166) <= input(10);
output(1, 167) <= input(11);
output(1, 168) <= input(12);
output(1, 169) <= input(13);
output(1, 170) <= input(14);
output(1, 171) <= input(15);
output(1, 172) <= input(32);
output(1, 173) <= input(34);
output(1, 174) <= input(36);
output(1, 175) <= input(38);
output(1, 176) <= input(20);
output(1, 177) <= input(21);
output(1, 178) <= input(22);
output(1, 179) <= input(23);
output(1, 180) <= input(24);
output(1, 181) <= input(25);
output(1, 182) <= input(26);
output(1, 183) <= input(27);
output(1, 184) <= input(28);
output(1, 185) <= input(29);
output(1, 186) <= input(30);
output(1, 187) <= input(31);
output(1, 188) <= input(33);
output(1, 189) <= input(35);
output(1, 190) <= input(37);
output(1, 191) <= input(39);
output(1, 192) <= input(5);
output(1, 193) <= input(6);
output(1, 194) <= input(7);
output(1, 195) <= input(8);
output(1, 196) <= input(9);
output(1, 197) <= input(10);
output(1, 198) <= input(11);
output(1, 199) <= input(12);
output(1, 200) <= input(13);
output(1, 201) <= input(14);
output(1, 202) <= input(15);
output(1, 203) <= input(32);
output(1, 204) <= input(34);
output(1, 205) <= input(36);
output(1, 206) <= input(38);
output(1, 207) <= input(40);
output(1, 208) <= input(21);
output(1, 209) <= input(22);
output(1, 210) <= input(23);
output(1, 211) <= input(24);
output(1, 212) <= input(25);
output(1, 213) <= input(26);
output(1, 214) <= input(27);
output(1, 215) <= input(28);
output(1, 216) <= input(29);
output(1, 217) <= input(30);
output(1, 218) <= input(31);
output(1, 219) <= input(33);
output(1, 220) <= input(35);
output(1, 221) <= input(37);
output(1, 222) <= input(39);
output(1, 223) <= input(41);
output(1, 224) <= input(6);
output(1, 225) <= input(7);
output(1, 226) <= input(8);
output(1, 227) <= input(9);
output(1, 228) <= input(10);
output(1, 229) <= input(11);
output(1, 230) <= input(12);
output(1, 231) <= input(13);
output(1, 232) <= input(14);
output(1, 233) <= input(15);
output(1, 234) <= input(32);
output(1, 235) <= input(34);
output(1, 236) <= input(36);
output(1, 237) <= input(38);
output(1, 238) <= input(40);
output(1, 239) <= input(42);
output(1, 240) <= input(22);
output(1, 241) <= input(23);
output(1, 242) <= input(24);
output(1, 243) <= input(25);
output(1, 244) <= input(26);
output(1, 245) <= input(27);
output(1, 246) <= input(28);
output(1, 247) <= input(29);
output(1, 248) <= input(30);
output(1, 249) <= input(31);
output(1, 250) <= input(33);
output(1, 251) <= input(35);
output(1, 252) <= input(37);
output(1, 253) <= input(39);
output(1, 254) <= input(41);
output(1, 255) <= input(43);
output(2, 0) <= input(46);
output(2, 1) <= input(16);
output(2, 2) <= input(17);
output(2, 3) <= input(18);
output(2, 4) <= input(19);
output(2, 5) <= input(20);
output(2, 6) <= input(21);
output(2, 7) <= input(22);
output(2, 8) <= input(23);
output(2, 9) <= input(24);
output(2, 10) <= input(25);
output(2, 11) <= input(26);
output(2, 12) <= input(27);
output(2, 13) <= input(28);
output(2, 14) <= input(29);
output(2, 15) <= input(30);
output(2, 16) <= input(0);
output(2, 17) <= input(1);
output(2, 18) <= input(2);
output(2, 19) <= input(3);
output(2, 20) <= input(4);
output(2, 21) <= input(5);
output(2, 22) <= input(6);
output(2, 23) <= input(7);
output(2, 24) <= input(8);
output(2, 25) <= input(9);
output(2, 26) <= input(10);
output(2, 27) <= input(11);
output(2, 28) <= input(12);
output(2, 29) <= input(13);
output(2, 30) <= input(14);
output(2, 31) <= input(15);
output(2, 32) <= input(16);
output(2, 33) <= input(17);
output(2, 34) <= input(18);
output(2, 35) <= input(19);
output(2, 36) <= input(20);
output(2, 37) <= input(21);
output(2, 38) <= input(22);
output(2, 39) <= input(23);
output(2, 40) <= input(24);
output(2, 41) <= input(25);
output(2, 42) <= input(26);
output(2, 43) <= input(27);
output(2, 44) <= input(28);
output(2, 45) <= input(29);
output(2, 46) <= input(30);
output(2, 47) <= input(31);
output(2, 48) <= input(1);
output(2, 49) <= input(2);
output(2, 50) <= input(3);
output(2, 51) <= input(4);
output(2, 52) <= input(5);
output(2, 53) <= input(6);
output(2, 54) <= input(7);
output(2, 55) <= input(8);
output(2, 56) <= input(9);
output(2, 57) <= input(10);
output(2, 58) <= input(11);
output(2, 59) <= input(12);
output(2, 60) <= input(13);
output(2, 61) <= input(14);
output(2, 62) <= input(15);
output(2, 63) <= input(32);
output(2, 64) <= input(1);
output(2, 65) <= input(2);
output(2, 66) <= input(3);
output(2, 67) <= input(4);
output(2, 68) <= input(5);
output(2, 69) <= input(6);
output(2, 70) <= input(7);
output(2, 71) <= input(8);
output(2, 72) <= input(9);
output(2, 73) <= input(10);
output(2, 74) <= input(11);
output(2, 75) <= input(12);
output(2, 76) <= input(13);
output(2, 77) <= input(14);
output(2, 78) <= input(15);
output(2, 79) <= input(32);
output(2, 80) <= input(17);
output(2, 81) <= input(18);
output(2, 82) <= input(19);
output(2, 83) <= input(20);
output(2, 84) <= input(21);
output(2, 85) <= input(22);
output(2, 86) <= input(23);
output(2, 87) <= input(24);
output(2, 88) <= input(25);
output(2, 89) <= input(26);
output(2, 90) <= input(27);
output(2, 91) <= input(28);
output(2, 92) <= input(29);
output(2, 93) <= input(30);
output(2, 94) <= input(31);
output(2, 95) <= input(33);
output(2, 96) <= input(2);
output(2, 97) <= input(3);
output(2, 98) <= input(4);
output(2, 99) <= input(5);
output(2, 100) <= input(6);
output(2, 101) <= input(7);
output(2, 102) <= input(8);
output(2, 103) <= input(9);
output(2, 104) <= input(10);
output(2, 105) <= input(11);
output(2, 106) <= input(12);
output(2, 107) <= input(13);
output(2, 108) <= input(14);
output(2, 109) <= input(15);
output(2, 110) <= input(32);
output(2, 111) <= input(34);
output(2, 112) <= input(18);
output(2, 113) <= input(19);
output(2, 114) <= input(20);
output(2, 115) <= input(21);
output(2, 116) <= input(22);
output(2, 117) <= input(23);
output(2, 118) <= input(24);
output(2, 119) <= input(25);
output(2, 120) <= input(26);
output(2, 121) <= input(27);
output(2, 122) <= input(28);
output(2, 123) <= input(29);
output(2, 124) <= input(30);
output(2, 125) <= input(31);
output(2, 126) <= input(33);
output(2, 127) <= input(35);
output(2, 128) <= input(18);
output(2, 129) <= input(19);
output(2, 130) <= input(20);
output(2, 131) <= input(21);
output(2, 132) <= input(22);
output(2, 133) <= input(23);
output(2, 134) <= input(24);
output(2, 135) <= input(25);
output(2, 136) <= input(26);
output(2, 137) <= input(27);
output(2, 138) <= input(28);
output(2, 139) <= input(29);
output(2, 140) <= input(30);
output(2, 141) <= input(31);
output(2, 142) <= input(33);
output(2, 143) <= input(35);
output(2, 144) <= input(3);
output(2, 145) <= input(4);
output(2, 146) <= input(5);
output(2, 147) <= input(6);
output(2, 148) <= input(7);
output(2, 149) <= input(8);
output(2, 150) <= input(9);
output(2, 151) <= input(10);
output(2, 152) <= input(11);
output(2, 153) <= input(12);
output(2, 154) <= input(13);
output(2, 155) <= input(14);
output(2, 156) <= input(15);
output(2, 157) <= input(32);
output(2, 158) <= input(34);
output(2, 159) <= input(36);
output(2, 160) <= input(19);
output(2, 161) <= input(20);
output(2, 162) <= input(21);
output(2, 163) <= input(22);
output(2, 164) <= input(23);
output(2, 165) <= input(24);
output(2, 166) <= input(25);
output(2, 167) <= input(26);
output(2, 168) <= input(27);
output(2, 169) <= input(28);
output(2, 170) <= input(29);
output(2, 171) <= input(30);
output(2, 172) <= input(31);
output(2, 173) <= input(33);
output(2, 174) <= input(35);
output(2, 175) <= input(37);
output(2, 176) <= input(4);
output(2, 177) <= input(5);
output(2, 178) <= input(6);
output(2, 179) <= input(7);
output(2, 180) <= input(8);
output(2, 181) <= input(9);
output(2, 182) <= input(10);
output(2, 183) <= input(11);
output(2, 184) <= input(12);
output(2, 185) <= input(13);
output(2, 186) <= input(14);
output(2, 187) <= input(15);
output(2, 188) <= input(32);
output(2, 189) <= input(34);
output(2, 190) <= input(36);
output(2, 191) <= input(38);
output(2, 192) <= input(4);
output(2, 193) <= input(5);
output(2, 194) <= input(6);
output(2, 195) <= input(7);
output(2, 196) <= input(8);
output(2, 197) <= input(9);
output(2, 198) <= input(10);
output(2, 199) <= input(11);
output(2, 200) <= input(12);
output(2, 201) <= input(13);
output(2, 202) <= input(14);
output(2, 203) <= input(15);
output(2, 204) <= input(32);
output(2, 205) <= input(34);
output(2, 206) <= input(36);
output(2, 207) <= input(38);
output(2, 208) <= input(20);
output(2, 209) <= input(21);
output(2, 210) <= input(22);
output(2, 211) <= input(23);
output(2, 212) <= input(24);
output(2, 213) <= input(25);
output(2, 214) <= input(26);
output(2, 215) <= input(27);
output(2, 216) <= input(28);
output(2, 217) <= input(29);
output(2, 218) <= input(30);
output(2, 219) <= input(31);
output(2, 220) <= input(33);
output(2, 221) <= input(35);
output(2, 222) <= input(37);
output(2, 223) <= input(39);
output(2, 224) <= input(5);
output(2, 225) <= input(6);
output(2, 226) <= input(7);
output(2, 227) <= input(8);
output(2, 228) <= input(9);
output(2, 229) <= input(10);
output(2, 230) <= input(11);
output(2, 231) <= input(12);
output(2, 232) <= input(13);
output(2, 233) <= input(14);
output(2, 234) <= input(15);
output(2, 235) <= input(32);
output(2, 236) <= input(34);
output(2, 237) <= input(36);
output(2, 238) <= input(38);
output(2, 239) <= input(40);
output(2, 240) <= input(21);
output(2, 241) <= input(22);
output(2, 242) <= input(23);
output(2, 243) <= input(24);
output(2, 244) <= input(25);
output(2, 245) <= input(26);
output(2, 246) <= input(27);
output(2, 247) <= input(28);
output(2, 248) <= input(29);
output(2, 249) <= input(30);
output(2, 250) <= input(31);
output(2, 251) <= input(33);
output(2, 252) <= input(35);
output(2, 253) <= input(37);
output(2, 254) <= input(39);
output(2, 255) <= input(41);
output(3, 0) <= input(46);
output(3, 1) <= input(16);
output(3, 2) <= input(17);
output(3, 3) <= input(18);
output(3, 4) <= input(19);
output(3, 5) <= input(20);
output(3, 6) <= input(21);
output(3, 7) <= input(22);
output(3, 8) <= input(23);
output(3, 9) <= input(24);
output(3, 10) <= input(25);
output(3, 11) <= input(26);
output(3, 12) <= input(27);
output(3, 13) <= input(28);
output(3, 14) <= input(29);
output(3, 15) <= input(30);
output(3, 16) <= input(0);
output(3, 17) <= input(1);
output(3, 18) <= input(2);
output(3, 19) <= input(3);
output(3, 20) <= input(4);
output(3, 21) <= input(5);
output(3, 22) <= input(6);
output(3, 23) <= input(7);
output(3, 24) <= input(8);
output(3, 25) <= input(9);
output(3, 26) <= input(10);
output(3, 27) <= input(11);
output(3, 28) <= input(12);
output(3, 29) <= input(13);
output(3, 30) <= input(14);
output(3, 31) <= input(15);
output(3, 32) <= input(0);
output(3, 33) <= input(1);
output(3, 34) <= input(2);
output(3, 35) <= input(3);
output(3, 36) <= input(4);
output(3, 37) <= input(5);
output(3, 38) <= input(6);
output(3, 39) <= input(7);
output(3, 40) <= input(8);
output(3, 41) <= input(9);
output(3, 42) <= input(10);
output(3, 43) <= input(11);
output(3, 44) <= input(12);
output(3, 45) <= input(13);
output(3, 46) <= input(14);
output(3, 47) <= input(15);
output(3, 48) <= input(16);
output(3, 49) <= input(17);
output(3, 50) <= input(18);
output(3, 51) <= input(19);
output(3, 52) <= input(20);
output(3, 53) <= input(21);
output(3, 54) <= input(22);
output(3, 55) <= input(23);
output(3, 56) <= input(24);
output(3, 57) <= input(25);
output(3, 58) <= input(26);
output(3, 59) <= input(27);
output(3, 60) <= input(28);
output(3, 61) <= input(29);
output(3, 62) <= input(30);
output(3, 63) <= input(31);
output(3, 64) <= input(1);
output(3, 65) <= input(2);
output(3, 66) <= input(3);
output(3, 67) <= input(4);
output(3, 68) <= input(5);
output(3, 69) <= input(6);
output(3, 70) <= input(7);
output(3, 71) <= input(8);
output(3, 72) <= input(9);
output(3, 73) <= input(10);
output(3, 74) <= input(11);
output(3, 75) <= input(12);
output(3, 76) <= input(13);
output(3, 77) <= input(14);
output(3, 78) <= input(15);
output(3, 79) <= input(32);
output(3, 80) <= input(1);
output(3, 81) <= input(2);
output(3, 82) <= input(3);
output(3, 83) <= input(4);
output(3, 84) <= input(5);
output(3, 85) <= input(6);
output(3, 86) <= input(7);
output(3, 87) <= input(8);
output(3, 88) <= input(9);
output(3, 89) <= input(10);
output(3, 90) <= input(11);
output(3, 91) <= input(12);
output(3, 92) <= input(13);
output(3, 93) <= input(14);
output(3, 94) <= input(15);
output(3, 95) <= input(32);
output(3, 96) <= input(17);
output(3, 97) <= input(18);
output(3, 98) <= input(19);
output(3, 99) <= input(20);
output(3, 100) <= input(21);
output(3, 101) <= input(22);
output(3, 102) <= input(23);
output(3, 103) <= input(24);
output(3, 104) <= input(25);
output(3, 105) <= input(26);
output(3, 106) <= input(27);
output(3, 107) <= input(28);
output(3, 108) <= input(29);
output(3, 109) <= input(30);
output(3, 110) <= input(31);
output(3, 111) <= input(33);
output(3, 112) <= input(2);
output(3, 113) <= input(3);
output(3, 114) <= input(4);
output(3, 115) <= input(5);
output(3, 116) <= input(6);
output(3, 117) <= input(7);
output(3, 118) <= input(8);
output(3, 119) <= input(9);
output(3, 120) <= input(10);
output(3, 121) <= input(11);
output(3, 122) <= input(12);
output(3, 123) <= input(13);
output(3, 124) <= input(14);
output(3, 125) <= input(15);
output(3, 126) <= input(32);
output(3, 127) <= input(34);
output(3, 128) <= input(2);
output(3, 129) <= input(3);
output(3, 130) <= input(4);
output(3, 131) <= input(5);
output(3, 132) <= input(6);
output(3, 133) <= input(7);
output(3, 134) <= input(8);
output(3, 135) <= input(9);
output(3, 136) <= input(10);
output(3, 137) <= input(11);
output(3, 138) <= input(12);
output(3, 139) <= input(13);
output(3, 140) <= input(14);
output(3, 141) <= input(15);
output(3, 142) <= input(32);
output(3, 143) <= input(34);
output(3, 144) <= input(18);
output(3, 145) <= input(19);
output(3, 146) <= input(20);
output(3, 147) <= input(21);
output(3, 148) <= input(22);
output(3, 149) <= input(23);
output(3, 150) <= input(24);
output(3, 151) <= input(25);
output(3, 152) <= input(26);
output(3, 153) <= input(27);
output(3, 154) <= input(28);
output(3, 155) <= input(29);
output(3, 156) <= input(30);
output(3, 157) <= input(31);
output(3, 158) <= input(33);
output(3, 159) <= input(35);
output(3, 160) <= input(18);
output(3, 161) <= input(19);
output(3, 162) <= input(20);
output(3, 163) <= input(21);
output(3, 164) <= input(22);
output(3, 165) <= input(23);
output(3, 166) <= input(24);
output(3, 167) <= input(25);
output(3, 168) <= input(26);
output(3, 169) <= input(27);
output(3, 170) <= input(28);
output(3, 171) <= input(29);
output(3, 172) <= input(30);
output(3, 173) <= input(31);
output(3, 174) <= input(33);
output(3, 175) <= input(35);
output(3, 176) <= input(3);
output(3, 177) <= input(4);
output(3, 178) <= input(5);
output(3, 179) <= input(6);
output(3, 180) <= input(7);
output(3, 181) <= input(8);
output(3, 182) <= input(9);
output(3, 183) <= input(10);
output(3, 184) <= input(11);
output(3, 185) <= input(12);
output(3, 186) <= input(13);
output(3, 187) <= input(14);
output(3, 188) <= input(15);
output(3, 189) <= input(32);
output(3, 190) <= input(34);
output(3, 191) <= input(36);
output(3, 192) <= input(19);
output(3, 193) <= input(20);
output(3, 194) <= input(21);
output(3, 195) <= input(22);
output(3, 196) <= input(23);
output(3, 197) <= input(24);
output(3, 198) <= input(25);
output(3, 199) <= input(26);
output(3, 200) <= input(27);
output(3, 201) <= input(28);
output(3, 202) <= input(29);
output(3, 203) <= input(30);
output(3, 204) <= input(31);
output(3, 205) <= input(33);
output(3, 206) <= input(35);
output(3, 207) <= input(37);
output(3, 208) <= input(19);
output(3, 209) <= input(20);
output(3, 210) <= input(21);
output(3, 211) <= input(22);
output(3, 212) <= input(23);
output(3, 213) <= input(24);
output(3, 214) <= input(25);
output(3, 215) <= input(26);
output(3, 216) <= input(27);
output(3, 217) <= input(28);
output(3, 218) <= input(29);
output(3, 219) <= input(30);
output(3, 220) <= input(31);
output(3, 221) <= input(33);
output(3, 222) <= input(35);
output(3, 223) <= input(37);
output(3, 224) <= input(4);
output(3, 225) <= input(5);
output(3, 226) <= input(6);
output(3, 227) <= input(7);
output(3, 228) <= input(8);
output(3, 229) <= input(9);
output(3, 230) <= input(10);
output(3, 231) <= input(11);
output(3, 232) <= input(12);
output(3, 233) <= input(13);
output(3, 234) <= input(14);
output(3, 235) <= input(15);
output(3, 236) <= input(32);
output(3, 237) <= input(34);
output(3, 238) <= input(36);
output(3, 239) <= input(38);
output(3, 240) <= input(20);
output(3, 241) <= input(21);
output(3, 242) <= input(22);
output(3, 243) <= input(23);
output(3, 244) <= input(24);
output(3, 245) <= input(25);
output(3, 246) <= input(26);
output(3, 247) <= input(27);
output(3, 248) <= input(28);
output(3, 249) <= input(29);
output(3, 250) <= input(30);
output(3, 251) <= input(31);
output(3, 252) <= input(33);
output(3, 253) <= input(35);
output(3, 254) <= input(37);
output(3, 255) <= input(39);
output(4, 0) <= input(46);
output(4, 1) <= input(16);
output(4, 2) <= input(17);
output(4, 3) <= input(18);
output(4, 4) <= input(19);
output(4, 5) <= input(20);
output(4, 6) <= input(21);
output(4, 7) <= input(22);
output(4, 8) <= input(23);
output(4, 9) <= input(24);
output(4, 10) <= input(25);
output(4, 11) <= input(26);
output(4, 12) <= input(27);
output(4, 13) <= input(28);
output(4, 14) <= input(29);
output(4, 15) <= input(30);
output(4, 16) <= input(0);
output(4, 17) <= input(1);
output(4, 18) <= input(2);
output(4, 19) <= input(3);
output(4, 20) <= input(4);
output(4, 21) <= input(5);
output(4, 22) <= input(6);
output(4, 23) <= input(7);
output(4, 24) <= input(8);
output(4, 25) <= input(9);
output(4, 26) <= input(10);
output(4, 27) <= input(11);
output(4, 28) <= input(12);
output(4, 29) <= input(13);
output(4, 30) <= input(14);
output(4, 31) <= input(15);
output(4, 32) <= input(0);
output(4, 33) <= input(1);
output(4, 34) <= input(2);
output(4, 35) <= input(3);
output(4, 36) <= input(4);
output(4, 37) <= input(5);
output(4, 38) <= input(6);
output(4, 39) <= input(7);
output(4, 40) <= input(8);
output(4, 41) <= input(9);
output(4, 42) <= input(10);
output(4, 43) <= input(11);
output(4, 44) <= input(12);
output(4, 45) <= input(13);
output(4, 46) <= input(14);
output(4, 47) <= input(15);
output(4, 48) <= input(16);
output(4, 49) <= input(17);
output(4, 50) <= input(18);
output(4, 51) <= input(19);
output(4, 52) <= input(20);
output(4, 53) <= input(21);
output(4, 54) <= input(22);
output(4, 55) <= input(23);
output(4, 56) <= input(24);
output(4, 57) <= input(25);
output(4, 58) <= input(26);
output(4, 59) <= input(27);
output(4, 60) <= input(28);
output(4, 61) <= input(29);
output(4, 62) <= input(30);
output(4, 63) <= input(31);
output(4, 64) <= input(16);
output(4, 65) <= input(17);
output(4, 66) <= input(18);
output(4, 67) <= input(19);
output(4, 68) <= input(20);
output(4, 69) <= input(21);
output(4, 70) <= input(22);
output(4, 71) <= input(23);
output(4, 72) <= input(24);
output(4, 73) <= input(25);
output(4, 74) <= input(26);
output(4, 75) <= input(27);
output(4, 76) <= input(28);
output(4, 77) <= input(29);
output(4, 78) <= input(30);
output(4, 79) <= input(31);
output(4, 80) <= input(1);
output(4, 81) <= input(2);
output(4, 82) <= input(3);
output(4, 83) <= input(4);
output(4, 84) <= input(5);
output(4, 85) <= input(6);
output(4, 86) <= input(7);
output(4, 87) <= input(8);
output(4, 88) <= input(9);
output(4, 89) <= input(10);
output(4, 90) <= input(11);
output(4, 91) <= input(12);
output(4, 92) <= input(13);
output(4, 93) <= input(14);
output(4, 94) <= input(15);
output(4, 95) <= input(32);
output(4, 96) <= input(1);
output(4, 97) <= input(2);
output(4, 98) <= input(3);
output(4, 99) <= input(4);
output(4, 100) <= input(5);
output(4, 101) <= input(6);
output(4, 102) <= input(7);
output(4, 103) <= input(8);
output(4, 104) <= input(9);
output(4, 105) <= input(10);
output(4, 106) <= input(11);
output(4, 107) <= input(12);
output(4, 108) <= input(13);
output(4, 109) <= input(14);
output(4, 110) <= input(15);
output(4, 111) <= input(32);
output(4, 112) <= input(17);
output(4, 113) <= input(18);
output(4, 114) <= input(19);
output(4, 115) <= input(20);
output(4, 116) <= input(21);
output(4, 117) <= input(22);
output(4, 118) <= input(23);
output(4, 119) <= input(24);
output(4, 120) <= input(25);
output(4, 121) <= input(26);
output(4, 122) <= input(27);
output(4, 123) <= input(28);
output(4, 124) <= input(29);
output(4, 125) <= input(30);
output(4, 126) <= input(31);
output(4, 127) <= input(33);
output(4, 128) <= input(17);
output(4, 129) <= input(18);
output(4, 130) <= input(19);
output(4, 131) <= input(20);
output(4, 132) <= input(21);
output(4, 133) <= input(22);
output(4, 134) <= input(23);
output(4, 135) <= input(24);
output(4, 136) <= input(25);
output(4, 137) <= input(26);
output(4, 138) <= input(27);
output(4, 139) <= input(28);
output(4, 140) <= input(29);
output(4, 141) <= input(30);
output(4, 142) <= input(31);
output(4, 143) <= input(33);
output(4, 144) <= input(2);
output(4, 145) <= input(3);
output(4, 146) <= input(4);
output(4, 147) <= input(5);
output(4, 148) <= input(6);
output(4, 149) <= input(7);
output(4, 150) <= input(8);
output(4, 151) <= input(9);
output(4, 152) <= input(10);
output(4, 153) <= input(11);
output(4, 154) <= input(12);
output(4, 155) <= input(13);
output(4, 156) <= input(14);
output(4, 157) <= input(15);
output(4, 158) <= input(32);
output(4, 159) <= input(34);
output(4, 160) <= input(2);
output(4, 161) <= input(3);
output(4, 162) <= input(4);
output(4, 163) <= input(5);
output(4, 164) <= input(6);
output(4, 165) <= input(7);
output(4, 166) <= input(8);
output(4, 167) <= input(9);
output(4, 168) <= input(10);
output(4, 169) <= input(11);
output(4, 170) <= input(12);
output(4, 171) <= input(13);
output(4, 172) <= input(14);
output(4, 173) <= input(15);
output(4, 174) <= input(32);
output(4, 175) <= input(34);
output(4, 176) <= input(18);
output(4, 177) <= input(19);
output(4, 178) <= input(20);
output(4, 179) <= input(21);
output(4, 180) <= input(22);
output(4, 181) <= input(23);
output(4, 182) <= input(24);
output(4, 183) <= input(25);
output(4, 184) <= input(26);
output(4, 185) <= input(27);
output(4, 186) <= input(28);
output(4, 187) <= input(29);
output(4, 188) <= input(30);
output(4, 189) <= input(31);
output(4, 190) <= input(33);
output(4, 191) <= input(35);
output(4, 192) <= input(18);
output(4, 193) <= input(19);
output(4, 194) <= input(20);
output(4, 195) <= input(21);
output(4, 196) <= input(22);
output(4, 197) <= input(23);
output(4, 198) <= input(24);
output(4, 199) <= input(25);
output(4, 200) <= input(26);
output(4, 201) <= input(27);
output(4, 202) <= input(28);
output(4, 203) <= input(29);
output(4, 204) <= input(30);
output(4, 205) <= input(31);
output(4, 206) <= input(33);
output(4, 207) <= input(35);
output(4, 208) <= input(3);
output(4, 209) <= input(4);
output(4, 210) <= input(5);
output(4, 211) <= input(6);
output(4, 212) <= input(7);
output(4, 213) <= input(8);
output(4, 214) <= input(9);
output(4, 215) <= input(10);
output(4, 216) <= input(11);
output(4, 217) <= input(12);
output(4, 218) <= input(13);
output(4, 219) <= input(14);
output(4, 220) <= input(15);
output(4, 221) <= input(32);
output(4, 222) <= input(34);
output(4, 223) <= input(36);
output(4, 224) <= input(3);
output(4, 225) <= input(4);
output(4, 226) <= input(5);
output(4, 227) <= input(6);
output(4, 228) <= input(7);
output(4, 229) <= input(8);
output(4, 230) <= input(9);
output(4, 231) <= input(10);
output(4, 232) <= input(11);
output(4, 233) <= input(12);
output(4, 234) <= input(13);
output(4, 235) <= input(14);
output(4, 236) <= input(15);
output(4, 237) <= input(32);
output(4, 238) <= input(34);
output(4, 239) <= input(36);
output(4, 240) <= input(19);
output(4, 241) <= input(20);
output(4, 242) <= input(21);
output(4, 243) <= input(22);
output(4, 244) <= input(23);
output(4, 245) <= input(24);
output(4, 246) <= input(25);
output(4, 247) <= input(26);
output(4, 248) <= input(27);
output(4, 249) <= input(28);
output(4, 250) <= input(29);
output(4, 251) <= input(30);
output(4, 252) <= input(31);
output(4, 253) <= input(33);
output(4, 254) <= input(35);
output(4, 255) <= input(37);
output(5, 0) <= input(46);
output(5, 1) <= input(16);
output(5, 2) <= input(17);
output(5, 3) <= input(18);
output(5, 4) <= input(19);
output(5, 5) <= input(20);
output(5, 6) <= input(21);
output(5, 7) <= input(22);
output(5, 8) <= input(23);
output(5, 9) <= input(24);
output(5, 10) <= input(25);
output(5, 11) <= input(26);
output(5, 12) <= input(27);
output(5, 13) <= input(28);
output(5, 14) <= input(29);
output(5, 15) <= input(30);
output(5, 16) <= input(46);
output(5, 17) <= input(16);
output(5, 18) <= input(17);
output(5, 19) <= input(18);
output(5, 20) <= input(19);
output(5, 21) <= input(20);
output(5, 22) <= input(21);
output(5, 23) <= input(22);
output(5, 24) <= input(23);
output(5, 25) <= input(24);
output(5, 26) <= input(25);
output(5, 27) <= input(26);
output(5, 28) <= input(27);
output(5, 29) <= input(28);
output(5, 30) <= input(29);
output(5, 31) <= input(30);
output(5, 32) <= input(0);
output(5, 33) <= input(1);
output(5, 34) <= input(2);
output(5, 35) <= input(3);
output(5, 36) <= input(4);
output(5, 37) <= input(5);
output(5, 38) <= input(6);
output(5, 39) <= input(7);
output(5, 40) <= input(8);
output(5, 41) <= input(9);
output(5, 42) <= input(10);
output(5, 43) <= input(11);
output(5, 44) <= input(12);
output(5, 45) <= input(13);
output(5, 46) <= input(14);
output(5, 47) <= input(15);
output(5, 48) <= input(0);
output(5, 49) <= input(1);
output(5, 50) <= input(2);
output(5, 51) <= input(3);
output(5, 52) <= input(4);
output(5, 53) <= input(5);
output(5, 54) <= input(6);
output(5, 55) <= input(7);
output(5, 56) <= input(8);
output(5, 57) <= input(9);
output(5, 58) <= input(10);
output(5, 59) <= input(11);
output(5, 60) <= input(12);
output(5, 61) <= input(13);
output(5, 62) <= input(14);
output(5, 63) <= input(15);
output(5, 64) <= input(0);
output(5, 65) <= input(1);
output(5, 66) <= input(2);
output(5, 67) <= input(3);
output(5, 68) <= input(4);
output(5, 69) <= input(5);
output(5, 70) <= input(6);
output(5, 71) <= input(7);
output(5, 72) <= input(8);
output(5, 73) <= input(9);
output(5, 74) <= input(10);
output(5, 75) <= input(11);
output(5, 76) <= input(12);
output(5, 77) <= input(13);
output(5, 78) <= input(14);
output(5, 79) <= input(15);
output(5, 80) <= input(16);
output(5, 81) <= input(17);
output(5, 82) <= input(18);
output(5, 83) <= input(19);
output(5, 84) <= input(20);
output(5, 85) <= input(21);
output(5, 86) <= input(22);
output(5, 87) <= input(23);
output(5, 88) <= input(24);
output(5, 89) <= input(25);
output(5, 90) <= input(26);
output(5, 91) <= input(27);
output(5, 92) <= input(28);
output(5, 93) <= input(29);
output(5, 94) <= input(30);
output(5, 95) <= input(31);
output(5, 96) <= input(16);
output(5, 97) <= input(17);
output(5, 98) <= input(18);
output(5, 99) <= input(19);
output(5, 100) <= input(20);
output(5, 101) <= input(21);
output(5, 102) <= input(22);
output(5, 103) <= input(23);
output(5, 104) <= input(24);
output(5, 105) <= input(25);
output(5, 106) <= input(26);
output(5, 107) <= input(27);
output(5, 108) <= input(28);
output(5, 109) <= input(29);
output(5, 110) <= input(30);
output(5, 111) <= input(31);
output(5, 112) <= input(1);
output(5, 113) <= input(2);
output(5, 114) <= input(3);
output(5, 115) <= input(4);
output(5, 116) <= input(5);
output(5, 117) <= input(6);
output(5, 118) <= input(7);
output(5, 119) <= input(8);
output(5, 120) <= input(9);
output(5, 121) <= input(10);
output(5, 122) <= input(11);
output(5, 123) <= input(12);
output(5, 124) <= input(13);
output(5, 125) <= input(14);
output(5, 126) <= input(15);
output(5, 127) <= input(32);
output(5, 128) <= input(1);
output(5, 129) <= input(2);
output(5, 130) <= input(3);
output(5, 131) <= input(4);
output(5, 132) <= input(5);
output(5, 133) <= input(6);
output(5, 134) <= input(7);
output(5, 135) <= input(8);
output(5, 136) <= input(9);
output(5, 137) <= input(10);
output(5, 138) <= input(11);
output(5, 139) <= input(12);
output(5, 140) <= input(13);
output(5, 141) <= input(14);
output(5, 142) <= input(15);
output(5, 143) <= input(32);
output(5, 144) <= input(1);
output(5, 145) <= input(2);
output(5, 146) <= input(3);
output(5, 147) <= input(4);
output(5, 148) <= input(5);
output(5, 149) <= input(6);
output(5, 150) <= input(7);
output(5, 151) <= input(8);
output(5, 152) <= input(9);
output(5, 153) <= input(10);
output(5, 154) <= input(11);
output(5, 155) <= input(12);
output(5, 156) <= input(13);
output(5, 157) <= input(14);
output(5, 158) <= input(15);
output(5, 159) <= input(32);
output(5, 160) <= input(17);
output(5, 161) <= input(18);
output(5, 162) <= input(19);
output(5, 163) <= input(20);
output(5, 164) <= input(21);
output(5, 165) <= input(22);
output(5, 166) <= input(23);
output(5, 167) <= input(24);
output(5, 168) <= input(25);
output(5, 169) <= input(26);
output(5, 170) <= input(27);
output(5, 171) <= input(28);
output(5, 172) <= input(29);
output(5, 173) <= input(30);
output(5, 174) <= input(31);
output(5, 175) <= input(33);
output(5, 176) <= input(17);
output(5, 177) <= input(18);
output(5, 178) <= input(19);
output(5, 179) <= input(20);
output(5, 180) <= input(21);
output(5, 181) <= input(22);
output(5, 182) <= input(23);
output(5, 183) <= input(24);
output(5, 184) <= input(25);
output(5, 185) <= input(26);
output(5, 186) <= input(27);
output(5, 187) <= input(28);
output(5, 188) <= input(29);
output(5, 189) <= input(30);
output(5, 190) <= input(31);
output(5, 191) <= input(33);
output(5, 192) <= input(17);
output(5, 193) <= input(18);
output(5, 194) <= input(19);
output(5, 195) <= input(20);
output(5, 196) <= input(21);
output(5, 197) <= input(22);
output(5, 198) <= input(23);
output(5, 199) <= input(24);
output(5, 200) <= input(25);
output(5, 201) <= input(26);
output(5, 202) <= input(27);
output(5, 203) <= input(28);
output(5, 204) <= input(29);
output(5, 205) <= input(30);
output(5, 206) <= input(31);
output(5, 207) <= input(33);
output(5, 208) <= input(2);
output(5, 209) <= input(3);
output(5, 210) <= input(4);
output(5, 211) <= input(5);
output(5, 212) <= input(6);
output(5, 213) <= input(7);
output(5, 214) <= input(8);
output(5, 215) <= input(9);
output(5, 216) <= input(10);
output(5, 217) <= input(11);
output(5, 218) <= input(12);
output(5, 219) <= input(13);
output(5, 220) <= input(14);
output(5, 221) <= input(15);
output(5, 222) <= input(32);
output(5, 223) <= input(34);
output(5, 224) <= input(2);
output(5, 225) <= input(3);
output(5, 226) <= input(4);
output(5, 227) <= input(5);
output(5, 228) <= input(6);
output(5, 229) <= input(7);
output(5, 230) <= input(8);
output(5, 231) <= input(9);
output(5, 232) <= input(10);
output(5, 233) <= input(11);
output(5, 234) <= input(12);
output(5, 235) <= input(13);
output(5, 236) <= input(14);
output(5, 237) <= input(15);
output(5, 238) <= input(32);
output(5, 239) <= input(34);
output(5, 240) <= input(18);
output(5, 241) <= input(19);
output(5, 242) <= input(20);
output(5, 243) <= input(21);
output(5, 244) <= input(22);
output(5, 245) <= input(23);
output(5, 246) <= input(24);
output(5, 247) <= input(25);
output(5, 248) <= input(26);
output(5, 249) <= input(27);
output(5, 250) <= input(28);
output(5, 251) <= input(29);
output(5, 252) <= input(30);
output(5, 253) <= input(31);
output(5, 254) <= input(33);
output(5, 255) <= input(35);
when "0010" =>
output(0, 0) <= input(0);
output(0, 1) <= input(1);
output(0, 2) <= input(2);
output(0, 3) <= input(3);
output(0, 4) <= input(4);
output(0, 5) <= input(5);
output(0, 6) <= input(6);
output(0, 7) <= input(7);
output(0, 8) <= input(8);
output(0, 9) <= input(9);
output(0, 10) <= input(10);
output(0, 11) <= input(11);
output(0, 12) <= input(12);
output(0, 13) <= input(13);
output(0, 14) <= input(14);
output(0, 15) <= input(15);
output(0, 16) <= input(0);
output(0, 17) <= input(1);
output(0, 18) <= input(2);
output(0, 19) <= input(3);
output(0, 20) <= input(4);
output(0, 21) <= input(5);
output(0, 22) <= input(6);
output(0, 23) <= input(7);
output(0, 24) <= input(8);
output(0, 25) <= input(9);
output(0, 26) <= input(10);
output(0, 27) <= input(11);
output(0, 28) <= input(12);
output(0, 29) <= input(13);
output(0, 30) <= input(14);
output(0, 31) <= input(15);
output(0, 32) <= input(0);
output(0, 33) <= input(1);
output(0, 34) <= input(2);
output(0, 35) <= input(3);
output(0, 36) <= input(4);
output(0, 37) <= input(5);
output(0, 38) <= input(6);
output(0, 39) <= input(7);
output(0, 40) <= input(8);
output(0, 41) <= input(9);
output(0, 42) <= input(10);
output(0, 43) <= input(11);
output(0, 44) <= input(12);
output(0, 45) <= input(13);
output(0, 46) <= input(14);
output(0, 47) <= input(15);
output(0, 48) <= input(16);
output(0, 49) <= input(17);
output(0, 50) <= input(18);
output(0, 51) <= input(19);
output(0, 52) <= input(20);
output(0, 53) <= input(21);
output(0, 54) <= input(22);
output(0, 55) <= input(23);
output(0, 56) <= input(24);
output(0, 57) <= input(25);
output(0, 58) <= input(26);
output(0, 59) <= input(27);
output(0, 60) <= input(28);
output(0, 61) <= input(29);
output(0, 62) <= input(30);
output(0, 63) <= input(31);
output(0, 64) <= input(16);
output(0, 65) <= input(17);
output(0, 66) <= input(18);
output(0, 67) <= input(19);
output(0, 68) <= input(20);
output(0, 69) <= input(21);
output(0, 70) <= input(22);
output(0, 71) <= input(23);
output(0, 72) <= input(24);
output(0, 73) <= input(25);
output(0, 74) <= input(26);
output(0, 75) <= input(27);
output(0, 76) <= input(28);
output(0, 77) <= input(29);
output(0, 78) <= input(30);
output(0, 79) <= input(31);
output(0, 80) <= input(16);
output(0, 81) <= input(17);
output(0, 82) <= input(18);
output(0, 83) <= input(19);
output(0, 84) <= input(20);
output(0, 85) <= input(21);
output(0, 86) <= input(22);
output(0, 87) <= input(23);
output(0, 88) <= input(24);
output(0, 89) <= input(25);
output(0, 90) <= input(26);
output(0, 91) <= input(27);
output(0, 92) <= input(28);
output(0, 93) <= input(29);
output(0, 94) <= input(30);
output(0, 95) <= input(31);
output(0, 96) <= input(16);
output(0, 97) <= input(17);
output(0, 98) <= input(18);
output(0, 99) <= input(19);
output(0, 100) <= input(20);
output(0, 101) <= input(21);
output(0, 102) <= input(22);
output(0, 103) <= input(23);
output(0, 104) <= input(24);
output(0, 105) <= input(25);
output(0, 106) <= input(26);
output(0, 107) <= input(27);
output(0, 108) <= input(28);
output(0, 109) <= input(29);
output(0, 110) <= input(30);
output(0, 111) <= input(31);
output(0, 112) <= input(1);
output(0, 113) <= input(2);
output(0, 114) <= input(3);
output(0, 115) <= input(4);
output(0, 116) <= input(5);
output(0, 117) <= input(6);
output(0, 118) <= input(7);
output(0, 119) <= input(8);
output(0, 120) <= input(9);
output(0, 121) <= input(10);
output(0, 122) <= input(11);
output(0, 123) <= input(12);
output(0, 124) <= input(13);
output(0, 125) <= input(14);
output(0, 126) <= input(15);
output(0, 127) <= input(32);
output(0, 128) <= input(1);
output(0, 129) <= input(2);
output(0, 130) <= input(3);
output(0, 131) <= input(4);
output(0, 132) <= input(5);
output(0, 133) <= input(6);
output(0, 134) <= input(7);
output(0, 135) <= input(8);
output(0, 136) <= input(9);
output(0, 137) <= input(10);
output(0, 138) <= input(11);
output(0, 139) <= input(12);
output(0, 140) <= input(13);
output(0, 141) <= input(14);
output(0, 142) <= input(15);
output(0, 143) <= input(32);
output(0, 144) <= input(1);
output(0, 145) <= input(2);
output(0, 146) <= input(3);
output(0, 147) <= input(4);
output(0, 148) <= input(5);
output(0, 149) <= input(6);
output(0, 150) <= input(7);
output(0, 151) <= input(8);
output(0, 152) <= input(9);
output(0, 153) <= input(10);
output(0, 154) <= input(11);
output(0, 155) <= input(12);
output(0, 156) <= input(13);
output(0, 157) <= input(14);
output(0, 158) <= input(15);
output(0, 159) <= input(32);
output(0, 160) <= input(1);
output(0, 161) <= input(2);
output(0, 162) <= input(3);
output(0, 163) <= input(4);
output(0, 164) <= input(5);
output(0, 165) <= input(6);
output(0, 166) <= input(7);
output(0, 167) <= input(8);
output(0, 168) <= input(9);
output(0, 169) <= input(10);
output(0, 170) <= input(11);
output(0, 171) <= input(12);
output(0, 172) <= input(13);
output(0, 173) <= input(14);
output(0, 174) <= input(15);
output(0, 175) <= input(32);
output(0, 176) <= input(17);
output(0, 177) <= input(18);
output(0, 178) <= input(19);
output(0, 179) <= input(20);
output(0, 180) <= input(21);
output(0, 181) <= input(22);
output(0, 182) <= input(23);
output(0, 183) <= input(24);
output(0, 184) <= input(25);
output(0, 185) <= input(26);
output(0, 186) <= input(27);
output(0, 187) <= input(28);
output(0, 188) <= input(29);
output(0, 189) <= input(30);
output(0, 190) <= input(31);
output(0, 191) <= input(33);
output(0, 192) <= input(17);
output(0, 193) <= input(18);
output(0, 194) <= input(19);
output(0, 195) <= input(20);
output(0, 196) <= input(21);
output(0, 197) <= input(22);
output(0, 198) <= input(23);
output(0, 199) <= input(24);
output(0, 200) <= input(25);
output(0, 201) <= input(26);
output(0, 202) <= input(27);
output(0, 203) <= input(28);
output(0, 204) <= input(29);
output(0, 205) <= input(30);
output(0, 206) <= input(31);
output(0, 207) <= input(33);
output(0, 208) <= input(17);
output(0, 209) <= input(18);
output(0, 210) <= input(19);
output(0, 211) <= input(20);
output(0, 212) <= input(21);
output(0, 213) <= input(22);
output(0, 214) <= input(23);
output(0, 215) <= input(24);
output(0, 216) <= input(25);
output(0, 217) <= input(26);
output(0, 218) <= input(27);
output(0, 219) <= input(28);
output(0, 220) <= input(29);
output(0, 221) <= input(30);
output(0, 222) <= input(31);
output(0, 223) <= input(33);
output(0, 224) <= input(17);
output(0, 225) <= input(18);
output(0, 226) <= input(19);
output(0, 227) <= input(20);
output(0, 228) <= input(21);
output(0, 229) <= input(22);
output(0, 230) <= input(23);
output(0, 231) <= input(24);
output(0, 232) <= input(25);
output(0, 233) <= input(26);
output(0, 234) <= input(27);
output(0, 235) <= input(28);
output(0, 236) <= input(29);
output(0, 237) <= input(30);
output(0, 238) <= input(31);
output(0, 239) <= input(33);
output(0, 240) <= input(2);
output(0, 241) <= input(3);
output(0, 242) <= input(4);
output(0, 243) <= input(5);
output(0, 244) <= input(6);
output(0, 245) <= input(7);
output(0, 246) <= input(8);
output(0, 247) <= input(9);
output(0, 248) <= input(10);
output(0, 249) <= input(11);
output(0, 250) <= input(12);
output(0, 251) <= input(13);
output(0, 252) <= input(14);
output(0, 253) <= input(15);
output(0, 254) <= input(32);
output(0, 255) <= input(34);
output(1, 0) <= input(0);
output(1, 1) <= input(1);
output(1, 2) <= input(2);
output(1, 3) <= input(3);
output(1, 4) <= input(4);
output(1, 5) <= input(5);
output(1, 6) <= input(6);
output(1, 7) <= input(7);
output(1, 8) <= input(8);
output(1, 9) <= input(9);
output(1, 10) <= input(10);
output(1, 11) <= input(11);
output(1, 12) <= input(12);
output(1, 13) <= input(13);
output(1, 14) <= input(14);
output(1, 15) <= input(15);
output(1, 16) <= input(0);
output(1, 17) <= input(1);
output(1, 18) <= input(2);
output(1, 19) <= input(3);
output(1, 20) <= input(4);
output(1, 21) <= input(5);
output(1, 22) <= input(6);
output(1, 23) <= input(7);
output(1, 24) <= input(8);
output(1, 25) <= input(9);
output(1, 26) <= input(10);
output(1, 27) <= input(11);
output(1, 28) <= input(12);
output(1, 29) <= input(13);
output(1, 30) <= input(14);
output(1, 31) <= input(15);
output(1, 32) <= input(0);
output(1, 33) <= input(1);
output(1, 34) <= input(2);
output(1, 35) <= input(3);
output(1, 36) <= input(4);
output(1, 37) <= input(5);
output(1, 38) <= input(6);
output(1, 39) <= input(7);
output(1, 40) <= input(8);
output(1, 41) <= input(9);
output(1, 42) <= input(10);
output(1, 43) <= input(11);
output(1, 44) <= input(12);
output(1, 45) <= input(13);
output(1, 46) <= input(14);
output(1, 47) <= input(15);
output(1, 48) <= input(0);
output(1, 49) <= input(1);
output(1, 50) <= input(2);
output(1, 51) <= input(3);
output(1, 52) <= input(4);
output(1, 53) <= input(5);
output(1, 54) <= input(6);
output(1, 55) <= input(7);
output(1, 56) <= input(8);
output(1, 57) <= input(9);
output(1, 58) <= input(10);
output(1, 59) <= input(11);
output(1, 60) <= input(12);
output(1, 61) <= input(13);
output(1, 62) <= input(14);
output(1, 63) <= input(15);
output(1, 64) <= input(0);
output(1, 65) <= input(1);
output(1, 66) <= input(2);
output(1, 67) <= input(3);
output(1, 68) <= input(4);
output(1, 69) <= input(5);
output(1, 70) <= input(6);
output(1, 71) <= input(7);
output(1, 72) <= input(8);
output(1, 73) <= input(9);
output(1, 74) <= input(10);
output(1, 75) <= input(11);
output(1, 76) <= input(12);
output(1, 77) <= input(13);
output(1, 78) <= input(14);
output(1, 79) <= input(15);
output(1, 80) <= input(16);
output(1, 81) <= input(17);
output(1, 82) <= input(18);
output(1, 83) <= input(19);
output(1, 84) <= input(20);
output(1, 85) <= input(21);
output(1, 86) <= input(22);
output(1, 87) <= input(23);
output(1, 88) <= input(24);
output(1, 89) <= input(25);
output(1, 90) <= input(26);
output(1, 91) <= input(27);
output(1, 92) <= input(28);
output(1, 93) <= input(29);
output(1, 94) <= input(30);
output(1, 95) <= input(31);
output(1, 96) <= input(16);
output(1, 97) <= input(17);
output(1, 98) <= input(18);
output(1, 99) <= input(19);
output(1, 100) <= input(20);
output(1, 101) <= input(21);
output(1, 102) <= input(22);
output(1, 103) <= input(23);
output(1, 104) <= input(24);
output(1, 105) <= input(25);
output(1, 106) <= input(26);
output(1, 107) <= input(27);
output(1, 108) <= input(28);
output(1, 109) <= input(29);
output(1, 110) <= input(30);
output(1, 111) <= input(31);
output(1, 112) <= input(16);
output(1, 113) <= input(17);
output(1, 114) <= input(18);
output(1, 115) <= input(19);
output(1, 116) <= input(20);
output(1, 117) <= input(21);
output(1, 118) <= input(22);
output(1, 119) <= input(23);
output(1, 120) <= input(24);
output(1, 121) <= input(25);
output(1, 122) <= input(26);
output(1, 123) <= input(27);
output(1, 124) <= input(28);
output(1, 125) <= input(29);
output(1, 126) <= input(30);
output(1, 127) <= input(31);
output(1, 128) <= input(16);
output(1, 129) <= input(17);
output(1, 130) <= input(18);
output(1, 131) <= input(19);
output(1, 132) <= input(20);
output(1, 133) <= input(21);
output(1, 134) <= input(22);
output(1, 135) <= input(23);
output(1, 136) <= input(24);
output(1, 137) <= input(25);
output(1, 138) <= input(26);
output(1, 139) <= input(27);
output(1, 140) <= input(28);
output(1, 141) <= input(29);
output(1, 142) <= input(30);
output(1, 143) <= input(31);
output(1, 144) <= input(16);
output(1, 145) <= input(17);
output(1, 146) <= input(18);
output(1, 147) <= input(19);
output(1, 148) <= input(20);
output(1, 149) <= input(21);
output(1, 150) <= input(22);
output(1, 151) <= input(23);
output(1, 152) <= input(24);
output(1, 153) <= input(25);
output(1, 154) <= input(26);
output(1, 155) <= input(27);
output(1, 156) <= input(28);
output(1, 157) <= input(29);
output(1, 158) <= input(30);
output(1, 159) <= input(31);
output(1, 160) <= input(1);
output(1, 161) <= input(2);
output(1, 162) <= input(3);
output(1, 163) <= input(4);
output(1, 164) <= input(5);
output(1, 165) <= input(6);
output(1, 166) <= input(7);
output(1, 167) <= input(8);
output(1, 168) <= input(9);
output(1, 169) <= input(10);
output(1, 170) <= input(11);
output(1, 171) <= input(12);
output(1, 172) <= input(13);
output(1, 173) <= input(14);
output(1, 174) <= input(15);
output(1, 175) <= input(32);
output(1, 176) <= input(1);
output(1, 177) <= input(2);
output(1, 178) <= input(3);
output(1, 179) <= input(4);
output(1, 180) <= input(5);
output(1, 181) <= input(6);
output(1, 182) <= input(7);
output(1, 183) <= input(8);
output(1, 184) <= input(9);
output(1, 185) <= input(10);
output(1, 186) <= input(11);
output(1, 187) <= input(12);
output(1, 188) <= input(13);
output(1, 189) <= input(14);
output(1, 190) <= input(15);
output(1, 191) <= input(32);
output(1, 192) <= input(1);
output(1, 193) <= input(2);
output(1, 194) <= input(3);
output(1, 195) <= input(4);
output(1, 196) <= input(5);
output(1, 197) <= input(6);
output(1, 198) <= input(7);
output(1, 199) <= input(8);
output(1, 200) <= input(9);
output(1, 201) <= input(10);
output(1, 202) <= input(11);
output(1, 203) <= input(12);
output(1, 204) <= input(13);
output(1, 205) <= input(14);
output(1, 206) <= input(15);
output(1, 207) <= input(32);
output(1, 208) <= input(1);
output(1, 209) <= input(2);
output(1, 210) <= input(3);
output(1, 211) <= input(4);
output(1, 212) <= input(5);
output(1, 213) <= input(6);
output(1, 214) <= input(7);
output(1, 215) <= input(8);
output(1, 216) <= input(9);
output(1, 217) <= input(10);
output(1, 218) <= input(11);
output(1, 219) <= input(12);
output(1, 220) <= input(13);
output(1, 221) <= input(14);
output(1, 222) <= input(15);
output(1, 223) <= input(32);
output(1, 224) <= input(1);
output(1, 225) <= input(2);
output(1, 226) <= input(3);
output(1, 227) <= input(4);
output(1, 228) <= input(5);
output(1, 229) <= input(6);
output(1, 230) <= input(7);
output(1, 231) <= input(8);
output(1, 232) <= input(9);
output(1, 233) <= input(10);
output(1, 234) <= input(11);
output(1, 235) <= input(12);
output(1, 236) <= input(13);
output(1, 237) <= input(14);
output(1, 238) <= input(15);
output(1, 239) <= input(32);
output(1, 240) <= input(17);
output(1, 241) <= input(18);
output(1, 242) <= input(19);
output(1, 243) <= input(20);
output(1, 244) <= input(21);
output(1, 245) <= input(22);
output(1, 246) <= input(23);
output(1, 247) <= input(24);
output(1, 248) <= input(25);
output(1, 249) <= input(26);
output(1, 250) <= input(27);
output(1, 251) <= input(28);
output(1, 252) <= input(29);
output(1, 253) <= input(30);
output(1, 254) <= input(31);
output(1, 255) <= input(33);
output(2, 0) <= input(0);
output(2, 1) <= input(1);
output(2, 2) <= input(2);
output(2, 3) <= input(3);
output(2, 4) <= input(4);
output(2, 5) <= input(5);
output(2, 6) <= input(6);
output(2, 7) <= input(7);
output(2, 8) <= input(8);
output(2, 9) <= input(9);
output(2, 10) <= input(10);
output(2, 11) <= input(11);
output(2, 12) <= input(12);
output(2, 13) <= input(13);
output(2, 14) <= input(14);
output(2, 15) <= input(15);
output(2, 16) <= input(0);
output(2, 17) <= input(1);
output(2, 18) <= input(2);
output(2, 19) <= input(3);
output(2, 20) <= input(4);
output(2, 21) <= input(5);
output(2, 22) <= input(6);
output(2, 23) <= input(7);
output(2, 24) <= input(8);
output(2, 25) <= input(9);
output(2, 26) <= input(10);
output(2, 27) <= input(11);
output(2, 28) <= input(12);
output(2, 29) <= input(13);
output(2, 30) <= input(14);
output(2, 31) <= input(15);
output(2, 32) <= input(0);
output(2, 33) <= input(1);
output(2, 34) <= input(2);
output(2, 35) <= input(3);
output(2, 36) <= input(4);
output(2, 37) <= input(5);
output(2, 38) <= input(6);
output(2, 39) <= input(7);
output(2, 40) <= input(8);
output(2, 41) <= input(9);
output(2, 42) <= input(10);
output(2, 43) <= input(11);
output(2, 44) <= input(12);
output(2, 45) <= input(13);
output(2, 46) <= input(14);
output(2, 47) <= input(15);
output(2, 48) <= input(0);
output(2, 49) <= input(1);
output(2, 50) <= input(2);
output(2, 51) <= input(3);
output(2, 52) <= input(4);
output(2, 53) <= input(5);
output(2, 54) <= input(6);
output(2, 55) <= input(7);
output(2, 56) <= input(8);
output(2, 57) <= input(9);
output(2, 58) <= input(10);
output(2, 59) <= input(11);
output(2, 60) <= input(12);
output(2, 61) <= input(13);
output(2, 62) <= input(14);
output(2, 63) <= input(15);
output(2, 64) <= input(0);
output(2, 65) <= input(1);
output(2, 66) <= input(2);
output(2, 67) <= input(3);
output(2, 68) <= input(4);
output(2, 69) <= input(5);
output(2, 70) <= input(6);
output(2, 71) <= input(7);
output(2, 72) <= input(8);
output(2, 73) <= input(9);
output(2, 74) <= input(10);
output(2, 75) <= input(11);
output(2, 76) <= input(12);
output(2, 77) <= input(13);
output(2, 78) <= input(14);
output(2, 79) <= input(15);
output(2, 80) <= input(0);
output(2, 81) <= input(1);
output(2, 82) <= input(2);
output(2, 83) <= input(3);
output(2, 84) <= input(4);
output(2, 85) <= input(5);
output(2, 86) <= input(6);
output(2, 87) <= input(7);
output(2, 88) <= input(8);
output(2, 89) <= input(9);
output(2, 90) <= input(10);
output(2, 91) <= input(11);
output(2, 92) <= input(12);
output(2, 93) <= input(13);
output(2, 94) <= input(14);
output(2, 95) <= input(15);
output(2, 96) <= input(0);
output(2, 97) <= input(1);
output(2, 98) <= input(2);
output(2, 99) <= input(3);
output(2, 100) <= input(4);
output(2, 101) <= input(5);
output(2, 102) <= input(6);
output(2, 103) <= input(7);
output(2, 104) <= input(8);
output(2, 105) <= input(9);
output(2, 106) <= input(10);
output(2, 107) <= input(11);
output(2, 108) <= input(12);
output(2, 109) <= input(13);
output(2, 110) <= input(14);
output(2, 111) <= input(15);
output(2, 112) <= input(16);
output(2, 113) <= input(17);
output(2, 114) <= input(18);
output(2, 115) <= input(19);
output(2, 116) <= input(20);
output(2, 117) <= input(21);
output(2, 118) <= input(22);
output(2, 119) <= input(23);
output(2, 120) <= input(24);
output(2, 121) <= input(25);
output(2, 122) <= input(26);
output(2, 123) <= input(27);
output(2, 124) <= input(28);
output(2, 125) <= input(29);
output(2, 126) <= input(30);
output(2, 127) <= input(31);
output(2, 128) <= input(16);
output(2, 129) <= input(17);
output(2, 130) <= input(18);
output(2, 131) <= input(19);
output(2, 132) <= input(20);
output(2, 133) <= input(21);
output(2, 134) <= input(22);
output(2, 135) <= input(23);
output(2, 136) <= input(24);
output(2, 137) <= input(25);
output(2, 138) <= input(26);
output(2, 139) <= input(27);
output(2, 140) <= input(28);
output(2, 141) <= input(29);
output(2, 142) <= input(30);
output(2, 143) <= input(31);
output(2, 144) <= input(16);
output(2, 145) <= input(17);
output(2, 146) <= input(18);
output(2, 147) <= input(19);
output(2, 148) <= input(20);
output(2, 149) <= input(21);
output(2, 150) <= input(22);
output(2, 151) <= input(23);
output(2, 152) <= input(24);
output(2, 153) <= input(25);
output(2, 154) <= input(26);
output(2, 155) <= input(27);
output(2, 156) <= input(28);
output(2, 157) <= input(29);
output(2, 158) <= input(30);
output(2, 159) <= input(31);
output(2, 160) <= input(16);
output(2, 161) <= input(17);
output(2, 162) <= input(18);
output(2, 163) <= input(19);
output(2, 164) <= input(20);
output(2, 165) <= input(21);
output(2, 166) <= input(22);
output(2, 167) <= input(23);
output(2, 168) <= input(24);
output(2, 169) <= input(25);
output(2, 170) <= input(26);
output(2, 171) <= input(27);
output(2, 172) <= input(28);
output(2, 173) <= input(29);
output(2, 174) <= input(30);
output(2, 175) <= input(31);
output(2, 176) <= input(16);
output(2, 177) <= input(17);
output(2, 178) <= input(18);
output(2, 179) <= input(19);
output(2, 180) <= input(20);
output(2, 181) <= input(21);
output(2, 182) <= input(22);
output(2, 183) <= input(23);
output(2, 184) <= input(24);
output(2, 185) <= input(25);
output(2, 186) <= input(26);
output(2, 187) <= input(27);
output(2, 188) <= input(28);
output(2, 189) <= input(29);
output(2, 190) <= input(30);
output(2, 191) <= input(31);
output(2, 192) <= input(16);
output(2, 193) <= input(17);
output(2, 194) <= input(18);
output(2, 195) <= input(19);
output(2, 196) <= input(20);
output(2, 197) <= input(21);
output(2, 198) <= input(22);
output(2, 199) <= input(23);
output(2, 200) <= input(24);
output(2, 201) <= input(25);
output(2, 202) <= input(26);
output(2, 203) <= input(27);
output(2, 204) <= input(28);
output(2, 205) <= input(29);
output(2, 206) <= input(30);
output(2, 207) <= input(31);
output(2, 208) <= input(16);
output(2, 209) <= input(17);
output(2, 210) <= input(18);
output(2, 211) <= input(19);
output(2, 212) <= input(20);
output(2, 213) <= input(21);
output(2, 214) <= input(22);
output(2, 215) <= input(23);
output(2, 216) <= input(24);
output(2, 217) <= input(25);
output(2, 218) <= input(26);
output(2, 219) <= input(27);
output(2, 220) <= input(28);
output(2, 221) <= input(29);
output(2, 222) <= input(30);
output(2, 223) <= input(31);
output(2, 224) <= input(16);
output(2, 225) <= input(17);
output(2, 226) <= input(18);
output(2, 227) <= input(19);
output(2, 228) <= input(20);
output(2, 229) <= input(21);
output(2, 230) <= input(22);
output(2, 231) <= input(23);
output(2, 232) <= input(24);
output(2, 233) <= input(25);
output(2, 234) <= input(26);
output(2, 235) <= input(27);
output(2, 236) <= input(28);
output(2, 237) <= input(29);
output(2, 238) <= input(30);
output(2, 239) <= input(31);
output(2, 240) <= input(1);
output(2, 241) <= input(2);
output(2, 242) <= input(3);
output(2, 243) <= input(4);
output(2, 244) <= input(5);
output(2, 245) <= input(6);
output(2, 246) <= input(7);
output(2, 247) <= input(8);
output(2, 248) <= input(9);
output(2, 249) <= input(10);
output(2, 250) <= input(11);
output(2, 251) <= input(12);
output(2, 252) <= input(13);
output(2, 253) <= input(14);
output(2, 254) <= input(15);
output(2, 255) <= input(32);
output(3, 0) <= input(0);
output(3, 1) <= input(1);
output(3, 2) <= input(2);
output(3, 3) <= input(3);
output(3, 4) <= input(4);
output(3, 5) <= input(5);
output(3, 6) <= input(6);
output(3, 7) <= input(7);
output(3, 8) <= input(8);
output(3, 9) <= input(9);
output(3, 10) <= input(10);
output(3, 11) <= input(11);
output(3, 12) <= input(12);
output(3, 13) <= input(13);
output(3, 14) <= input(14);
output(3, 15) <= input(15);
output(3, 16) <= input(0);
output(3, 17) <= input(1);
output(3, 18) <= input(2);
output(3, 19) <= input(3);
output(3, 20) <= input(4);
output(3, 21) <= input(5);
output(3, 22) <= input(6);
output(3, 23) <= input(7);
output(3, 24) <= input(8);
output(3, 25) <= input(9);
output(3, 26) <= input(10);
output(3, 27) <= input(11);
output(3, 28) <= input(12);
output(3, 29) <= input(13);
output(3, 30) <= input(14);
output(3, 31) <= input(15);
output(3, 32) <= input(0);
output(3, 33) <= input(1);
output(3, 34) <= input(2);
output(3, 35) <= input(3);
output(3, 36) <= input(4);
output(3, 37) <= input(5);
output(3, 38) <= input(6);
output(3, 39) <= input(7);
output(3, 40) <= input(8);
output(3, 41) <= input(9);
output(3, 42) <= input(10);
output(3, 43) <= input(11);
output(3, 44) <= input(12);
output(3, 45) <= input(13);
output(3, 46) <= input(14);
output(3, 47) <= input(15);
output(3, 48) <= input(0);
output(3, 49) <= input(1);
output(3, 50) <= input(2);
output(3, 51) <= input(3);
output(3, 52) <= input(4);
output(3, 53) <= input(5);
output(3, 54) <= input(6);
output(3, 55) <= input(7);
output(3, 56) <= input(8);
output(3, 57) <= input(9);
output(3, 58) <= input(10);
output(3, 59) <= input(11);
output(3, 60) <= input(12);
output(3, 61) <= input(13);
output(3, 62) <= input(14);
output(3, 63) <= input(15);
output(3, 64) <= input(0);
output(3, 65) <= input(1);
output(3, 66) <= input(2);
output(3, 67) <= input(3);
output(3, 68) <= input(4);
output(3, 69) <= input(5);
output(3, 70) <= input(6);
output(3, 71) <= input(7);
output(3, 72) <= input(8);
output(3, 73) <= input(9);
output(3, 74) <= input(10);
output(3, 75) <= input(11);
output(3, 76) <= input(12);
output(3, 77) <= input(13);
output(3, 78) <= input(14);
output(3, 79) <= input(15);
output(3, 80) <= input(0);
output(3, 81) <= input(1);
output(3, 82) <= input(2);
output(3, 83) <= input(3);
output(3, 84) <= input(4);
output(3, 85) <= input(5);
output(3, 86) <= input(6);
output(3, 87) <= input(7);
output(3, 88) <= input(8);
output(3, 89) <= input(9);
output(3, 90) <= input(10);
output(3, 91) <= input(11);
output(3, 92) <= input(12);
output(3, 93) <= input(13);
output(3, 94) <= input(14);
output(3, 95) <= input(15);
output(3, 96) <= input(0);
output(3, 97) <= input(1);
output(3, 98) <= input(2);
output(3, 99) <= input(3);
output(3, 100) <= input(4);
output(3, 101) <= input(5);
output(3, 102) <= input(6);
output(3, 103) <= input(7);
output(3, 104) <= input(8);
output(3, 105) <= input(9);
output(3, 106) <= input(10);
output(3, 107) <= input(11);
output(3, 108) <= input(12);
output(3, 109) <= input(13);
output(3, 110) <= input(14);
output(3, 111) <= input(15);
output(3, 112) <= input(0);
output(3, 113) <= input(1);
output(3, 114) <= input(2);
output(3, 115) <= input(3);
output(3, 116) <= input(4);
output(3, 117) <= input(5);
output(3, 118) <= input(6);
output(3, 119) <= input(7);
output(3, 120) <= input(8);
output(3, 121) <= input(9);
output(3, 122) <= input(10);
output(3, 123) <= input(11);
output(3, 124) <= input(12);
output(3, 125) <= input(13);
output(3, 126) <= input(14);
output(3, 127) <= input(15);
output(3, 128) <= input(0);
output(3, 129) <= input(1);
output(3, 130) <= input(2);
output(3, 131) <= input(3);
output(3, 132) <= input(4);
output(3, 133) <= input(5);
output(3, 134) <= input(6);
output(3, 135) <= input(7);
output(3, 136) <= input(8);
output(3, 137) <= input(9);
output(3, 138) <= input(10);
output(3, 139) <= input(11);
output(3, 140) <= input(12);
output(3, 141) <= input(13);
output(3, 142) <= input(14);
output(3, 143) <= input(15);
output(3, 144) <= input(0);
output(3, 145) <= input(1);
output(3, 146) <= input(2);
output(3, 147) <= input(3);
output(3, 148) <= input(4);
output(3, 149) <= input(5);
output(3, 150) <= input(6);
output(3, 151) <= input(7);
output(3, 152) <= input(8);
output(3, 153) <= input(9);
output(3, 154) <= input(10);
output(3, 155) <= input(11);
output(3, 156) <= input(12);
output(3, 157) <= input(13);
output(3, 158) <= input(14);
output(3, 159) <= input(15);
output(3, 160) <= input(0);
output(3, 161) <= input(1);
output(3, 162) <= input(2);
output(3, 163) <= input(3);
output(3, 164) <= input(4);
output(3, 165) <= input(5);
output(3, 166) <= input(6);
output(3, 167) <= input(7);
output(3, 168) <= input(8);
output(3, 169) <= input(9);
output(3, 170) <= input(10);
output(3, 171) <= input(11);
output(3, 172) <= input(12);
output(3, 173) <= input(13);
output(3, 174) <= input(14);
output(3, 175) <= input(15);
output(3, 176) <= input(0);
output(3, 177) <= input(1);
output(3, 178) <= input(2);
output(3, 179) <= input(3);
output(3, 180) <= input(4);
output(3, 181) <= input(5);
output(3, 182) <= input(6);
output(3, 183) <= input(7);
output(3, 184) <= input(8);
output(3, 185) <= input(9);
output(3, 186) <= input(10);
output(3, 187) <= input(11);
output(3, 188) <= input(12);
output(3, 189) <= input(13);
output(3, 190) <= input(14);
output(3, 191) <= input(15);
output(3, 192) <= input(0);
output(3, 193) <= input(1);
output(3, 194) <= input(2);
output(3, 195) <= input(3);
output(3, 196) <= input(4);
output(3, 197) <= input(5);
output(3, 198) <= input(6);
output(3, 199) <= input(7);
output(3, 200) <= input(8);
output(3, 201) <= input(9);
output(3, 202) <= input(10);
output(3, 203) <= input(11);
output(3, 204) <= input(12);
output(3, 205) <= input(13);
output(3, 206) <= input(14);
output(3, 207) <= input(15);
output(3, 208) <= input(0);
output(3, 209) <= input(1);
output(3, 210) <= input(2);
output(3, 211) <= input(3);
output(3, 212) <= input(4);
output(3, 213) <= input(5);
output(3, 214) <= input(6);
output(3, 215) <= input(7);
output(3, 216) <= input(8);
output(3, 217) <= input(9);
output(3, 218) <= input(10);
output(3, 219) <= input(11);
output(3, 220) <= input(12);
output(3, 221) <= input(13);
output(3, 222) <= input(14);
output(3, 223) <= input(15);
output(3, 224) <= input(0);
output(3, 225) <= input(1);
output(3, 226) <= input(2);
output(3, 227) <= input(3);
output(3, 228) <= input(4);
output(3, 229) <= input(5);
output(3, 230) <= input(6);
output(3, 231) <= input(7);
output(3, 232) <= input(8);
output(3, 233) <= input(9);
output(3, 234) <= input(10);
output(3, 235) <= input(11);
output(3, 236) <= input(12);
output(3, 237) <= input(13);
output(3, 238) <= input(14);
output(3, 239) <= input(15);
output(3, 240) <= input(16);
output(3, 241) <= input(17);
output(3, 242) <= input(18);
output(3, 243) <= input(19);
output(3, 244) <= input(20);
output(3, 245) <= input(21);
output(3, 246) <= input(22);
output(3, 247) <= input(23);
output(3, 248) <= input(24);
output(3, 249) <= input(25);
output(3, 250) <= input(26);
output(3, 251) <= input(27);
output(3, 252) <= input(28);
output(3, 253) <= input(29);
output(3, 254) <= input(30);
output(3, 255) <= input(31);
output(4, 0) <= input(0);
output(4, 1) <= input(1);
output(4, 2) <= input(2);
output(4, 3) <= input(3);
output(4, 4) <= input(4);
output(4, 5) <= input(5);
output(4, 6) <= input(6);
output(4, 7) <= input(7);
output(4, 8) <= input(8);
output(4, 9) <= input(9);
output(4, 10) <= input(10);
output(4, 11) <= input(11);
output(4, 12) <= input(12);
output(4, 13) <= input(13);
output(4, 14) <= input(14);
output(4, 15) <= input(15);
output(4, 16) <= input(0);
output(4, 17) <= input(1);
output(4, 18) <= input(2);
output(4, 19) <= input(3);
output(4, 20) <= input(4);
output(4, 21) <= input(5);
output(4, 22) <= input(6);
output(4, 23) <= input(7);
output(4, 24) <= input(8);
output(4, 25) <= input(9);
output(4, 26) <= input(10);
output(4, 27) <= input(11);
output(4, 28) <= input(12);
output(4, 29) <= input(13);
output(4, 30) <= input(14);
output(4, 31) <= input(15);
output(4, 32) <= input(0);
output(4, 33) <= input(1);
output(4, 34) <= input(2);
output(4, 35) <= input(3);
output(4, 36) <= input(4);
output(4, 37) <= input(5);
output(4, 38) <= input(6);
output(4, 39) <= input(7);
output(4, 40) <= input(8);
output(4, 41) <= input(9);
output(4, 42) <= input(10);
output(4, 43) <= input(11);
output(4, 44) <= input(12);
output(4, 45) <= input(13);
output(4, 46) <= input(14);
output(4, 47) <= input(15);
output(4, 48) <= input(0);
output(4, 49) <= input(1);
output(4, 50) <= input(2);
output(4, 51) <= input(3);
output(4, 52) <= input(4);
output(4, 53) <= input(5);
output(4, 54) <= input(6);
output(4, 55) <= input(7);
output(4, 56) <= input(8);
output(4, 57) <= input(9);
output(4, 58) <= input(10);
output(4, 59) <= input(11);
output(4, 60) <= input(12);
output(4, 61) <= input(13);
output(4, 62) <= input(14);
output(4, 63) <= input(15);
output(4, 64) <= input(0);
output(4, 65) <= input(1);
output(4, 66) <= input(2);
output(4, 67) <= input(3);
output(4, 68) <= input(4);
output(4, 69) <= input(5);
output(4, 70) <= input(6);
output(4, 71) <= input(7);
output(4, 72) <= input(8);
output(4, 73) <= input(9);
output(4, 74) <= input(10);
output(4, 75) <= input(11);
output(4, 76) <= input(12);
output(4, 77) <= input(13);
output(4, 78) <= input(14);
output(4, 79) <= input(15);
output(4, 80) <= input(0);
output(4, 81) <= input(1);
output(4, 82) <= input(2);
output(4, 83) <= input(3);
output(4, 84) <= input(4);
output(4, 85) <= input(5);
output(4, 86) <= input(6);
output(4, 87) <= input(7);
output(4, 88) <= input(8);
output(4, 89) <= input(9);
output(4, 90) <= input(10);
output(4, 91) <= input(11);
output(4, 92) <= input(12);
output(4, 93) <= input(13);
output(4, 94) <= input(14);
output(4, 95) <= input(15);
output(4, 96) <= input(0);
output(4, 97) <= input(1);
output(4, 98) <= input(2);
output(4, 99) <= input(3);
output(4, 100) <= input(4);
output(4, 101) <= input(5);
output(4, 102) <= input(6);
output(4, 103) <= input(7);
output(4, 104) <= input(8);
output(4, 105) <= input(9);
output(4, 106) <= input(10);
output(4, 107) <= input(11);
output(4, 108) <= input(12);
output(4, 109) <= input(13);
output(4, 110) <= input(14);
output(4, 111) <= input(15);
output(4, 112) <= input(0);
output(4, 113) <= input(1);
output(4, 114) <= input(2);
output(4, 115) <= input(3);
output(4, 116) <= input(4);
output(4, 117) <= input(5);
output(4, 118) <= input(6);
output(4, 119) <= input(7);
output(4, 120) <= input(8);
output(4, 121) <= input(9);
output(4, 122) <= input(10);
output(4, 123) <= input(11);
output(4, 124) <= input(12);
output(4, 125) <= input(13);
output(4, 126) <= input(14);
output(4, 127) <= input(15);
output(4, 128) <= input(0);
output(4, 129) <= input(1);
output(4, 130) <= input(2);
output(4, 131) <= input(3);
output(4, 132) <= input(4);
output(4, 133) <= input(5);
output(4, 134) <= input(6);
output(4, 135) <= input(7);
output(4, 136) <= input(8);
output(4, 137) <= input(9);
output(4, 138) <= input(10);
output(4, 139) <= input(11);
output(4, 140) <= input(12);
output(4, 141) <= input(13);
output(4, 142) <= input(14);
output(4, 143) <= input(15);
output(4, 144) <= input(0);
output(4, 145) <= input(1);
output(4, 146) <= input(2);
output(4, 147) <= input(3);
output(4, 148) <= input(4);
output(4, 149) <= input(5);
output(4, 150) <= input(6);
output(4, 151) <= input(7);
output(4, 152) <= input(8);
output(4, 153) <= input(9);
output(4, 154) <= input(10);
output(4, 155) <= input(11);
output(4, 156) <= input(12);
output(4, 157) <= input(13);
output(4, 158) <= input(14);
output(4, 159) <= input(15);
output(4, 160) <= input(0);
output(4, 161) <= input(1);
output(4, 162) <= input(2);
output(4, 163) <= input(3);
output(4, 164) <= input(4);
output(4, 165) <= input(5);
output(4, 166) <= input(6);
output(4, 167) <= input(7);
output(4, 168) <= input(8);
output(4, 169) <= input(9);
output(4, 170) <= input(10);
output(4, 171) <= input(11);
output(4, 172) <= input(12);
output(4, 173) <= input(13);
output(4, 174) <= input(14);
output(4, 175) <= input(15);
output(4, 176) <= input(0);
output(4, 177) <= input(1);
output(4, 178) <= input(2);
output(4, 179) <= input(3);
output(4, 180) <= input(4);
output(4, 181) <= input(5);
output(4, 182) <= input(6);
output(4, 183) <= input(7);
output(4, 184) <= input(8);
output(4, 185) <= input(9);
output(4, 186) <= input(10);
output(4, 187) <= input(11);
output(4, 188) <= input(12);
output(4, 189) <= input(13);
output(4, 190) <= input(14);
output(4, 191) <= input(15);
output(4, 192) <= input(0);
output(4, 193) <= input(1);
output(4, 194) <= input(2);
output(4, 195) <= input(3);
output(4, 196) <= input(4);
output(4, 197) <= input(5);
output(4, 198) <= input(6);
output(4, 199) <= input(7);
output(4, 200) <= input(8);
output(4, 201) <= input(9);
output(4, 202) <= input(10);
output(4, 203) <= input(11);
output(4, 204) <= input(12);
output(4, 205) <= input(13);
output(4, 206) <= input(14);
output(4, 207) <= input(15);
output(4, 208) <= input(0);
output(4, 209) <= input(1);
output(4, 210) <= input(2);
output(4, 211) <= input(3);
output(4, 212) <= input(4);
output(4, 213) <= input(5);
output(4, 214) <= input(6);
output(4, 215) <= input(7);
output(4, 216) <= input(8);
output(4, 217) <= input(9);
output(4, 218) <= input(10);
output(4, 219) <= input(11);
output(4, 220) <= input(12);
output(4, 221) <= input(13);
output(4, 222) <= input(14);
output(4, 223) <= input(15);
output(4, 224) <= input(0);
output(4, 225) <= input(1);
output(4, 226) <= input(2);
output(4, 227) <= input(3);
output(4, 228) <= input(4);
output(4, 229) <= input(5);
output(4, 230) <= input(6);
output(4, 231) <= input(7);
output(4, 232) <= input(8);
output(4, 233) <= input(9);
output(4, 234) <= input(10);
output(4, 235) <= input(11);
output(4, 236) <= input(12);
output(4, 237) <= input(13);
output(4, 238) <= input(14);
output(4, 239) <= input(15);
output(4, 240) <= input(0);
output(4, 241) <= input(1);
output(4, 242) <= input(2);
output(4, 243) <= input(3);
output(4, 244) <= input(4);
output(4, 245) <= input(5);
output(4, 246) <= input(6);
output(4, 247) <= input(7);
output(4, 248) <= input(8);
output(4, 249) <= input(9);
output(4, 250) <= input(10);
output(4, 251) <= input(11);
output(4, 252) <= input(12);
output(4, 253) <= input(13);
output(4, 254) <= input(14);
output(4, 255) <= input(15);
output(5, 0) <= input(35);
output(5, 1) <= input(16);
output(5, 2) <= input(17);
output(5, 3) <= input(18);
output(5, 4) <= input(19);
output(5, 5) <= input(20);
output(5, 6) <= input(21);
output(5, 7) <= input(22);
output(5, 8) <= input(23);
output(5, 9) <= input(24);
output(5, 10) <= input(25);
output(5, 11) <= input(26);
output(5, 12) <= input(27);
output(5, 13) <= input(28);
output(5, 14) <= input(29);
output(5, 15) <= input(30);
output(5, 16) <= input(35);
output(5, 17) <= input(16);
output(5, 18) <= input(17);
output(5, 19) <= input(18);
output(5, 20) <= input(19);
output(5, 21) <= input(20);
output(5, 22) <= input(21);
output(5, 23) <= input(22);
output(5, 24) <= input(23);
output(5, 25) <= input(24);
output(5, 26) <= input(25);
output(5, 27) <= input(26);
output(5, 28) <= input(27);
output(5, 29) <= input(28);
output(5, 30) <= input(29);
output(5, 31) <= input(30);
output(5, 32) <= input(35);
output(5, 33) <= input(16);
output(5, 34) <= input(17);
output(5, 35) <= input(18);
output(5, 36) <= input(19);
output(5, 37) <= input(20);
output(5, 38) <= input(21);
output(5, 39) <= input(22);
output(5, 40) <= input(23);
output(5, 41) <= input(24);
output(5, 42) <= input(25);
output(5, 43) <= input(26);
output(5, 44) <= input(27);
output(5, 45) <= input(28);
output(5, 46) <= input(29);
output(5, 47) <= input(30);
output(5, 48) <= input(35);
output(5, 49) <= input(16);
output(5, 50) <= input(17);
output(5, 51) <= input(18);
output(5, 52) <= input(19);
output(5, 53) <= input(20);
output(5, 54) <= input(21);
output(5, 55) <= input(22);
output(5, 56) <= input(23);
output(5, 57) <= input(24);
output(5, 58) <= input(25);
output(5, 59) <= input(26);
output(5, 60) <= input(27);
output(5, 61) <= input(28);
output(5, 62) <= input(29);
output(5, 63) <= input(30);
output(5, 64) <= input(35);
output(5, 65) <= input(16);
output(5, 66) <= input(17);
output(5, 67) <= input(18);
output(5, 68) <= input(19);
output(5, 69) <= input(20);
output(5, 70) <= input(21);
output(5, 71) <= input(22);
output(5, 72) <= input(23);
output(5, 73) <= input(24);
output(5, 74) <= input(25);
output(5, 75) <= input(26);
output(5, 76) <= input(27);
output(5, 77) <= input(28);
output(5, 78) <= input(29);
output(5, 79) <= input(30);
output(5, 80) <= input(35);
output(5, 81) <= input(16);
output(5, 82) <= input(17);
output(5, 83) <= input(18);
output(5, 84) <= input(19);
output(5, 85) <= input(20);
output(5, 86) <= input(21);
output(5, 87) <= input(22);
output(5, 88) <= input(23);
output(5, 89) <= input(24);
output(5, 90) <= input(25);
output(5, 91) <= input(26);
output(5, 92) <= input(27);
output(5, 93) <= input(28);
output(5, 94) <= input(29);
output(5, 95) <= input(30);
output(5, 96) <= input(35);
output(5, 97) <= input(16);
output(5, 98) <= input(17);
output(5, 99) <= input(18);
output(5, 100) <= input(19);
output(5, 101) <= input(20);
output(5, 102) <= input(21);
output(5, 103) <= input(22);
output(5, 104) <= input(23);
output(5, 105) <= input(24);
output(5, 106) <= input(25);
output(5, 107) <= input(26);
output(5, 108) <= input(27);
output(5, 109) <= input(28);
output(5, 110) <= input(29);
output(5, 111) <= input(30);
output(5, 112) <= input(35);
output(5, 113) <= input(16);
output(5, 114) <= input(17);
output(5, 115) <= input(18);
output(5, 116) <= input(19);
output(5, 117) <= input(20);
output(5, 118) <= input(21);
output(5, 119) <= input(22);
output(5, 120) <= input(23);
output(5, 121) <= input(24);
output(5, 122) <= input(25);
output(5, 123) <= input(26);
output(5, 124) <= input(27);
output(5, 125) <= input(28);
output(5, 126) <= input(29);
output(5, 127) <= input(30);
output(5, 128) <= input(35);
output(5, 129) <= input(16);
output(5, 130) <= input(17);
output(5, 131) <= input(18);
output(5, 132) <= input(19);
output(5, 133) <= input(20);
output(5, 134) <= input(21);
output(5, 135) <= input(22);
output(5, 136) <= input(23);
output(5, 137) <= input(24);
output(5, 138) <= input(25);
output(5, 139) <= input(26);
output(5, 140) <= input(27);
output(5, 141) <= input(28);
output(5, 142) <= input(29);
output(5, 143) <= input(30);
output(5, 144) <= input(35);
output(5, 145) <= input(16);
output(5, 146) <= input(17);
output(5, 147) <= input(18);
output(5, 148) <= input(19);
output(5, 149) <= input(20);
output(5, 150) <= input(21);
output(5, 151) <= input(22);
output(5, 152) <= input(23);
output(5, 153) <= input(24);
output(5, 154) <= input(25);
output(5, 155) <= input(26);
output(5, 156) <= input(27);
output(5, 157) <= input(28);
output(5, 158) <= input(29);
output(5, 159) <= input(30);
output(5, 160) <= input(35);
output(5, 161) <= input(16);
output(5, 162) <= input(17);
output(5, 163) <= input(18);
output(5, 164) <= input(19);
output(5, 165) <= input(20);
output(5, 166) <= input(21);
output(5, 167) <= input(22);
output(5, 168) <= input(23);
output(5, 169) <= input(24);
output(5, 170) <= input(25);
output(5, 171) <= input(26);
output(5, 172) <= input(27);
output(5, 173) <= input(28);
output(5, 174) <= input(29);
output(5, 175) <= input(30);
output(5, 176) <= input(35);
output(5, 177) <= input(16);
output(5, 178) <= input(17);
output(5, 179) <= input(18);
output(5, 180) <= input(19);
output(5, 181) <= input(20);
output(5, 182) <= input(21);
output(5, 183) <= input(22);
output(5, 184) <= input(23);
output(5, 185) <= input(24);
output(5, 186) <= input(25);
output(5, 187) <= input(26);
output(5, 188) <= input(27);
output(5, 189) <= input(28);
output(5, 190) <= input(29);
output(5, 191) <= input(30);
output(5, 192) <= input(35);
output(5, 193) <= input(16);
output(5, 194) <= input(17);
output(5, 195) <= input(18);
output(5, 196) <= input(19);
output(5, 197) <= input(20);
output(5, 198) <= input(21);
output(5, 199) <= input(22);
output(5, 200) <= input(23);
output(5, 201) <= input(24);
output(5, 202) <= input(25);
output(5, 203) <= input(26);
output(5, 204) <= input(27);
output(5, 205) <= input(28);
output(5, 206) <= input(29);
output(5, 207) <= input(30);
output(5, 208) <= input(35);
output(5, 209) <= input(16);
output(5, 210) <= input(17);
output(5, 211) <= input(18);
output(5, 212) <= input(19);
output(5, 213) <= input(20);
output(5, 214) <= input(21);
output(5, 215) <= input(22);
output(5, 216) <= input(23);
output(5, 217) <= input(24);
output(5, 218) <= input(25);
output(5, 219) <= input(26);
output(5, 220) <= input(27);
output(5, 221) <= input(28);
output(5, 222) <= input(29);
output(5, 223) <= input(30);
output(5, 224) <= input(35);
output(5, 225) <= input(16);
output(5, 226) <= input(17);
output(5, 227) <= input(18);
output(5, 228) <= input(19);
output(5, 229) <= input(20);
output(5, 230) <= input(21);
output(5, 231) <= input(22);
output(5, 232) <= input(23);
output(5, 233) <= input(24);
output(5, 234) <= input(25);
output(5, 235) <= input(26);
output(5, 236) <= input(27);
output(5, 237) <= input(28);
output(5, 238) <= input(29);
output(5, 239) <= input(30);
output(5, 240) <= input(35);
output(5, 241) <= input(16);
output(5, 242) <= input(17);
output(5, 243) <= input(18);
output(5, 244) <= input(19);
output(5, 245) <= input(20);
output(5, 246) <= input(21);
output(5, 247) <= input(22);
output(5, 248) <= input(23);
output(5, 249) <= input(24);
output(5, 250) <= input(25);
output(5, 251) <= input(26);
output(5, 252) <= input(27);
output(5, 253) <= input(28);
output(5, 254) <= input(29);
output(5, 255) <= input(30);
output(6, 0) <= input(35);
output(6, 1) <= input(16);
output(6, 2) <= input(17);
output(6, 3) <= input(18);
output(6, 4) <= input(19);
output(6, 5) <= input(20);
output(6, 6) <= input(21);
output(6, 7) <= input(22);
output(6, 8) <= input(23);
output(6, 9) <= input(24);
output(6, 10) <= input(25);
output(6, 11) <= input(26);
output(6, 12) <= input(27);
output(6, 13) <= input(28);
output(6, 14) <= input(29);
output(6, 15) <= input(30);
output(6, 16) <= input(35);
output(6, 17) <= input(16);
output(6, 18) <= input(17);
output(6, 19) <= input(18);
output(6, 20) <= input(19);
output(6, 21) <= input(20);
output(6, 22) <= input(21);
output(6, 23) <= input(22);
output(6, 24) <= input(23);
output(6, 25) <= input(24);
output(6, 26) <= input(25);
output(6, 27) <= input(26);
output(6, 28) <= input(27);
output(6, 29) <= input(28);
output(6, 30) <= input(29);
output(6, 31) <= input(30);
output(6, 32) <= input(35);
output(6, 33) <= input(16);
output(6, 34) <= input(17);
output(6, 35) <= input(18);
output(6, 36) <= input(19);
output(6, 37) <= input(20);
output(6, 38) <= input(21);
output(6, 39) <= input(22);
output(6, 40) <= input(23);
output(6, 41) <= input(24);
output(6, 42) <= input(25);
output(6, 43) <= input(26);
output(6, 44) <= input(27);
output(6, 45) <= input(28);
output(6, 46) <= input(29);
output(6, 47) <= input(30);
output(6, 48) <= input(35);
output(6, 49) <= input(16);
output(6, 50) <= input(17);
output(6, 51) <= input(18);
output(6, 52) <= input(19);
output(6, 53) <= input(20);
output(6, 54) <= input(21);
output(6, 55) <= input(22);
output(6, 56) <= input(23);
output(6, 57) <= input(24);
output(6, 58) <= input(25);
output(6, 59) <= input(26);
output(6, 60) <= input(27);
output(6, 61) <= input(28);
output(6, 62) <= input(29);
output(6, 63) <= input(30);
output(6, 64) <= input(35);
output(6, 65) <= input(16);
output(6, 66) <= input(17);
output(6, 67) <= input(18);
output(6, 68) <= input(19);
output(6, 69) <= input(20);
output(6, 70) <= input(21);
output(6, 71) <= input(22);
output(6, 72) <= input(23);
output(6, 73) <= input(24);
output(6, 74) <= input(25);
output(6, 75) <= input(26);
output(6, 76) <= input(27);
output(6, 77) <= input(28);
output(6, 78) <= input(29);
output(6, 79) <= input(30);
output(6, 80) <= input(35);
output(6, 81) <= input(16);
output(6, 82) <= input(17);
output(6, 83) <= input(18);
output(6, 84) <= input(19);
output(6, 85) <= input(20);
output(6, 86) <= input(21);
output(6, 87) <= input(22);
output(6, 88) <= input(23);
output(6, 89) <= input(24);
output(6, 90) <= input(25);
output(6, 91) <= input(26);
output(6, 92) <= input(27);
output(6, 93) <= input(28);
output(6, 94) <= input(29);
output(6, 95) <= input(30);
output(6, 96) <= input(35);
output(6, 97) <= input(16);
output(6, 98) <= input(17);
output(6, 99) <= input(18);
output(6, 100) <= input(19);
output(6, 101) <= input(20);
output(6, 102) <= input(21);
output(6, 103) <= input(22);
output(6, 104) <= input(23);
output(6, 105) <= input(24);
output(6, 106) <= input(25);
output(6, 107) <= input(26);
output(6, 108) <= input(27);
output(6, 109) <= input(28);
output(6, 110) <= input(29);
output(6, 111) <= input(30);
output(6, 112) <= input(35);
output(6, 113) <= input(16);
output(6, 114) <= input(17);
output(6, 115) <= input(18);
output(6, 116) <= input(19);
output(6, 117) <= input(20);
output(6, 118) <= input(21);
output(6, 119) <= input(22);
output(6, 120) <= input(23);
output(6, 121) <= input(24);
output(6, 122) <= input(25);
output(6, 123) <= input(26);
output(6, 124) <= input(27);
output(6, 125) <= input(28);
output(6, 126) <= input(29);
output(6, 127) <= input(30);
output(6, 128) <= input(36);
output(6, 129) <= input(0);
output(6, 130) <= input(1);
output(6, 131) <= input(2);
output(6, 132) <= input(3);
output(6, 133) <= input(4);
output(6, 134) <= input(5);
output(6, 135) <= input(6);
output(6, 136) <= input(7);
output(6, 137) <= input(8);
output(6, 138) <= input(9);
output(6, 139) <= input(10);
output(6, 140) <= input(11);
output(6, 141) <= input(12);
output(6, 142) <= input(13);
output(6, 143) <= input(14);
output(6, 144) <= input(36);
output(6, 145) <= input(0);
output(6, 146) <= input(1);
output(6, 147) <= input(2);
output(6, 148) <= input(3);
output(6, 149) <= input(4);
output(6, 150) <= input(5);
output(6, 151) <= input(6);
output(6, 152) <= input(7);
output(6, 153) <= input(8);
output(6, 154) <= input(9);
output(6, 155) <= input(10);
output(6, 156) <= input(11);
output(6, 157) <= input(12);
output(6, 158) <= input(13);
output(6, 159) <= input(14);
output(6, 160) <= input(36);
output(6, 161) <= input(0);
output(6, 162) <= input(1);
output(6, 163) <= input(2);
output(6, 164) <= input(3);
output(6, 165) <= input(4);
output(6, 166) <= input(5);
output(6, 167) <= input(6);
output(6, 168) <= input(7);
output(6, 169) <= input(8);
output(6, 170) <= input(9);
output(6, 171) <= input(10);
output(6, 172) <= input(11);
output(6, 173) <= input(12);
output(6, 174) <= input(13);
output(6, 175) <= input(14);
output(6, 176) <= input(36);
output(6, 177) <= input(0);
output(6, 178) <= input(1);
output(6, 179) <= input(2);
output(6, 180) <= input(3);
output(6, 181) <= input(4);
output(6, 182) <= input(5);
output(6, 183) <= input(6);
output(6, 184) <= input(7);
output(6, 185) <= input(8);
output(6, 186) <= input(9);
output(6, 187) <= input(10);
output(6, 188) <= input(11);
output(6, 189) <= input(12);
output(6, 190) <= input(13);
output(6, 191) <= input(14);
output(6, 192) <= input(36);
output(6, 193) <= input(0);
output(6, 194) <= input(1);
output(6, 195) <= input(2);
output(6, 196) <= input(3);
output(6, 197) <= input(4);
output(6, 198) <= input(5);
output(6, 199) <= input(6);
output(6, 200) <= input(7);
output(6, 201) <= input(8);
output(6, 202) <= input(9);
output(6, 203) <= input(10);
output(6, 204) <= input(11);
output(6, 205) <= input(12);
output(6, 206) <= input(13);
output(6, 207) <= input(14);
output(6, 208) <= input(36);
output(6, 209) <= input(0);
output(6, 210) <= input(1);
output(6, 211) <= input(2);
output(6, 212) <= input(3);
output(6, 213) <= input(4);
output(6, 214) <= input(5);
output(6, 215) <= input(6);
output(6, 216) <= input(7);
output(6, 217) <= input(8);
output(6, 218) <= input(9);
output(6, 219) <= input(10);
output(6, 220) <= input(11);
output(6, 221) <= input(12);
output(6, 222) <= input(13);
output(6, 223) <= input(14);
output(6, 224) <= input(36);
output(6, 225) <= input(0);
output(6, 226) <= input(1);
output(6, 227) <= input(2);
output(6, 228) <= input(3);
output(6, 229) <= input(4);
output(6, 230) <= input(5);
output(6, 231) <= input(6);
output(6, 232) <= input(7);
output(6, 233) <= input(8);
output(6, 234) <= input(9);
output(6, 235) <= input(10);
output(6, 236) <= input(11);
output(6, 237) <= input(12);
output(6, 238) <= input(13);
output(6, 239) <= input(14);
output(6, 240) <= input(36);
output(6, 241) <= input(0);
output(6, 242) <= input(1);
output(6, 243) <= input(2);
output(6, 244) <= input(3);
output(6, 245) <= input(4);
output(6, 246) <= input(5);
output(6, 247) <= input(6);
output(6, 248) <= input(7);
output(6, 249) <= input(8);
output(6, 250) <= input(9);
output(6, 251) <= input(10);
output(6, 252) <= input(11);
output(6, 253) <= input(12);
output(6, 254) <= input(13);
output(6, 255) <= input(14);
output(7, 0) <= input(35);
output(7, 1) <= input(16);
output(7, 2) <= input(17);
output(7, 3) <= input(18);
output(7, 4) <= input(19);
output(7, 5) <= input(20);
output(7, 6) <= input(21);
output(7, 7) <= input(22);
output(7, 8) <= input(23);
output(7, 9) <= input(24);
output(7, 10) <= input(25);
output(7, 11) <= input(26);
output(7, 12) <= input(27);
output(7, 13) <= input(28);
output(7, 14) <= input(29);
output(7, 15) <= input(30);
output(7, 16) <= input(35);
output(7, 17) <= input(16);
output(7, 18) <= input(17);
output(7, 19) <= input(18);
output(7, 20) <= input(19);
output(7, 21) <= input(20);
output(7, 22) <= input(21);
output(7, 23) <= input(22);
output(7, 24) <= input(23);
output(7, 25) <= input(24);
output(7, 26) <= input(25);
output(7, 27) <= input(26);
output(7, 28) <= input(27);
output(7, 29) <= input(28);
output(7, 30) <= input(29);
output(7, 31) <= input(30);
output(7, 32) <= input(35);
output(7, 33) <= input(16);
output(7, 34) <= input(17);
output(7, 35) <= input(18);
output(7, 36) <= input(19);
output(7, 37) <= input(20);
output(7, 38) <= input(21);
output(7, 39) <= input(22);
output(7, 40) <= input(23);
output(7, 41) <= input(24);
output(7, 42) <= input(25);
output(7, 43) <= input(26);
output(7, 44) <= input(27);
output(7, 45) <= input(28);
output(7, 46) <= input(29);
output(7, 47) <= input(30);
output(7, 48) <= input(35);
output(7, 49) <= input(16);
output(7, 50) <= input(17);
output(7, 51) <= input(18);
output(7, 52) <= input(19);
output(7, 53) <= input(20);
output(7, 54) <= input(21);
output(7, 55) <= input(22);
output(7, 56) <= input(23);
output(7, 57) <= input(24);
output(7, 58) <= input(25);
output(7, 59) <= input(26);
output(7, 60) <= input(27);
output(7, 61) <= input(28);
output(7, 62) <= input(29);
output(7, 63) <= input(30);
output(7, 64) <= input(35);
output(7, 65) <= input(16);
output(7, 66) <= input(17);
output(7, 67) <= input(18);
output(7, 68) <= input(19);
output(7, 69) <= input(20);
output(7, 70) <= input(21);
output(7, 71) <= input(22);
output(7, 72) <= input(23);
output(7, 73) <= input(24);
output(7, 74) <= input(25);
output(7, 75) <= input(26);
output(7, 76) <= input(27);
output(7, 77) <= input(28);
output(7, 78) <= input(29);
output(7, 79) <= input(30);
output(7, 80) <= input(36);
output(7, 81) <= input(0);
output(7, 82) <= input(1);
output(7, 83) <= input(2);
output(7, 84) <= input(3);
output(7, 85) <= input(4);
output(7, 86) <= input(5);
output(7, 87) <= input(6);
output(7, 88) <= input(7);
output(7, 89) <= input(8);
output(7, 90) <= input(9);
output(7, 91) <= input(10);
output(7, 92) <= input(11);
output(7, 93) <= input(12);
output(7, 94) <= input(13);
output(7, 95) <= input(14);
output(7, 96) <= input(36);
output(7, 97) <= input(0);
output(7, 98) <= input(1);
output(7, 99) <= input(2);
output(7, 100) <= input(3);
output(7, 101) <= input(4);
output(7, 102) <= input(5);
output(7, 103) <= input(6);
output(7, 104) <= input(7);
output(7, 105) <= input(8);
output(7, 106) <= input(9);
output(7, 107) <= input(10);
output(7, 108) <= input(11);
output(7, 109) <= input(12);
output(7, 110) <= input(13);
output(7, 111) <= input(14);
output(7, 112) <= input(36);
output(7, 113) <= input(0);
output(7, 114) <= input(1);
output(7, 115) <= input(2);
output(7, 116) <= input(3);
output(7, 117) <= input(4);
output(7, 118) <= input(5);
output(7, 119) <= input(6);
output(7, 120) <= input(7);
output(7, 121) <= input(8);
output(7, 122) <= input(9);
output(7, 123) <= input(10);
output(7, 124) <= input(11);
output(7, 125) <= input(12);
output(7, 126) <= input(13);
output(7, 127) <= input(14);
output(7, 128) <= input(36);
output(7, 129) <= input(0);
output(7, 130) <= input(1);
output(7, 131) <= input(2);
output(7, 132) <= input(3);
output(7, 133) <= input(4);
output(7, 134) <= input(5);
output(7, 135) <= input(6);
output(7, 136) <= input(7);
output(7, 137) <= input(8);
output(7, 138) <= input(9);
output(7, 139) <= input(10);
output(7, 140) <= input(11);
output(7, 141) <= input(12);
output(7, 142) <= input(13);
output(7, 143) <= input(14);
output(7, 144) <= input(36);
output(7, 145) <= input(0);
output(7, 146) <= input(1);
output(7, 147) <= input(2);
output(7, 148) <= input(3);
output(7, 149) <= input(4);
output(7, 150) <= input(5);
output(7, 151) <= input(6);
output(7, 152) <= input(7);
output(7, 153) <= input(8);
output(7, 154) <= input(9);
output(7, 155) <= input(10);
output(7, 156) <= input(11);
output(7, 157) <= input(12);
output(7, 158) <= input(13);
output(7, 159) <= input(14);
output(7, 160) <= input(37);
output(7, 161) <= input(35);
output(7, 162) <= input(16);
output(7, 163) <= input(17);
output(7, 164) <= input(18);
output(7, 165) <= input(19);
output(7, 166) <= input(20);
output(7, 167) <= input(21);
output(7, 168) <= input(22);
output(7, 169) <= input(23);
output(7, 170) <= input(24);
output(7, 171) <= input(25);
output(7, 172) <= input(26);
output(7, 173) <= input(27);
output(7, 174) <= input(28);
output(7, 175) <= input(29);
output(7, 176) <= input(37);
output(7, 177) <= input(35);
output(7, 178) <= input(16);
output(7, 179) <= input(17);
output(7, 180) <= input(18);
output(7, 181) <= input(19);
output(7, 182) <= input(20);
output(7, 183) <= input(21);
output(7, 184) <= input(22);
output(7, 185) <= input(23);
output(7, 186) <= input(24);
output(7, 187) <= input(25);
output(7, 188) <= input(26);
output(7, 189) <= input(27);
output(7, 190) <= input(28);
output(7, 191) <= input(29);
output(7, 192) <= input(37);
output(7, 193) <= input(35);
output(7, 194) <= input(16);
output(7, 195) <= input(17);
output(7, 196) <= input(18);
output(7, 197) <= input(19);
output(7, 198) <= input(20);
output(7, 199) <= input(21);
output(7, 200) <= input(22);
output(7, 201) <= input(23);
output(7, 202) <= input(24);
output(7, 203) <= input(25);
output(7, 204) <= input(26);
output(7, 205) <= input(27);
output(7, 206) <= input(28);
output(7, 207) <= input(29);
output(7, 208) <= input(37);
output(7, 209) <= input(35);
output(7, 210) <= input(16);
output(7, 211) <= input(17);
output(7, 212) <= input(18);
output(7, 213) <= input(19);
output(7, 214) <= input(20);
output(7, 215) <= input(21);
output(7, 216) <= input(22);
output(7, 217) <= input(23);
output(7, 218) <= input(24);
output(7, 219) <= input(25);
output(7, 220) <= input(26);
output(7, 221) <= input(27);
output(7, 222) <= input(28);
output(7, 223) <= input(29);
output(7, 224) <= input(37);
output(7, 225) <= input(35);
output(7, 226) <= input(16);
output(7, 227) <= input(17);
output(7, 228) <= input(18);
output(7, 229) <= input(19);
output(7, 230) <= input(20);
output(7, 231) <= input(21);
output(7, 232) <= input(22);
output(7, 233) <= input(23);
output(7, 234) <= input(24);
output(7, 235) <= input(25);
output(7, 236) <= input(26);
output(7, 237) <= input(27);
output(7, 238) <= input(28);
output(7, 239) <= input(29);
output(7, 240) <= input(37);
output(7, 241) <= input(35);
output(7, 242) <= input(16);
output(7, 243) <= input(17);
output(7, 244) <= input(18);
output(7, 245) <= input(19);
output(7, 246) <= input(20);
output(7, 247) <= input(21);
output(7, 248) <= input(22);
output(7, 249) <= input(23);
output(7, 250) <= input(24);
output(7, 251) <= input(25);
output(7, 252) <= input(26);
output(7, 253) <= input(27);
output(7, 254) <= input(28);
output(7, 255) <= input(29);
when "0011" =>
output(0, 0) <= input(0);
output(0, 1) <= input(1);
output(0, 2) <= input(2);
output(0, 3) <= input(3);
output(0, 4) <= input(4);
output(0, 5) <= input(5);
output(0, 6) <= input(6);
output(0, 7) <= input(7);
output(0, 8) <= input(8);
output(0, 9) <= input(9);
output(0, 10) <= input(10);
output(0, 11) <= input(11);
output(0, 12) <= input(12);
output(0, 13) <= input(13);
output(0, 14) <= input(14);
output(0, 15) <= input(15);
output(0, 16) <= input(0);
output(0, 17) <= input(1);
output(0, 18) <= input(2);
output(0, 19) <= input(3);
output(0, 20) <= input(4);
output(0, 21) <= input(5);
output(0, 22) <= input(6);
output(0, 23) <= input(7);
output(0, 24) <= input(8);
output(0, 25) <= input(9);
output(0, 26) <= input(10);
output(0, 27) <= input(11);
output(0, 28) <= input(12);
output(0, 29) <= input(13);
output(0, 30) <= input(14);
output(0, 31) <= input(15);
output(0, 32) <= input(0);
output(0, 33) <= input(1);
output(0, 34) <= input(2);
output(0, 35) <= input(3);
output(0, 36) <= input(4);
output(0, 37) <= input(5);
output(0, 38) <= input(6);
output(0, 39) <= input(7);
output(0, 40) <= input(8);
output(0, 41) <= input(9);
output(0, 42) <= input(10);
output(0, 43) <= input(11);
output(0, 44) <= input(12);
output(0, 45) <= input(13);
output(0, 46) <= input(14);
output(0, 47) <= input(15);
output(0, 48) <= input(0);
output(0, 49) <= input(1);
output(0, 50) <= input(2);
output(0, 51) <= input(3);
output(0, 52) <= input(4);
output(0, 53) <= input(5);
output(0, 54) <= input(6);
output(0, 55) <= input(7);
output(0, 56) <= input(8);
output(0, 57) <= input(9);
output(0, 58) <= input(10);
output(0, 59) <= input(11);
output(0, 60) <= input(12);
output(0, 61) <= input(13);
output(0, 62) <= input(14);
output(0, 63) <= input(15);
output(0, 64) <= input(16);
output(0, 65) <= input(17);
output(0, 66) <= input(18);
output(0, 67) <= input(19);
output(0, 68) <= input(20);
output(0, 69) <= input(21);
output(0, 70) <= input(22);
output(0, 71) <= input(23);
output(0, 72) <= input(24);
output(0, 73) <= input(25);
output(0, 74) <= input(26);
output(0, 75) <= input(27);
output(0, 76) <= input(28);
output(0, 77) <= input(29);
output(0, 78) <= input(30);
output(0, 79) <= input(31);
output(0, 80) <= input(16);
output(0, 81) <= input(17);
output(0, 82) <= input(18);
output(0, 83) <= input(19);
output(0, 84) <= input(20);
output(0, 85) <= input(21);
output(0, 86) <= input(22);
output(0, 87) <= input(23);
output(0, 88) <= input(24);
output(0, 89) <= input(25);
output(0, 90) <= input(26);
output(0, 91) <= input(27);
output(0, 92) <= input(28);
output(0, 93) <= input(29);
output(0, 94) <= input(30);
output(0, 95) <= input(31);
output(0, 96) <= input(16);
output(0, 97) <= input(17);
output(0, 98) <= input(18);
output(0, 99) <= input(19);
output(0, 100) <= input(20);
output(0, 101) <= input(21);
output(0, 102) <= input(22);
output(0, 103) <= input(23);
output(0, 104) <= input(24);
output(0, 105) <= input(25);
output(0, 106) <= input(26);
output(0, 107) <= input(27);
output(0, 108) <= input(28);
output(0, 109) <= input(29);
output(0, 110) <= input(30);
output(0, 111) <= input(31);
output(0, 112) <= input(16);
output(0, 113) <= input(17);
output(0, 114) <= input(18);
output(0, 115) <= input(19);
output(0, 116) <= input(20);
output(0, 117) <= input(21);
output(0, 118) <= input(22);
output(0, 119) <= input(23);
output(0, 120) <= input(24);
output(0, 121) <= input(25);
output(0, 122) <= input(26);
output(0, 123) <= input(27);
output(0, 124) <= input(28);
output(0, 125) <= input(29);
output(0, 126) <= input(30);
output(0, 127) <= input(31);
output(0, 128) <= input(32);
output(0, 129) <= input(0);
output(0, 130) <= input(1);
output(0, 131) <= input(2);
output(0, 132) <= input(3);
output(0, 133) <= input(4);
output(0, 134) <= input(5);
output(0, 135) <= input(6);
output(0, 136) <= input(7);
output(0, 137) <= input(8);
output(0, 138) <= input(9);
output(0, 139) <= input(10);
output(0, 140) <= input(11);
output(0, 141) <= input(12);
output(0, 142) <= input(13);
output(0, 143) <= input(14);
output(0, 144) <= input(32);
output(0, 145) <= input(0);
output(0, 146) <= input(1);
output(0, 147) <= input(2);
output(0, 148) <= input(3);
output(0, 149) <= input(4);
output(0, 150) <= input(5);
output(0, 151) <= input(6);
output(0, 152) <= input(7);
output(0, 153) <= input(8);
output(0, 154) <= input(9);
output(0, 155) <= input(10);
output(0, 156) <= input(11);
output(0, 157) <= input(12);
output(0, 158) <= input(13);
output(0, 159) <= input(14);
output(0, 160) <= input(32);
output(0, 161) <= input(0);
output(0, 162) <= input(1);
output(0, 163) <= input(2);
output(0, 164) <= input(3);
output(0, 165) <= input(4);
output(0, 166) <= input(5);
output(0, 167) <= input(6);
output(0, 168) <= input(7);
output(0, 169) <= input(8);
output(0, 170) <= input(9);
output(0, 171) <= input(10);
output(0, 172) <= input(11);
output(0, 173) <= input(12);
output(0, 174) <= input(13);
output(0, 175) <= input(14);
output(0, 176) <= input(32);
output(0, 177) <= input(0);
output(0, 178) <= input(1);
output(0, 179) <= input(2);
output(0, 180) <= input(3);
output(0, 181) <= input(4);
output(0, 182) <= input(5);
output(0, 183) <= input(6);
output(0, 184) <= input(7);
output(0, 185) <= input(8);
output(0, 186) <= input(9);
output(0, 187) <= input(10);
output(0, 188) <= input(11);
output(0, 189) <= input(12);
output(0, 190) <= input(13);
output(0, 191) <= input(14);
output(0, 192) <= input(33);
output(0, 193) <= input(16);
output(0, 194) <= input(17);
output(0, 195) <= input(18);
output(0, 196) <= input(19);
output(0, 197) <= input(20);
output(0, 198) <= input(21);
output(0, 199) <= input(22);
output(0, 200) <= input(23);
output(0, 201) <= input(24);
output(0, 202) <= input(25);
output(0, 203) <= input(26);
output(0, 204) <= input(27);
output(0, 205) <= input(28);
output(0, 206) <= input(29);
output(0, 207) <= input(30);
output(0, 208) <= input(33);
output(0, 209) <= input(16);
output(0, 210) <= input(17);
output(0, 211) <= input(18);
output(0, 212) <= input(19);
output(0, 213) <= input(20);
output(0, 214) <= input(21);
output(0, 215) <= input(22);
output(0, 216) <= input(23);
output(0, 217) <= input(24);
output(0, 218) <= input(25);
output(0, 219) <= input(26);
output(0, 220) <= input(27);
output(0, 221) <= input(28);
output(0, 222) <= input(29);
output(0, 223) <= input(30);
output(0, 224) <= input(33);
output(0, 225) <= input(16);
output(0, 226) <= input(17);
output(0, 227) <= input(18);
output(0, 228) <= input(19);
output(0, 229) <= input(20);
output(0, 230) <= input(21);
output(0, 231) <= input(22);
output(0, 232) <= input(23);
output(0, 233) <= input(24);
output(0, 234) <= input(25);
output(0, 235) <= input(26);
output(0, 236) <= input(27);
output(0, 237) <= input(28);
output(0, 238) <= input(29);
output(0, 239) <= input(30);
output(0, 240) <= input(33);
output(0, 241) <= input(16);
output(0, 242) <= input(17);
output(0, 243) <= input(18);
output(0, 244) <= input(19);
output(0, 245) <= input(20);
output(0, 246) <= input(21);
output(0, 247) <= input(22);
output(0, 248) <= input(23);
output(0, 249) <= input(24);
output(0, 250) <= input(25);
output(0, 251) <= input(26);
output(0, 252) <= input(27);
output(0, 253) <= input(28);
output(0, 254) <= input(29);
output(0, 255) <= input(30);
output(1, 0) <= input(0);
output(1, 1) <= input(1);
output(1, 2) <= input(2);
output(1, 3) <= input(3);
output(1, 4) <= input(4);
output(1, 5) <= input(5);
output(1, 6) <= input(6);
output(1, 7) <= input(7);
output(1, 8) <= input(8);
output(1, 9) <= input(9);
output(1, 10) <= input(10);
output(1, 11) <= input(11);
output(1, 12) <= input(12);
output(1, 13) <= input(13);
output(1, 14) <= input(14);
output(1, 15) <= input(15);
output(1, 16) <= input(0);
output(1, 17) <= input(1);
output(1, 18) <= input(2);
output(1, 19) <= input(3);
output(1, 20) <= input(4);
output(1, 21) <= input(5);
output(1, 22) <= input(6);
output(1, 23) <= input(7);
output(1, 24) <= input(8);
output(1, 25) <= input(9);
output(1, 26) <= input(10);
output(1, 27) <= input(11);
output(1, 28) <= input(12);
output(1, 29) <= input(13);
output(1, 30) <= input(14);
output(1, 31) <= input(15);
output(1, 32) <= input(16);
output(1, 33) <= input(17);
output(1, 34) <= input(18);
output(1, 35) <= input(19);
output(1, 36) <= input(20);
output(1, 37) <= input(21);
output(1, 38) <= input(22);
output(1, 39) <= input(23);
output(1, 40) <= input(24);
output(1, 41) <= input(25);
output(1, 42) <= input(26);
output(1, 43) <= input(27);
output(1, 44) <= input(28);
output(1, 45) <= input(29);
output(1, 46) <= input(30);
output(1, 47) <= input(31);
output(1, 48) <= input(16);
output(1, 49) <= input(17);
output(1, 50) <= input(18);
output(1, 51) <= input(19);
output(1, 52) <= input(20);
output(1, 53) <= input(21);
output(1, 54) <= input(22);
output(1, 55) <= input(23);
output(1, 56) <= input(24);
output(1, 57) <= input(25);
output(1, 58) <= input(26);
output(1, 59) <= input(27);
output(1, 60) <= input(28);
output(1, 61) <= input(29);
output(1, 62) <= input(30);
output(1, 63) <= input(31);
output(1, 64) <= input(16);
output(1, 65) <= input(17);
output(1, 66) <= input(18);
output(1, 67) <= input(19);
output(1, 68) <= input(20);
output(1, 69) <= input(21);
output(1, 70) <= input(22);
output(1, 71) <= input(23);
output(1, 72) <= input(24);
output(1, 73) <= input(25);
output(1, 74) <= input(26);
output(1, 75) <= input(27);
output(1, 76) <= input(28);
output(1, 77) <= input(29);
output(1, 78) <= input(30);
output(1, 79) <= input(31);
output(1, 80) <= input(32);
output(1, 81) <= input(0);
output(1, 82) <= input(1);
output(1, 83) <= input(2);
output(1, 84) <= input(3);
output(1, 85) <= input(4);
output(1, 86) <= input(5);
output(1, 87) <= input(6);
output(1, 88) <= input(7);
output(1, 89) <= input(8);
output(1, 90) <= input(9);
output(1, 91) <= input(10);
output(1, 92) <= input(11);
output(1, 93) <= input(12);
output(1, 94) <= input(13);
output(1, 95) <= input(14);
output(1, 96) <= input(32);
output(1, 97) <= input(0);
output(1, 98) <= input(1);
output(1, 99) <= input(2);
output(1, 100) <= input(3);
output(1, 101) <= input(4);
output(1, 102) <= input(5);
output(1, 103) <= input(6);
output(1, 104) <= input(7);
output(1, 105) <= input(8);
output(1, 106) <= input(9);
output(1, 107) <= input(10);
output(1, 108) <= input(11);
output(1, 109) <= input(12);
output(1, 110) <= input(13);
output(1, 111) <= input(14);
output(1, 112) <= input(32);
output(1, 113) <= input(0);
output(1, 114) <= input(1);
output(1, 115) <= input(2);
output(1, 116) <= input(3);
output(1, 117) <= input(4);
output(1, 118) <= input(5);
output(1, 119) <= input(6);
output(1, 120) <= input(7);
output(1, 121) <= input(8);
output(1, 122) <= input(9);
output(1, 123) <= input(10);
output(1, 124) <= input(11);
output(1, 125) <= input(12);
output(1, 126) <= input(13);
output(1, 127) <= input(14);
output(1, 128) <= input(33);
output(1, 129) <= input(16);
output(1, 130) <= input(17);
output(1, 131) <= input(18);
output(1, 132) <= input(19);
output(1, 133) <= input(20);
output(1, 134) <= input(21);
output(1, 135) <= input(22);
output(1, 136) <= input(23);
output(1, 137) <= input(24);
output(1, 138) <= input(25);
output(1, 139) <= input(26);
output(1, 140) <= input(27);
output(1, 141) <= input(28);
output(1, 142) <= input(29);
output(1, 143) <= input(30);
output(1, 144) <= input(33);
output(1, 145) <= input(16);
output(1, 146) <= input(17);
output(1, 147) <= input(18);
output(1, 148) <= input(19);
output(1, 149) <= input(20);
output(1, 150) <= input(21);
output(1, 151) <= input(22);
output(1, 152) <= input(23);
output(1, 153) <= input(24);
output(1, 154) <= input(25);
output(1, 155) <= input(26);
output(1, 156) <= input(27);
output(1, 157) <= input(28);
output(1, 158) <= input(29);
output(1, 159) <= input(30);
output(1, 160) <= input(34);
output(1, 161) <= input(32);
output(1, 162) <= input(0);
output(1, 163) <= input(1);
output(1, 164) <= input(2);
output(1, 165) <= input(3);
output(1, 166) <= input(4);
output(1, 167) <= input(5);
output(1, 168) <= input(6);
output(1, 169) <= input(7);
output(1, 170) <= input(8);
output(1, 171) <= input(9);
output(1, 172) <= input(10);
output(1, 173) <= input(11);
output(1, 174) <= input(12);
output(1, 175) <= input(13);
output(1, 176) <= input(34);
output(1, 177) <= input(32);
output(1, 178) <= input(0);
output(1, 179) <= input(1);
output(1, 180) <= input(2);
output(1, 181) <= input(3);
output(1, 182) <= input(4);
output(1, 183) <= input(5);
output(1, 184) <= input(6);
output(1, 185) <= input(7);
output(1, 186) <= input(8);
output(1, 187) <= input(9);
output(1, 188) <= input(10);
output(1, 189) <= input(11);
output(1, 190) <= input(12);
output(1, 191) <= input(13);
output(1, 192) <= input(34);
output(1, 193) <= input(32);
output(1, 194) <= input(0);
output(1, 195) <= input(1);
output(1, 196) <= input(2);
output(1, 197) <= input(3);
output(1, 198) <= input(4);
output(1, 199) <= input(5);
output(1, 200) <= input(6);
output(1, 201) <= input(7);
output(1, 202) <= input(8);
output(1, 203) <= input(9);
output(1, 204) <= input(10);
output(1, 205) <= input(11);
output(1, 206) <= input(12);
output(1, 207) <= input(13);
output(1, 208) <= input(35);
output(1, 209) <= input(33);
output(1, 210) <= input(16);
output(1, 211) <= input(17);
output(1, 212) <= input(18);
output(1, 213) <= input(19);
output(1, 214) <= input(20);
output(1, 215) <= input(21);
output(1, 216) <= input(22);
output(1, 217) <= input(23);
output(1, 218) <= input(24);
output(1, 219) <= input(25);
output(1, 220) <= input(26);
output(1, 221) <= input(27);
output(1, 222) <= input(28);
output(1, 223) <= input(29);
output(1, 224) <= input(35);
output(1, 225) <= input(33);
output(1, 226) <= input(16);
output(1, 227) <= input(17);
output(1, 228) <= input(18);
output(1, 229) <= input(19);
output(1, 230) <= input(20);
output(1, 231) <= input(21);
output(1, 232) <= input(22);
output(1, 233) <= input(23);
output(1, 234) <= input(24);
output(1, 235) <= input(25);
output(1, 236) <= input(26);
output(1, 237) <= input(27);
output(1, 238) <= input(28);
output(1, 239) <= input(29);
output(1, 240) <= input(35);
output(1, 241) <= input(33);
output(1, 242) <= input(16);
output(1, 243) <= input(17);
output(1, 244) <= input(18);
output(1, 245) <= input(19);
output(1, 246) <= input(20);
output(1, 247) <= input(21);
output(1, 248) <= input(22);
output(1, 249) <= input(23);
output(1, 250) <= input(24);
output(1, 251) <= input(25);
output(1, 252) <= input(26);
output(1, 253) <= input(27);
output(1, 254) <= input(28);
output(1, 255) <= input(29);
output(2, 0) <= input(0);
output(2, 1) <= input(1);
output(2, 2) <= input(2);
output(2, 3) <= input(3);
output(2, 4) <= input(4);
output(2, 5) <= input(5);
output(2, 6) <= input(6);
output(2, 7) <= input(7);
output(2, 8) <= input(8);
output(2, 9) <= input(9);
output(2, 10) <= input(10);
output(2, 11) <= input(11);
output(2, 12) <= input(12);
output(2, 13) <= input(13);
output(2, 14) <= input(14);
output(2, 15) <= input(15);
output(2, 16) <= input(0);
output(2, 17) <= input(1);
output(2, 18) <= input(2);
output(2, 19) <= input(3);
output(2, 20) <= input(4);
output(2, 21) <= input(5);
output(2, 22) <= input(6);
output(2, 23) <= input(7);
output(2, 24) <= input(8);
output(2, 25) <= input(9);
output(2, 26) <= input(10);
output(2, 27) <= input(11);
output(2, 28) <= input(12);
output(2, 29) <= input(13);
output(2, 30) <= input(14);
output(2, 31) <= input(15);
output(2, 32) <= input(16);
output(2, 33) <= input(17);
output(2, 34) <= input(18);
output(2, 35) <= input(19);
output(2, 36) <= input(20);
output(2, 37) <= input(21);
output(2, 38) <= input(22);
output(2, 39) <= input(23);
output(2, 40) <= input(24);
output(2, 41) <= input(25);
output(2, 42) <= input(26);
output(2, 43) <= input(27);
output(2, 44) <= input(28);
output(2, 45) <= input(29);
output(2, 46) <= input(30);
output(2, 47) <= input(31);
output(2, 48) <= input(16);
output(2, 49) <= input(17);
output(2, 50) <= input(18);
output(2, 51) <= input(19);
output(2, 52) <= input(20);
output(2, 53) <= input(21);
output(2, 54) <= input(22);
output(2, 55) <= input(23);
output(2, 56) <= input(24);
output(2, 57) <= input(25);
output(2, 58) <= input(26);
output(2, 59) <= input(27);
output(2, 60) <= input(28);
output(2, 61) <= input(29);
output(2, 62) <= input(30);
output(2, 63) <= input(31);
output(2, 64) <= input(32);
output(2, 65) <= input(0);
output(2, 66) <= input(1);
output(2, 67) <= input(2);
output(2, 68) <= input(3);
output(2, 69) <= input(4);
output(2, 70) <= input(5);
output(2, 71) <= input(6);
output(2, 72) <= input(7);
output(2, 73) <= input(8);
output(2, 74) <= input(9);
output(2, 75) <= input(10);
output(2, 76) <= input(11);
output(2, 77) <= input(12);
output(2, 78) <= input(13);
output(2, 79) <= input(14);
output(2, 80) <= input(32);
output(2, 81) <= input(0);
output(2, 82) <= input(1);
output(2, 83) <= input(2);
output(2, 84) <= input(3);
output(2, 85) <= input(4);
output(2, 86) <= input(5);
output(2, 87) <= input(6);
output(2, 88) <= input(7);
output(2, 89) <= input(8);
output(2, 90) <= input(9);
output(2, 91) <= input(10);
output(2, 92) <= input(11);
output(2, 93) <= input(12);
output(2, 94) <= input(13);
output(2, 95) <= input(14);
output(2, 96) <= input(33);
output(2, 97) <= input(16);
output(2, 98) <= input(17);
output(2, 99) <= input(18);
output(2, 100) <= input(19);
output(2, 101) <= input(20);
output(2, 102) <= input(21);
output(2, 103) <= input(22);
output(2, 104) <= input(23);
output(2, 105) <= input(24);
output(2, 106) <= input(25);
output(2, 107) <= input(26);
output(2, 108) <= input(27);
output(2, 109) <= input(28);
output(2, 110) <= input(29);
output(2, 111) <= input(30);
output(2, 112) <= input(33);
output(2, 113) <= input(16);
output(2, 114) <= input(17);
output(2, 115) <= input(18);
output(2, 116) <= input(19);
output(2, 117) <= input(20);
output(2, 118) <= input(21);
output(2, 119) <= input(22);
output(2, 120) <= input(23);
output(2, 121) <= input(24);
output(2, 122) <= input(25);
output(2, 123) <= input(26);
output(2, 124) <= input(27);
output(2, 125) <= input(28);
output(2, 126) <= input(29);
output(2, 127) <= input(30);
output(2, 128) <= input(34);
output(2, 129) <= input(32);
output(2, 130) <= input(0);
output(2, 131) <= input(1);
output(2, 132) <= input(2);
output(2, 133) <= input(3);
output(2, 134) <= input(4);
output(2, 135) <= input(5);
output(2, 136) <= input(6);
output(2, 137) <= input(7);
output(2, 138) <= input(8);
output(2, 139) <= input(9);
output(2, 140) <= input(10);
output(2, 141) <= input(11);
output(2, 142) <= input(12);
output(2, 143) <= input(13);
output(2, 144) <= input(34);
output(2, 145) <= input(32);
output(2, 146) <= input(0);
output(2, 147) <= input(1);
output(2, 148) <= input(2);
output(2, 149) <= input(3);
output(2, 150) <= input(4);
output(2, 151) <= input(5);
output(2, 152) <= input(6);
output(2, 153) <= input(7);
output(2, 154) <= input(8);
output(2, 155) <= input(9);
output(2, 156) <= input(10);
output(2, 157) <= input(11);
output(2, 158) <= input(12);
output(2, 159) <= input(13);
output(2, 160) <= input(35);
output(2, 161) <= input(33);
output(2, 162) <= input(16);
output(2, 163) <= input(17);
output(2, 164) <= input(18);
output(2, 165) <= input(19);
output(2, 166) <= input(20);
output(2, 167) <= input(21);
output(2, 168) <= input(22);
output(2, 169) <= input(23);
output(2, 170) <= input(24);
output(2, 171) <= input(25);
output(2, 172) <= input(26);
output(2, 173) <= input(27);
output(2, 174) <= input(28);
output(2, 175) <= input(29);
output(2, 176) <= input(35);
output(2, 177) <= input(33);
output(2, 178) <= input(16);
output(2, 179) <= input(17);
output(2, 180) <= input(18);
output(2, 181) <= input(19);
output(2, 182) <= input(20);
output(2, 183) <= input(21);
output(2, 184) <= input(22);
output(2, 185) <= input(23);
output(2, 186) <= input(24);
output(2, 187) <= input(25);
output(2, 188) <= input(26);
output(2, 189) <= input(27);
output(2, 190) <= input(28);
output(2, 191) <= input(29);
output(2, 192) <= input(36);
output(2, 193) <= input(34);
output(2, 194) <= input(32);
output(2, 195) <= input(0);
output(2, 196) <= input(1);
output(2, 197) <= input(2);
output(2, 198) <= input(3);
output(2, 199) <= input(4);
output(2, 200) <= input(5);
output(2, 201) <= input(6);
output(2, 202) <= input(7);
output(2, 203) <= input(8);
output(2, 204) <= input(9);
output(2, 205) <= input(10);
output(2, 206) <= input(11);
output(2, 207) <= input(12);
output(2, 208) <= input(36);
output(2, 209) <= input(34);
output(2, 210) <= input(32);
output(2, 211) <= input(0);
output(2, 212) <= input(1);
output(2, 213) <= input(2);
output(2, 214) <= input(3);
output(2, 215) <= input(4);
output(2, 216) <= input(5);
output(2, 217) <= input(6);
output(2, 218) <= input(7);
output(2, 219) <= input(8);
output(2, 220) <= input(9);
output(2, 221) <= input(10);
output(2, 222) <= input(11);
output(2, 223) <= input(12);
output(2, 224) <= input(37);
output(2, 225) <= input(35);
output(2, 226) <= input(33);
output(2, 227) <= input(16);
output(2, 228) <= input(17);
output(2, 229) <= input(18);
output(2, 230) <= input(19);
output(2, 231) <= input(20);
output(2, 232) <= input(21);
output(2, 233) <= input(22);
output(2, 234) <= input(23);
output(2, 235) <= input(24);
output(2, 236) <= input(25);
output(2, 237) <= input(26);
output(2, 238) <= input(27);
output(2, 239) <= input(28);
output(2, 240) <= input(37);
output(2, 241) <= input(35);
output(2, 242) <= input(33);
output(2, 243) <= input(16);
output(2, 244) <= input(17);
output(2, 245) <= input(18);
output(2, 246) <= input(19);
output(2, 247) <= input(20);
output(2, 248) <= input(21);
output(2, 249) <= input(22);
output(2, 250) <= input(23);
output(2, 251) <= input(24);
output(2, 252) <= input(25);
output(2, 253) <= input(26);
output(2, 254) <= input(27);
output(2, 255) <= input(28);
when "0100" =>
output(0, 0) <= input(0);
output(0, 1) <= input(1);
output(0, 2) <= input(2);
output(0, 3) <= input(3);
output(0, 4) <= input(4);
output(0, 5) <= input(5);
output(0, 6) <= input(6);
output(0, 7) <= input(7);
output(0, 8) <= input(8);
output(0, 9) <= input(9);
output(0, 10) <= input(10);
output(0, 11) <= input(11);
output(0, 12) <= input(12);
output(0, 13) <= input(13);
output(0, 14) <= input(14);
output(0, 15) <= input(15);
output(0, 16) <= input(16);
output(0, 17) <= input(17);
output(0, 18) <= input(18);
output(0, 19) <= input(19);
output(0, 20) <= input(20);
output(0, 21) <= input(21);
output(0, 22) <= input(22);
output(0, 23) <= input(23);
output(0, 24) <= input(24);
output(0, 25) <= input(25);
output(0, 26) <= input(26);
output(0, 27) <= input(27);
output(0, 28) <= input(28);
output(0, 29) <= input(29);
output(0, 30) <= input(30);
output(0, 31) <= input(31);
output(0, 32) <= input(16);
output(0, 33) <= input(17);
output(0, 34) <= input(18);
output(0, 35) <= input(19);
output(0, 36) <= input(20);
output(0, 37) <= input(21);
output(0, 38) <= input(22);
output(0, 39) <= input(23);
output(0, 40) <= input(24);
output(0, 41) <= input(25);
output(0, 42) <= input(26);
output(0, 43) <= input(27);
output(0, 44) <= input(28);
output(0, 45) <= input(29);
output(0, 46) <= input(30);
output(0, 47) <= input(31);
output(0, 48) <= input(32);
output(0, 49) <= input(0);
output(0, 50) <= input(1);
output(0, 51) <= input(2);
output(0, 52) <= input(3);
output(0, 53) <= input(4);
output(0, 54) <= input(5);
output(0, 55) <= input(6);
output(0, 56) <= input(7);
output(0, 57) <= input(8);
output(0, 58) <= input(9);
output(0, 59) <= input(10);
output(0, 60) <= input(11);
output(0, 61) <= input(12);
output(0, 62) <= input(13);
output(0, 63) <= input(14);
output(0, 64) <= input(33);
output(0, 65) <= input(16);
output(0, 66) <= input(17);
output(0, 67) <= input(18);
output(0, 68) <= input(19);
output(0, 69) <= input(20);
output(0, 70) <= input(21);
output(0, 71) <= input(22);
output(0, 72) <= input(23);
output(0, 73) <= input(24);
output(0, 74) <= input(25);
output(0, 75) <= input(26);
output(0, 76) <= input(27);
output(0, 77) <= input(28);
output(0, 78) <= input(29);
output(0, 79) <= input(30);
output(0, 80) <= input(33);
output(0, 81) <= input(16);
output(0, 82) <= input(17);
output(0, 83) <= input(18);
output(0, 84) <= input(19);
output(0, 85) <= input(20);
output(0, 86) <= input(21);
output(0, 87) <= input(22);
output(0, 88) <= input(23);
output(0, 89) <= input(24);
output(0, 90) <= input(25);
output(0, 91) <= input(26);
output(0, 92) <= input(27);
output(0, 93) <= input(28);
output(0, 94) <= input(29);
output(0, 95) <= input(30);
output(0, 96) <= input(34);
output(0, 97) <= input(32);
output(0, 98) <= input(0);
output(0, 99) <= input(1);
output(0, 100) <= input(2);
output(0, 101) <= input(3);
output(0, 102) <= input(4);
output(0, 103) <= input(5);
output(0, 104) <= input(6);
output(0, 105) <= input(7);
output(0, 106) <= input(8);
output(0, 107) <= input(9);
output(0, 108) <= input(10);
output(0, 109) <= input(11);
output(0, 110) <= input(12);
output(0, 111) <= input(13);
output(0, 112) <= input(34);
output(0, 113) <= input(32);
output(0, 114) <= input(0);
output(0, 115) <= input(1);
output(0, 116) <= input(2);
output(0, 117) <= input(3);
output(0, 118) <= input(4);
output(0, 119) <= input(5);
output(0, 120) <= input(6);
output(0, 121) <= input(7);
output(0, 122) <= input(8);
output(0, 123) <= input(9);
output(0, 124) <= input(10);
output(0, 125) <= input(11);
output(0, 126) <= input(12);
output(0, 127) <= input(13);
output(0, 128) <= input(35);
output(0, 129) <= input(33);
output(0, 130) <= input(16);
output(0, 131) <= input(17);
output(0, 132) <= input(18);
output(0, 133) <= input(19);
output(0, 134) <= input(20);
output(0, 135) <= input(21);
output(0, 136) <= input(22);
output(0, 137) <= input(23);
output(0, 138) <= input(24);
output(0, 139) <= input(25);
output(0, 140) <= input(26);
output(0, 141) <= input(27);
output(0, 142) <= input(28);
output(0, 143) <= input(29);
output(0, 144) <= input(36);
output(0, 145) <= input(34);
output(0, 146) <= input(32);
output(0, 147) <= input(0);
output(0, 148) <= input(1);
output(0, 149) <= input(2);
output(0, 150) <= input(3);
output(0, 151) <= input(4);
output(0, 152) <= input(5);
output(0, 153) <= input(6);
output(0, 154) <= input(7);
output(0, 155) <= input(8);
output(0, 156) <= input(9);
output(0, 157) <= input(10);
output(0, 158) <= input(11);
output(0, 159) <= input(12);
output(0, 160) <= input(36);
output(0, 161) <= input(34);
output(0, 162) <= input(32);
output(0, 163) <= input(0);
output(0, 164) <= input(1);
output(0, 165) <= input(2);
output(0, 166) <= input(3);
output(0, 167) <= input(4);
output(0, 168) <= input(5);
output(0, 169) <= input(6);
output(0, 170) <= input(7);
output(0, 171) <= input(8);
output(0, 172) <= input(9);
output(0, 173) <= input(10);
output(0, 174) <= input(11);
output(0, 175) <= input(12);
output(0, 176) <= input(37);
output(0, 177) <= input(35);
output(0, 178) <= input(33);
output(0, 179) <= input(16);
output(0, 180) <= input(17);
output(0, 181) <= input(18);
output(0, 182) <= input(19);
output(0, 183) <= input(20);
output(0, 184) <= input(21);
output(0, 185) <= input(22);
output(0, 186) <= input(23);
output(0, 187) <= input(24);
output(0, 188) <= input(25);
output(0, 189) <= input(26);
output(0, 190) <= input(27);
output(0, 191) <= input(28);
output(0, 192) <= input(38);
output(0, 193) <= input(36);
output(0, 194) <= input(34);
output(0, 195) <= input(32);
output(0, 196) <= input(0);
output(0, 197) <= input(1);
output(0, 198) <= input(2);
output(0, 199) <= input(3);
output(0, 200) <= input(4);
output(0, 201) <= input(5);
output(0, 202) <= input(6);
output(0, 203) <= input(7);
output(0, 204) <= input(8);
output(0, 205) <= input(9);
output(0, 206) <= input(10);
output(0, 207) <= input(11);
output(0, 208) <= input(38);
output(0, 209) <= input(36);
output(0, 210) <= input(34);
output(0, 211) <= input(32);
output(0, 212) <= input(0);
output(0, 213) <= input(1);
output(0, 214) <= input(2);
output(0, 215) <= input(3);
output(0, 216) <= input(4);
output(0, 217) <= input(5);
output(0, 218) <= input(6);
output(0, 219) <= input(7);
output(0, 220) <= input(8);
output(0, 221) <= input(9);
output(0, 222) <= input(10);
output(0, 223) <= input(11);
output(0, 224) <= input(39);
output(0, 225) <= input(37);
output(0, 226) <= input(35);
output(0, 227) <= input(33);
output(0, 228) <= input(16);
output(0, 229) <= input(17);
output(0, 230) <= input(18);
output(0, 231) <= input(19);
output(0, 232) <= input(20);
output(0, 233) <= input(21);
output(0, 234) <= input(22);
output(0, 235) <= input(23);
output(0, 236) <= input(24);
output(0, 237) <= input(25);
output(0, 238) <= input(26);
output(0, 239) <= input(27);
output(0, 240) <= input(39);
output(0, 241) <= input(37);
output(0, 242) <= input(35);
output(0, 243) <= input(33);
output(0, 244) <= input(16);
output(0, 245) <= input(17);
output(0, 246) <= input(18);
output(0, 247) <= input(19);
output(0, 248) <= input(20);
output(0, 249) <= input(21);
output(0, 250) <= input(22);
output(0, 251) <= input(23);
output(0, 252) <= input(24);
output(0, 253) <= input(25);
output(0, 254) <= input(26);
output(0, 255) <= input(27);
output(1, 0) <= input(0);
output(1, 1) <= input(1);
output(1, 2) <= input(2);
output(1, 3) <= input(3);
output(1, 4) <= input(4);
output(1, 5) <= input(5);
output(1, 6) <= input(6);
output(1, 7) <= input(7);
output(1, 8) <= input(8);
output(1, 9) <= input(9);
output(1, 10) <= input(10);
output(1, 11) <= input(11);
output(1, 12) <= input(12);
output(1, 13) <= input(13);
output(1, 14) <= input(14);
output(1, 15) <= input(15);
output(1, 16) <= input(16);
output(1, 17) <= input(17);
output(1, 18) <= input(18);
output(1, 19) <= input(19);
output(1, 20) <= input(20);
output(1, 21) <= input(21);
output(1, 22) <= input(22);
output(1, 23) <= input(23);
output(1, 24) <= input(24);
output(1, 25) <= input(25);
output(1, 26) <= input(26);
output(1, 27) <= input(27);
output(1, 28) <= input(28);
output(1, 29) <= input(29);
output(1, 30) <= input(30);
output(1, 31) <= input(31);
output(1, 32) <= input(32);
output(1, 33) <= input(0);
output(1, 34) <= input(1);
output(1, 35) <= input(2);
output(1, 36) <= input(3);
output(1, 37) <= input(4);
output(1, 38) <= input(5);
output(1, 39) <= input(6);
output(1, 40) <= input(7);
output(1, 41) <= input(8);
output(1, 42) <= input(9);
output(1, 43) <= input(10);
output(1, 44) <= input(11);
output(1, 45) <= input(12);
output(1, 46) <= input(13);
output(1, 47) <= input(14);
output(1, 48) <= input(32);
output(1, 49) <= input(0);
output(1, 50) <= input(1);
output(1, 51) <= input(2);
output(1, 52) <= input(3);
output(1, 53) <= input(4);
output(1, 54) <= input(5);
output(1, 55) <= input(6);
output(1, 56) <= input(7);
output(1, 57) <= input(8);
output(1, 58) <= input(9);
output(1, 59) <= input(10);
output(1, 60) <= input(11);
output(1, 61) <= input(12);
output(1, 62) <= input(13);
output(1, 63) <= input(14);
output(1, 64) <= input(33);
output(1, 65) <= input(16);
output(1, 66) <= input(17);
output(1, 67) <= input(18);
output(1, 68) <= input(19);
output(1, 69) <= input(20);
output(1, 70) <= input(21);
output(1, 71) <= input(22);
output(1, 72) <= input(23);
output(1, 73) <= input(24);
output(1, 74) <= input(25);
output(1, 75) <= input(26);
output(1, 76) <= input(27);
output(1, 77) <= input(28);
output(1, 78) <= input(29);
output(1, 79) <= input(30);
output(1, 80) <= input(34);
output(1, 81) <= input(32);
output(1, 82) <= input(0);
output(1, 83) <= input(1);
output(1, 84) <= input(2);
output(1, 85) <= input(3);
output(1, 86) <= input(4);
output(1, 87) <= input(5);
output(1, 88) <= input(6);
output(1, 89) <= input(7);
output(1, 90) <= input(8);
output(1, 91) <= input(9);
output(1, 92) <= input(10);
output(1, 93) <= input(11);
output(1, 94) <= input(12);
output(1, 95) <= input(13);
output(1, 96) <= input(35);
output(1, 97) <= input(33);
output(1, 98) <= input(16);
output(1, 99) <= input(17);
output(1, 100) <= input(18);
output(1, 101) <= input(19);
output(1, 102) <= input(20);
output(1, 103) <= input(21);
output(1, 104) <= input(22);
output(1, 105) <= input(23);
output(1, 106) <= input(24);
output(1, 107) <= input(25);
output(1, 108) <= input(26);
output(1, 109) <= input(27);
output(1, 110) <= input(28);
output(1, 111) <= input(29);
output(1, 112) <= input(35);
output(1, 113) <= input(33);
output(1, 114) <= input(16);
output(1, 115) <= input(17);
output(1, 116) <= input(18);
output(1, 117) <= input(19);
output(1, 118) <= input(20);
output(1, 119) <= input(21);
output(1, 120) <= input(22);
output(1, 121) <= input(23);
output(1, 122) <= input(24);
output(1, 123) <= input(25);
output(1, 124) <= input(26);
output(1, 125) <= input(27);
output(1, 126) <= input(28);
output(1, 127) <= input(29);
output(1, 128) <= input(36);
output(1, 129) <= input(34);
output(1, 130) <= input(32);
output(1, 131) <= input(0);
output(1, 132) <= input(1);
output(1, 133) <= input(2);
output(1, 134) <= input(3);
output(1, 135) <= input(4);
output(1, 136) <= input(5);
output(1, 137) <= input(6);
output(1, 138) <= input(7);
output(1, 139) <= input(8);
output(1, 140) <= input(9);
output(1, 141) <= input(10);
output(1, 142) <= input(11);
output(1, 143) <= input(12);
output(1, 144) <= input(37);
output(1, 145) <= input(35);
output(1, 146) <= input(33);
output(1, 147) <= input(16);
output(1, 148) <= input(17);
output(1, 149) <= input(18);
output(1, 150) <= input(19);
output(1, 151) <= input(20);
output(1, 152) <= input(21);
output(1, 153) <= input(22);
output(1, 154) <= input(23);
output(1, 155) <= input(24);
output(1, 156) <= input(25);
output(1, 157) <= input(26);
output(1, 158) <= input(27);
output(1, 159) <= input(28);
output(1, 160) <= input(38);
output(1, 161) <= input(36);
output(1, 162) <= input(34);
output(1, 163) <= input(32);
output(1, 164) <= input(0);
output(1, 165) <= input(1);
output(1, 166) <= input(2);
output(1, 167) <= input(3);
output(1, 168) <= input(4);
output(1, 169) <= input(5);
output(1, 170) <= input(6);
output(1, 171) <= input(7);
output(1, 172) <= input(8);
output(1, 173) <= input(9);
output(1, 174) <= input(10);
output(1, 175) <= input(11);
output(1, 176) <= input(38);
output(1, 177) <= input(36);
output(1, 178) <= input(34);
output(1, 179) <= input(32);
output(1, 180) <= input(0);
output(1, 181) <= input(1);
output(1, 182) <= input(2);
output(1, 183) <= input(3);
output(1, 184) <= input(4);
output(1, 185) <= input(5);
output(1, 186) <= input(6);
output(1, 187) <= input(7);
output(1, 188) <= input(8);
output(1, 189) <= input(9);
output(1, 190) <= input(10);
output(1, 191) <= input(11);
output(1, 192) <= input(39);
output(1, 193) <= input(37);
output(1, 194) <= input(35);
output(1, 195) <= input(33);
output(1, 196) <= input(16);
output(1, 197) <= input(17);
output(1, 198) <= input(18);
output(1, 199) <= input(19);
output(1, 200) <= input(20);
output(1, 201) <= input(21);
output(1, 202) <= input(22);
output(1, 203) <= input(23);
output(1, 204) <= input(24);
output(1, 205) <= input(25);
output(1, 206) <= input(26);
output(1, 207) <= input(27);
output(1, 208) <= input(40);
output(1, 209) <= input(38);
output(1, 210) <= input(36);
output(1, 211) <= input(34);
output(1, 212) <= input(32);
output(1, 213) <= input(0);
output(1, 214) <= input(1);
output(1, 215) <= input(2);
output(1, 216) <= input(3);
output(1, 217) <= input(4);
output(1, 218) <= input(5);
output(1, 219) <= input(6);
output(1, 220) <= input(7);
output(1, 221) <= input(8);
output(1, 222) <= input(9);
output(1, 223) <= input(10);
output(1, 224) <= input(41);
output(1, 225) <= input(39);
output(1, 226) <= input(37);
output(1, 227) <= input(35);
output(1, 228) <= input(33);
output(1, 229) <= input(16);
output(1, 230) <= input(17);
output(1, 231) <= input(18);
output(1, 232) <= input(19);
output(1, 233) <= input(20);
output(1, 234) <= input(21);
output(1, 235) <= input(22);
output(1, 236) <= input(23);
output(1, 237) <= input(24);
output(1, 238) <= input(25);
output(1, 239) <= input(26);
output(1, 240) <= input(41);
output(1, 241) <= input(39);
output(1, 242) <= input(37);
output(1, 243) <= input(35);
output(1, 244) <= input(33);
output(1, 245) <= input(16);
output(1, 246) <= input(17);
output(1, 247) <= input(18);
output(1, 248) <= input(19);
output(1, 249) <= input(20);
output(1, 250) <= input(21);
output(1, 251) <= input(22);
output(1, 252) <= input(23);
output(1, 253) <= input(24);
output(1, 254) <= input(25);
output(1, 255) <= input(26);
output(2, 0) <= input(0);
output(2, 1) <= input(1);
output(2, 2) <= input(2);
output(2, 3) <= input(3);
output(2, 4) <= input(4);
output(2, 5) <= input(5);
output(2, 6) <= input(6);
output(2, 7) <= input(7);
output(2, 8) <= input(8);
output(2, 9) <= input(9);
output(2, 10) <= input(10);
output(2, 11) <= input(11);
output(2, 12) <= input(12);
output(2, 13) <= input(13);
output(2, 14) <= input(14);
output(2, 15) <= input(15);
output(2, 16) <= input(16);
output(2, 17) <= input(17);
output(2, 18) <= input(18);
output(2, 19) <= input(19);
output(2, 20) <= input(20);
output(2, 21) <= input(21);
output(2, 22) <= input(22);
output(2, 23) <= input(23);
output(2, 24) <= input(24);
output(2, 25) <= input(25);
output(2, 26) <= input(26);
output(2, 27) <= input(27);
output(2, 28) <= input(28);
output(2, 29) <= input(29);
output(2, 30) <= input(30);
output(2, 31) <= input(31);
output(2, 32) <= input(32);
output(2, 33) <= input(0);
output(2, 34) <= input(1);
output(2, 35) <= input(2);
output(2, 36) <= input(3);
output(2, 37) <= input(4);
output(2, 38) <= input(5);
output(2, 39) <= input(6);
output(2, 40) <= input(7);
output(2, 41) <= input(8);
output(2, 42) <= input(9);
output(2, 43) <= input(10);
output(2, 44) <= input(11);
output(2, 45) <= input(12);
output(2, 46) <= input(13);
output(2, 47) <= input(14);
output(2, 48) <= input(33);
output(2, 49) <= input(16);
output(2, 50) <= input(17);
output(2, 51) <= input(18);
output(2, 52) <= input(19);
output(2, 53) <= input(20);
output(2, 54) <= input(21);
output(2, 55) <= input(22);
output(2, 56) <= input(23);
output(2, 57) <= input(24);
output(2, 58) <= input(25);
output(2, 59) <= input(26);
output(2, 60) <= input(27);
output(2, 61) <= input(28);
output(2, 62) <= input(29);
output(2, 63) <= input(30);
output(2, 64) <= input(34);
output(2, 65) <= input(32);
output(2, 66) <= input(0);
output(2, 67) <= input(1);
output(2, 68) <= input(2);
output(2, 69) <= input(3);
output(2, 70) <= input(4);
output(2, 71) <= input(5);
output(2, 72) <= input(6);
output(2, 73) <= input(7);
output(2, 74) <= input(8);
output(2, 75) <= input(9);
output(2, 76) <= input(10);
output(2, 77) <= input(11);
output(2, 78) <= input(12);
output(2, 79) <= input(13);
output(2, 80) <= input(35);
output(2, 81) <= input(33);
output(2, 82) <= input(16);
output(2, 83) <= input(17);
output(2, 84) <= input(18);
output(2, 85) <= input(19);
output(2, 86) <= input(20);
output(2, 87) <= input(21);
output(2, 88) <= input(22);
output(2, 89) <= input(23);
output(2, 90) <= input(24);
output(2, 91) <= input(25);
output(2, 92) <= input(26);
output(2, 93) <= input(27);
output(2, 94) <= input(28);
output(2, 95) <= input(29);
output(2, 96) <= input(36);
output(2, 97) <= input(34);
output(2, 98) <= input(32);
output(2, 99) <= input(0);
output(2, 100) <= input(1);
output(2, 101) <= input(2);
output(2, 102) <= input(3);
output(2, 103) <= input(4);
output(2, 104) <= input(5);
output(2, 105) <= input(6);
output(2, 106) <= input(7);
output(2, 107) <= input(8);
output(2, 108) <= input(9);
output(2, 109) <= input(10);
output(2, 110) <= input(11);
output(2, 111) <= input(12);
output(2, 112) <= input(36);
output(2, 113) <= input(34);
output(2, 114) <= input(32);
output(2, 115) <= input(0);
output(2, 116) <= input(1);
output(2, 117) <= input(2);
output(2, 118) <= input(3);
output(2, 119) <= input(4);
output(2, 120) <= input(5);
output(2, 121) <= input(6);
output(2, 122) <= input(7);
output(2, 123) <= input(8);
output(2, 124) <= input(9);
output(2, 125) <= input(10);
output(2, 126) <= input(11);
output(2, 127) <= input(12);
output(2, 128) <= input(37);
output(2, 129) <= input(35);
output(2, 130) <= input(33);
output(2, 131) <= input(16);
output(2, 132) <= input(17);
output(2, 133) <= input(18);
output(2, 134) <= input(19);
output(2, 135) <= input(20);
output(2, 136) <= input(21);
output(2, 137) <= input(22);
output(2, 138) <= input(23);
output(2, 139) <= input(24);
output(2, 140) <= input(25);
output(2, 141) <= input(26);
output(2, 142) <= input(27);
output(2, 143) <= input(28);
output(2, 144) <= input(38);
output(2, 145) <= input(36);
output(2, 146) <= input(34);
output(2, 147) <= input(32);
output(2, 148) <= input(0);
output(2, 149) <= input(1);
output(2, 150) <= input(2);
output(2, 151) <= input(3);
output(2, 152) <= input(4);
output(2, 153) <= input(5);
output(2, 154) <= input(6);
output(2, 155) <= input(7);
output(2, 156) <= input(8);
output(2, 157) <= input(9);
output(2, 158) <= input(10);
output(2, 159) <= input(11);
output(2, 160) <= input(39);
output(2, 161) <= input(37);
output(2, 162) <= input(35);
output(2, 163) <= input(33);
output(2, 164) <= input(16);
output(2, 165) <= input(17);
output(2, 166) <= input(18);
output(2, 167) <= input(19);
output(2, 168) <= input(20);
output(2, 169) <= input(21);
output(2, 170) <= input(22);
output(2, 171) <= input(23);
output(2, 172) <= input(24);
output(2, 173) <= input(25);
output(2, 174) <= input(26);
output(2, 175) <= input(27);
output(2, 176) <= input(40);
output(2, 177) <= input(38);
output(2, 178) <= input(36);
output(2, 179) <= input(34);
output(2, 180) <= input(32);
output(2, 181) <= input(0);
output(2, 182) <= input(1);
output(2, 183) <= input(2);
output(2, 184) <= input(3);
output(2, 185) <= input(4);
output(2, 186) <= input(5);
output(2, 187) <= input(6);
output(2, 188) <= input(7);
output(2, 189) <= input(8);
output(2, 190) <= input(9);
output(2, 191) <= input(10);
output(2, 192) <= input(41);
output(2, 193) <= input(39);
output(2, 194) <= input(37);
output(2, 195) <= input(35);
output(2, 196) <= input(33);
output(2, 197) <= input(16);
output(2, 198) <= input(17);
output(2, 199) <= input(18);
output(2, 200) <= input(19);
output(2, 201) <= input(20);
output(2, 202) <= input(21);
output(2, 203) <= input(22);
output(2, 204) <= input(23);
output(2, 205) <= input(24);
output(2, 206) <= input(25);
output(2, 207) <= input(26);
output(2, 208) <= input(42);
output(2, 209) <= input(40);
output(2, 210) <= input(38);
output(2, 211) <= input(36);
output(2, 212) <= input(34);
output(2, 213) <= input(32);
output(2, 214) <= input(0);
output(2, 215) <= input(1);
output(2, 216) <= input(2);
output(2, 217) <= input(3);
output(2, 218) <= input(4);
output(2, 219) <= input(5);
output(2, 220) <= input(6);
output(2, 221) <= input(7);
output(2, 222) <= input(8);
output(2, 223) <= input(9);
output(2, 224) <= input(43);
output(2, 225) <= input(41);
output(2, 226) <= input(39);
output(2, 227) <= input(37);
output(2, 228) <= input(35);
output(2, 229) <= input(33);
output(2, 230) <= input(16);
output(2, 231) <= input(17);
output(2, 232) <= input(18);
output(2, 233) <= input(19);
output(2, 234) <= input(20);
output(2, 235) <= input(21);
output(2, 236) <= input(22);
output(2, 237) <= input(23);
output(2, 238) <= input(24);
output(2, 239) <= input(25);
output(2, 240) <= input(43);
output(2, 241) <= input(41);
output(2, 242) <= input(39);
output(2, 243) <= input(37);
output(2, 244) <= input(35);
output(2, 245) <= input(33);
output(2, 246) <= input(16);
output(2, 247) <= input(17);
output(2, 248) <= input(18);
output(2, 249) <= input(19);
output(2, 250) <= input(20);
output(2, 251) <= input(21);
output(2, 252) <= input(22);
output(2, 253) <= input(23);
output(2, 254) <= input(24);
output(2, 255) <= input(25);
when "0101" =>
output(0, 0) <= input(0);
output(0, 1) <= input(1);
output(0, 2) <= input(2);
output(0, 3) <= input(3);
output(0, 4) <= input(4);
output(0, 5) <= input(5);
output(0, 6) <= input(6);
output(0, 7) <= input(7);
output(0, 8) <= input(8);
output(0, 9) <= input(9);
output(0, 10) <= input(10);
output(0, 11) <= input(11);
output(0, 12) <= input(12);
output(0, 13) <= input(13);
output(0, 14) <= input(14);
output(0, 15) <= input(15);
output(0, 16) <= input(16);
output(0, 17) <= input(17);
output(0, 18) <= input(18);
output(0, 19) <= input(19);
output(0, 20) <= input(20);
output(0, 21) <= input(21);
output(0, 22) <= input(22);
output(0, 23) <= input(23);
output(0, 24) <= input(24);
output(0, 25) <= input(25);
output(0, 26) <= input(26);
output(0, 27) <= input(27);
output(0, 28) <= input(28);
output(0, 29) <= input(29);
output(0, 30) <= input(30);
output(0, 31) <= input(31);
output(0, 32) <= input(32);
output(0, 33) <= input(0);
output(0, 34) <= input(1);
output(0, 35) <= input(2);
output(0, 36) <= input(3);
output(0, 37) <= input(4);
output(0, 38) <= input(5);
output(0, 39) <= input(6);
output(0, 40) <= input(7);
output(0, 41) <= input(8);
output(0, 42) <= input(9);
output(0, 43) <= input(10);
output(0, 44) <= input(11);
output(0, 45) <= input(12);
output(0, 46) <= input(13);
output(0, 47) <= input(14);
output(0, 48) <= input(33);
output(0, 49) <= input(16);
output(0, 50) <= input(17);
output(0, 51) <= input(18);
output(0, 52) <= input(19);
output(0, 53) <= input(20);
output(0, 54) <= input(21);
output(0, 55) <= input(22);
output(0, 56) <= input(23);
output(0, 57) <= input(24);
output(0, 58) <= input(25);
output(0, 59) <= input(26);
output(0, 60) <= input(27);
output(0, 61) <= input(28);
output(0, 62) <= input(29);
output(0, 63) <= input(30);
output(0, 64) <= input(34);
output(0, 65) <= input(32);
output(0, 66) <= input(0);
output(0, 67) <= input(1);
output(0, 68) <= input(2);
output(0, 69) <= input(3);
output(0, 70) <= input(4);
output(0, 71) <= input(5);
output(0, 72) <= input(6);
output(0, 73) <= input(7);
output(0, 74) <= input(8);
output(0, 75) <= input(9);
output(0, 76) <= input(10);
output(0, 77) <= input(11);
output(0, 78) <= input(12);
output(0, 79) <= input(13);
output(0, 80) <= input(35);
output(0, 81) <= input(33);
output(0, 82) <= input(16);
output(0, 83) <= input(17);
output(0, 84) <= input(18);
output(0, 85) <= input(19);
output(0, 86) <= input(20);
output(0, 87) <= input(21);
output(0, 88) <= input(22);
output(0, 89) <= input(23);
output(0, 90) <= input(24);
output(0, 91) <= input(25);
output(0, 92) <= input(26);
output(0, 93) <= input(27);
output(0, 94) <= input(28);
output(0, 95) <= input(29);
output(0, 96) <= input(36);
output(0, 97) <= input(34);
output(0, 98) <= input(32);
output(0, 99) <= input(0);
output(0, 100) <= input(1);
output(0, 101) <= input(2);
output(0, 102) <= input(3);
output(0, 103) <= input(4);
output(0, 104) <= input(5);
output(0, 105) <= input(6);
output(0, 106) <= input(7);
output(0, 107) <= input(8);
output(0, 108) <= input(9);
output(0, 109) <= input(10);
output(0, 110) <= input(11);
output(0, 111) <= input(12);
output(0, 112) <= input(37);
output(0, 113) <= input(35);
output(0, 114) <= input(33);
output(0, 115) <= input(16);
output(0, 116) <= input(17);
output(0, 117) <= input(18);
output(0, 118) <= input(19);
output(0, 119) <= input(20);
output(0, 120) <= input(21);
output(0, 121) <= input(22);
output(0, 122) <= input(23);
output(0, 123) <= input(24);
output(0, 124) <= input(25);
output(0, 125) <= input(26);
output(0, 126) <= input(27);
output(0, 127) <= input(28);
output(0, 128) <= input(38);
output(0, 129) <= input(36);
output(0, 130) <= input(34);
output(0, 131) <= input(32);
output(0, 132) <= input(0);
output(0, 133) <= input(1);
output(0, 134) <= input(2);
output(0, 135) <= input(3);
output(0, 136) <= input(4);
output(0, 137) <= input(5);
output(0, 138) <= input(6);
output(0, 139) <= input(7);
output(0, 140) <= input(8);
output(0, 141) <= input(9);
output(0, 142) <= input(10);
output(0, 143) <= input(11);
output(0, 144) <= input(39);
output(0, 145) <= input(37);
output(0, 146) <= input(35);
output(0, 147) <= input(33);
output(0, 148) <= input(16);
output(0, 149) <= input(17);
output(0, 150) <= input(18);
output(0, 151) <= input(19);
output(0, 152) <= input(20);
output(0, 153) <= input(21);
output(0, 154) <= input(22);
output(0, 155) <= input(23);
output(0, 156) <= input(24);
output(0, 157) <= input(25);
output(0, 158) <= input(26);
output(0, 159) <= input(27);
output(0, 160) <= input(40);
output(0, 161) <= input(38);
output(0, 162) <= input(36);
output(0, 163) <= input(34);
output(0, 164) <= input(32);
output(0, 165) <= input(0);
output(0, 166) <= input(1);
output(0, 167) <= input(2);
output(0, 168) <= input(3);
output(0, 169) <= input(4);
output(0, 170) <= input(5);
output(0, 171) <= input(6);
output(0, 172) <= input(7);
output(0, 173) <= input(8);
output(0, 174) <= input(9);
output(0, 175) <= input(10);
output(0, 176) <= input(41);
output(0, 177) <= input(39);
output(0, 178) <= input(37);
output(0, 179) <= input(35);
output(0, 180) <= input(33);
output(0, 181) <= input(16);
output(0, 182) <= input(17);
output(0, 183) <= input(18);
output(0, 184) <= input(19);
output(0, 185) <= input(20);
output(0, 186) <= input(21);
output(0, 187) <= input(22);
output(0, 188) <= input(23);
output(0, 189) <= input(24);
output(0, 190) <= input(25);
output(0, 191) <= input(26);
output(0, 192) <= input(42);
output(0, 193) <= input(40);
output(0, 194) <= input(38);
output(0, 195) <= input(36);
output(0, 196) <= input(34);
output(0, 197) <= input(32);
output(0, 198) <= input(0);
output(0, 199) <= input(1);
output(0, 200) <= input(2);
output(0, 201) <= input(3);
output(0, 202) <= input(4);
output(0, 203) <= input(5);
output(0, 204) <= input(6);
output(0, 205) <= input(7);
output(0, 206) <= input(8);
output(0, 207) <= input(9);
output(0, 208) <= input(43);
output(0, 209) <= input(41);
output(0, 210) <= input(39);
output(0, 211) <= input(37);
output(0, 212) <= input(35);
output(0, 213) <= input(33);
output(0, 214) <= input(16);
output(0, 215) <= input(17);
output(0, 216) <= input(18);
output(0, 217) <= input(19);
output(0, 218) <= input(20);
output(0, 219) <= input(21);
output(0, 220) <= input(22);
output(0, 221) <= input(23);
output(0, 222) <= input(24);
output(0, 223) <= input(25);
output(0, 224) <= input(44);
output(0, 225) <= input(42);
output(0, 226) <= input(40);
output(0, 227) <= input(38);
output(0, 228) <= input(36);
output(0, 229) <= input(34);
output(0, 230) <= input(32);
output(0, 231) <= input(0);
output(0, 232) <= input(1);
output(0, 233) <= input(2);
output(0, 234) <= input(3);
output(0, 235) <= input(4);
output(0, 236) <= input(5);
output(0, 237) <= input(6);
output(0, 238) <= input(7);
output(0, 239) <= input(8);
output(0, 240) <= input(45);
output(0, 241) <= input(43);
output(0, 242) <= input(41);
output(0, 243) <= input(39);
output(0, 244) <= input(37);
output(0, 245) <= input(35);
output(0, 246) <= input(33);
output(0, 247) <= input(16);
output(0, 248) <= input(17);
output(0, 249) <= input(18);
output(0, 250) <= input(19);
output(0, 251) <= input(20);
output(0, 252) <= input(21);
output(0, 253) <= input(22);
output(0, 254) <= input(23);
output(0, 255) <= input(24);
output(1, 0) <= input(16);
output(1, 1) <= input(17);
output(1, 2) <= input(18);
output(1, 3) <= input(19);
output(1, 4) <= input(20);
output(1, 5) <= input(21);
output(1, 6) <= input(22);
output(1, 7) <= input(23);
output(1, 8) <= input(24);
output(1, 9) <= input(25);
output(1, 10) <= input(26);
output(1, 11) <= input(27);
output(1, 12) <= input(28);
output(1, 13) <= input(29);
output(1, 14) <= input(30);
output(1, 15) <= input(31);
output(1, 16) <= input(32);
output(1, 17) <= input(0);
output(1, 18) <= input(1);
output(1, 19) <= input(2);
output(1, 20) <= input(3);
output(1, 21) <= input(4);
output(1, 22) <= input(5);
output(1, 23) <= input(6);
output(1, 24) <= input(7);
output(1, 25) <= input(8);
output(1, 26) <= input(9);
output(1, 27) <= input(10);
output(1, 28) <= input(11);
output(1, 29) <= input(12);
output(1, 30) <= input(13);
output(1, 31) <= input(14);
output(1, 32) <= input(33);
output(1, 33) <= input(16);
output(1, 34) <= input(17);
output(1, 35) <= input(18);
output(1, 36) <= input(19);
output(1, 37) <= input(20);
output(1, 38) <= input(21);
output(1, 39) <= input(22);
output(1, 40) <= input(23);
output(1, 41) <= input(24);
output(1, 42) <= input(25);
output(1, 43) <= input(26);
output(1, 44) <= input(27);
output(1, 45) <= input(28);
output(1, 46) <= input(29);
output(1, 47) <= input(30);
output(1, 48) <= input(34);
output(1, 49) <= input(32);
output(1, 50) <= input(0);
output(1, 51) <= input(1);
output(1, 52) <= input(2);
output(1, 53) <= input(3);
output(1, 54) <= input(4);
output(1, 55) <= input(5);
output(1, 56) <= input(6);
output(1, 57) <= input(7);
output(1, 58) <= input(8);
output(1, 59) <= input(9);
output(1, 60) <= input(10);
output(1, 61) <= input(11);
output(1, 62) <= input(12);
output(1, 63) <= input(13);
output(1, 64) <= input(35);
output(1, 65) <= input(33);
output(1, 66) <= input(16);
output(1, 67) <= input(17);
output(1, 68) <= input(18);
output(1, 69) <= input(19);
output(1, 70) <= input(20);
output(1, 71) <= input(21);
output(1, 72) <= input(22);
output(1, 73) <= input(23);
output(1, 74) <= input(24);
output(1, 75) <= input(25);
output(1, 76) <= input(26);
output(1, 77) <= input(27);
output(1, 78) <= input(28);
output(1, 79) <= input(29);
output(1, 80) <= input(36);
output(1, 81) <= input(34);
output(1, 82) <= input(32);
output(1, 83) <= input(0);
output(1, 84) <= input(1);
output(1, 85) <= input(2);
output(1, 86) <= input(3);
output(1, 87) <= input(4);
output(1, 88) <= input(5);
output(1, 89) <= input(6);
output(1, 90) <= input(7);
output(1, 91) <= input(8);
output(1, 92) <= input(9);
output(1, 93) <= input(10);
output(1, 94) <= input(11);
output(1, 95) <= input(12);
output(1, 96) <= input(37);
output(1, 97) <= input(35);
output(1, 98) <= input(33);
output(1, 99) <= input(16);
output(1, 100) <= input(17);
output(1, 101) <= input(18);
output(1, 102) <= input(19);
output(1, 103) <= input(20);
output(1, 104) <= input(21);
output(1, 105) <= input(22);
output(1, 106) <= input(23);
output(1, 107) <= input(24);
output(1, 108) <= input(25);
output(1, 109) <= input(26);
output(1, 110) <= input(27);
output(1, 111) <= input(28);
output(1, 112) <= input(38);
output(1, 113) <= input(36);
output(1, 114) <= input(34);
output(1, 115) <= input(32);
output(1, 116) <= input(0);
output(1, 117) <= input(1);
output(1, 118) <= input(2);
output(1, 119) <= input(3);
output(1, 120) <= input(4);
output(1, 121) <= input(5);
output(1, 122) <= input(6);
output(1, 123) <= input(7);
output(1, 124) <= input(8);
output(1, 125) <= input(9);
output(1, 126) <= input(10);
output(1, 127) <= input(11);
output(1, 128) <= input(40);
output(1, 129) <= input(38);
output(1, 130) <= input(36);
output(1, 131) <= input(34);
output(1, 132) <= input(32);
output(1, 133) <= input(0);
output(1, 134) <= input(1);
output(1, 135) <= input(2);
output(1, 136) <= input(3);
output(1, 137) <= input(4);
output(1, 138) <= input(5);
output(1, 139) <= input(6);
output(1, 140) <= input(7);
output(1, 141) <= input(8);
output(1, 142) <= input(9);
output(1, 143) <= input(10);
output(1, 144) <= input(41);
output(1, 145) <= input(39);
output(1, 146) <= input(37);
output(1, 147) <= input(35);
output(1, 148) <= input(33);
output(1, 149) <= input(16);
output(1, 150) <= input(17);
output(1, 151) <= input(18);
output(1, 152) <= input(19);
output(1, 153) <= input(20);
output(1, 154) <= input(21);
output(1, 155) <= input(22);
output(1, 156) <= input(23);
output(1, 157) <= input(24);
output(1, 158) <= input(25);
output(1, 159) <= input(26);
output(1, 160) <= input(42);
output(1, 161) <= input(40);
output(1, 162) <= input(38);
output(1, 163) <= input(36);
output(1, 164) <= input(34);
output(1, 165) <= input(32);
output(1, 166) <= input(0);
output(1, 167) <= input(1);
output(1, 168) <= input(2);
output(1, 169) <= input(3);
output(1, 170) <= input(4);
output(1, 171) <= input(5);
output(1, 172) <= input(6);
output(1, 173) <= input(7);
output(1, 174) <= input(8);
output(1, 175) <= input(9);
output(1, 176) <= input(43);
output(1, 177) <= input(41);
output(1, 178) <= input(39);
output(1, 179) <= input(37);
output(1, 180) <= input(35);
output(1, 181) <= input(33);
output(1, 182) <= input(16);
output(1, 183) <= input(17);
output(1, 184) <= input(18);
output(1, 185) <= input(19);
output(1, 186) <= input(20);
output(1, 187) <= input(21);
output(1, 188) <= input(22);
output(1, 189) <= input(23);
output(1, 190) <= input(24);
output(1, 191) <= input(25);
output(1, 192) <= input(44);
output(1, 193) <= input(42);
output(1, 194) <= input(40);
output(1, 195) <= input(38);
output(1, 196) <= input(36);
output(1, 197) <= input(34);
output(1, 198) <= input(32);
output(1, 199) <= input(0);
output(1, 200) <= input(1);
output(1, 201) <= input(2);
output(1, 202) <= input(3);
output(1, 203) <= input(4);
output(1, 204) <= input(5);
output(1, 205) <= input(6);
output(1, 206) <= input(7);
output(1, 207) <= input(8);
output(1, 208) <= input(45);
output(1, 209) <= input(43);
output(1, 210) <= input(41);
output(1, 211) <= input(39);
output(1, 212) <= input(37);
output(1, 213) <= input(35);
output(1, 214) <= input(33);
output(1, 215) <= input(16);
output(1, 216) <= input(17);
output(1, 217) <= input(18);
output(1, 218) <= input(19);
output(1, 219) <= input(20);
output(1, 220) <= input(21);
output(1, 221) <= input(22);
output(1, 222) <= input(23);
output(1, 223) <= input(24);
output(1, 224) <= input(46);
output(1, 225) <= input(44);
output(1, 226) <= input(42);
output(1, 227) <= input(40);
output(1, 228) <= input(38);
output(1, 229) <= input(36);
output(1, 230) <= input(34);
output(1, 231) <= input(32);
output(1, 232) <= input(0);
output(1, 233) <= input(1);
output(1, 234) <= input(2);
output(1, 235) <= input(3);
output(1, 236) <= input(4);
output(1, 237) <= input(5);
output(1, 238) <= input(6);
output(1, 239) <= input(7);
output(1, 240) <= input(47);
output(1, 241) <= input(45);
output(1, 242) <= input(43);
output(1, 243) <= input(41);
output(1, 244) <= input(39);
output(1, 245) <= input(37);
output(1, 246) <= input(35);
output(1, 247) <= input(33);
output(1, 248) <= input(16);
output(1, 249) <= input(17);
output(1, 250) <= input(18);
output(1, 251) <= input(19);
output(1, 252) <= input(20);
output(1, 253) <= input(21);
output(1, 254) <= input(22);
output(1, 255) <= input(23);
when "0110" =>
output(0, 0) <= input(0);
output(0, 1) <= input(1);
output(0, 2) <= input(2);
output(0, 3) <= input(3);
output(0, 4) <= input(4);
output(0, 5) <= input(5);
output(0, 6) <= input(6);
output(0, 7) <= input(7);
output(0, 8) <= input(8);
output(0, 9) <= input(9);
output(0, 10) <= input(10);
output(0, 11) <= input(11);
output(0, 12) <= input(12);
output(0, 13) <= input(13);
output(0, 14) <= input(14);
output(0, 15) <= input(15);
output(0, 16) <= input(16);
output(0, 17) <= input(17);
output(0, 18) <= input(18);
output(0, 19) <= input(19);
output(0, 20) <= input(20);
output(0, 21) <= input(21);
output(0, 22) <= input(22);
output(0, 23) <= input(23);
output(0, 24) <= input(24);
output(0, 25) <= input(25);
output(0, 26) <= input(26);
output(0, 27) <= input(27);
output(0, 28) <= input(28);
output(0, 29) <= input(29);
output(0, 30) <= input(30);
output(0, 31) <= input(31);
output(0, 32) <= input(32);
output(0, 33) <= input(0);
output(0, 34) <= input(1);
output(0, 35) <= input(2);
output(0, 36) <= input(3);
output(0, 37) <= input(4);
output(0, 38) <= input(5);
output(0, 39) <= input(6);
output(0, 40) <= input(7);
output(0, 41) <= input(8);
output(0, 42) <= input(9);
output(0, 43) <= input(10);
output(0, 44) <= input(11);
output(0, 45) <= input(12);
output(0, 46) <= input(13);
output(0, 47) <= input(14);
output(0, 48) <= input(33);
output(0, 49) <= input(16);
output(0, 50) <= input(17);
output(0, 51) <= input(18);
output(0, 52) <= input(19);
output(0, 53) <= input(20);
output(0, 54) <= input(21);
output(0, 55) <= input(22);
output(0, 56) <= input(23);
output(0, 57) <= input(24);
output(0, 58) <= input(25);
output(0, 59) <= input(26);
output(0, 60) <= input(27);
output(0, 61) <= input(28);
output(0, 62) <= input(29);
output(0, 63) <= input(30);
output(0, 64) <= input(34);
output(0, 65) <= input(33);
output(0, 66) <= input(16);
output(0, 67) <= input(17);
output(0, 68) <= input(18);
output(0, 69) <= input(19);
output(0, 70) <= input(20);
output(0, 71) <= input(21);
output(0, 72) <= input(22);
output(0, 73) <= input(23);
output(0, 74) <= input(24);
output(0, 75) <= input(25);
output(0, 76) <= input(26);
output(0, 77) <= input(27);
output(0, 78) <= input(28);
output(0, 79) <= input(29);
output(0, 80) <= input(35);
output(0, 81) <= input(36);
output(0, 82) <= input(32);
output(0, 83) <= input(0);
output(0, 84) <= input(1);
output(0, 85) <= input(2);
output(0, 86) <= input(3);
output(0, 87) <= input(4);
output(0, 88) <= input(5);
output(0, 89) <= input(6);
output(0, 90) <= input(7);
output(0, 91) <= input(8);
output(0, 92) <= input(9);
output(0, 93) <= input(10);
output(0, 94) <= input(11);
output(0, 95) <= input(12);
output(0, 96) <= input(37);
output(0, 97) <= input(34);
output(0, 98) <= input(33);
output(0, 99) <= input(16);
output(0, 100) <= input(17);
output(0, 101) <= input(18);
output(0, 102) <= input(19);
output(0, 103) <= input(20);
output(0, 104) <= input(21);
output(0, 105) <= input(22);
output(0, 106) <= input(23);
output(0, 107) <= input(24);
output(0, 108) <= input(25);
output(0, 109) <= input(26);
output(0, 110) <= input(27);
output(0, 111) <= input(28);
output(0, 112) <= input(38);
output(0, 113) <= input(35);
output(0, 114) <= input(36);
output(0, 115) <= input(32);
output(0, 116) <= input(0);
output(0, 117) <= input(1);
output(0, 118) <= input(2);
output(0, 119) <= input(3);
output(0, 120) <= input(4);
output(0, 121) <= input(5);
output(0, 122) <= input(6);
output(0, 123) <= input(7);
output(0, 124) <= input(8);
output(0, 125) <= input(9);
output(0, 126) <= input(10);
output(0, 127) <= input(11);
output(0, 128) <= input(39);
output(0, 129) <= input(38);
output(0, 130) <= input(35);
output(0, 131) <= input(36);
output(0, 132) <= input(32);
output(0, 133) <= input(0);
output(0, 134) <= input(1);
output(0, 135) <= input(2);
output(0, 136) <= input(3);
output(0, 137) <= input(4);
output(0, 138) <= input(5);
output(0, 139) <= input(6);
output(0, 140) <= input(7);
output(0, 141) <= input(8);
output(0, 142) <= input(9);
output(0, 143) <= input(10);
output(0, 144) <= input(40);
output(0, 145) <= input(41);
output(0, 146) <= input(37);
output(0, 147) <= input(34);
output(0, 148) <= input(33);
output(0, 149) <= input(16);
output(0, 150) <= input(17);
output(0, 151) <= input(18);
output(0, 152) <= input(19);
output(0, 153) <= input(20);
output(0, 154) <= input(21);
output(0, 155) <= input(22);
output(0, 156) <= input(23);
output(0, 157) <= input(24);
output(0, 158) <= input(25);
output(0, 159) <= input(26);
output(0, 160) <= input(42);
output(0, 161) <= input(39);
output(0, 162) <= input(38);
output(0, 163) <= input(35);
output(0, 164) <= input(36);
output(0, 165) <= input(32);
output(0, 166) <= input(0);
output(0, 167) <= input(1);
output(0, 168) <= input(2);
output(0, 169) <= input(3);
output(0, 170) <= input(4);
output(0, 171) <= input(5);
output(0, 172) <= input(6);
output(0, 173) <= input(7);
output(0, 174) <= input(8);
output(0, 175) <= input(9);
output(0, 176) <= input(43);
output(0, 177) <= input(40);
output(0, 178) <= input(41);
output(0, 179) <= input(37);
output(0, 180) <= input(34);
output(0, 181) <= input(33);
output(0, 182) <= input(16);
output(0, 183) <= input(17);
output(0, 184) <= input(18);
output(0, 185) <= input(19);
output(0, 186) <= input(20);
output(0, 187) <= input(21);
output(0, 188) <= input(22);
output(0, 189) <= input(23);
output(0, 190) <= input(24);
output(0, 191) <= input(25);
output(0, 192) <= input(44);
output(0, 193) <= input(43);
output(0, 194) <= input(40);
output(0, 195) <= input(41);
output(0, 196) <= input(37);
output(0, 197) <= input(34);
output(0, 198) <= input(33);
output(0, 199) <= input(16);
output(0, 200) <= input(17);
output(0, 201) <= input(18);
output(0, 202) <= input(19);
output(0, 203) <= input(20);
output(0, 204) <= input(21);
output(0, 205) <= input(22);
output(0, 206) <= input(23);
output(0, 207) <= input(24);
output(0, 208) <= input(45);
output(0, 209) <= input(46);
output(0, 210) <= input(42);
output(0, 211) <= input(39);
output(0, 212) <= input(38);
output(0, 213) <= input(35);
output(0, 214) <= input(36);
output(0, 215) <= input(32);
output(0, 216) <= input(0);
output(0, 217) <= input(1);
output(0, 218) <= input(2);
output(0, 219) <= input(3);
output(0, 220) <= input(4);
output(0, 221) <= input(5);
output(0, 222) <= input(6);
output(0, 223) <= input(7);
output(0, 224) <= input(47);
output(0, 225) <= input(44);
output(0, 226) <= input(43);
output(0, 227) <= input(40);
output(0, 228) <= input(41);
output(0, 229) <= input(37);
output(0, 230) <= input(34);
output(0, 231) <= input(33);
output(0, 232) <= input(16);
output(0, 233) <= input(17);
output(0, 234) <= input(18);
output(0, 235) <= input(19);
output(0, 236) <= input(20);
output(0, 237) <= input(21);
output(0, 238) <= input(22);
output(0, 239) <= input(23);
output(0, 240) <= input(48);
output(0, 241) <= input(45);
output(0, 242) <= input(46);
output(0, 243) <= input(42);
output(0, 244) <= input(39);
output(0, 245) <= input(38);
output(0, 246) <= input(35);
output(0, 247) <= input(36);
output(0, 248) <= input(32);
output(0, 249) <= input(0);
output(0, 250) <= input(1);
output(0, 251) <= input(2);
output(0, 252) <= input(3);
output(0, 253) <= input(4);
output(0, 254) <= input(5);
output(0, 255) <= input(6);
output(1, 0) <= input(0);
output(1, 1) <= input(1);
output(1, 2) <= input(2);
output(1, 3) <= input(3);
output(1, 4) <= input(4);
output(1, 5) <= input(5);
output(1, 6) <= input(6);
output(1, 7) <= input(7);
output(1, 8) <= input(8);
output(1, 9) <= input(9);
output(1, 10) <= input(10);
output(1, 11) <= input(11);
output(1, 12) <= input(12);
output(1, 13) <= input(13);
output(1, 14) <= input(14);
output(1, 15) <= input(15);
output(1, 16) <= input(16);
output(1, 17) <= input(17);
output(1, 18) <= input(18);
output(1, 19) <= input(19);
output(1, 20) <= input(20);
output(1, 21) <= input(21);
output(1, 22) <= input(22);
output(1, 23) <= input(23);
output(1, 24) <= input(24);
output(1, 25) <= input(25);
output(1, 26) <= input(26);
output(1, 27) <= input(27);
output(1, 28) <= input(28);
output(1, 29) <= input(29);
output(1, 30) <= input(30);
output(1, 31) <= input(31);
output(1, 32) <= input(33);
output(1, 33) <= input(16);
output(1, 34) <= input(17);
output(1, 35) <= input(18);
output(1, 36) <= input(19);
output(1, 37) <= input(20);
output(1, 38) <= input(21);
output(1, 39) <= input(22);
output(1, 40) <= input(23);
output(1, 41) <= input(24);
output(1, 42) <= input(25);
output(1, 43) <= input(26);
output(1, 44) <= input(27);
output(1, 45) <= input(28);
output(1, 46) <= input(29);
output(1, 47) <= input(30);
output(1, 48) <= input(36);
output(1, 49) <= input(32);
output(1, 50) <= input(0);
output(1, 51) <= input(1);
output(1, 52) <= input(2);
output(1, 53) <= input(3);
output(1, 54) <= input(4);
output(1, 55) <= input(5);
output(1, 56) <= input(6);
output(1, 57) <= input(7);
output(1, 58) <= input(8);
output(1, 59) <= input(9);
output(1, 60) <= input(10);
output(1, 61) <= input(11);
output(1, 62) <= input(12);
output(1, 63) <= input(13);
output(1, 64) <= input(35);
output(1, 65) <= input(36);
output(1, 66) <= input(32);
output(1, 67) <= input(0);
output(1, 68) <= input(1);
output(1, 69) <= input(2);
output(1, 70) <= input(3);
output(1, 71) <= input(4);
output(1, 72) <= input(5);
output(1, 73) <= input(6);
output(1, 74) <= input(7);
output(1, 75) <= input(8);
output(1, 76) <= input(9);
output(1, 77) <= input(10);
output(1, 78) <= input(11);
output(1, 79) <= input(12);
output(1, 80) <= input(37);
output(1, 81) <= input(34);
output(1, 82) <= input(33);
output(1, 83) <= input(16);
output(1, 84) <= input(17);
output(1, 85) <= input(18);
output(1, 86) <= input(19);
output(1, 87) <= input(20);
output(1, 88) <= input(21);
output(1, 89) <= input(22);
output(1, 90) <= input(23);
output(1, 91) <= input(24);
output(1, 92) <= input(25);
output(1, 93) <= input(26);
output(1, 94) <= input(27);
output(1, 95) <= input(28);
output(1, 96) <= input(41);
output(1, 97) <= input(37);
output(1, 98) <= input(34);
output(1, 99) <= input(33);
output(1, 100) <= input(16);
output(1, 101) <= input(17);
output(1, 102) <= input(18);
output(1, 103) <= input(19);
output(1, 104) <= input(20);
output(1, 105) <= input(21);
output(1, 106) <= input(22);
output(1, 107) <= input(23);
output(1, 108) <= input(24);
output(1, 109) <= input(25);
output(1, 110) <= input(26);
output(1, 111) <= input(27);
output(1, 112) <= input(39);
output(1, 113) <= input(38);
output(1, 114) <= input(35);
output(1, 115) <= input(36);
output(1, 116) <= input(32);
output(1, 117) <= input(0);
output(1, 118) <= input(1);
output(1, 119) <= input(2);
output(1, 120) <= input(3);
output(1, 121) <= input(4);
output(1, 122) <= input(5);
output(1, 123) <= input(6);
output(1, 124) <= input(7);
output(1, 125) <= input(8);
output(1, 126) <= input(9);
output(1, 127) <= input(10);
output(1, 128) <= input(40);
output(1, 129) <= input(41);
output(1, 130) <= input(37);
output(1, 131) <= input(34);
output(1, 132) <= input(33);
output(1, 133) <= input(16);
output(1, 134) <= input(17);
output(1, 135) <= input(18);
output(1, 136) <= input(19);
output(1, 137) <= input(20);
output(1, 138) <= input(21);
output(1, 139) <= input(22);
output(1, 140) <= input(23);
output(1, 141) <= input(24);
output(1, 142) <= input(25);
output(1, 143) <= input(26);
output(1, 144) <= input(43);
output(1, 145) <= input(40);
output(1, 146) <= input(41);
output(1, 147) <= input(37);
output(1, 148) <= input(34);
output(1, 149) <= input(33);
output(1, 150) <= input(16);
output(1, 151) <= input(17);
output(1, 152) <= input(18);
output(1, 153) <= input(19);
output(1, 154) <= input(20);
output(1, 155) <= input(21);
output(1, 156) <= input(22);
output(1, 157) <= input(23);
output(1, 158) <= input(24);
output(1, 159) <= input(25);
output(1, 160) <= input(46);
output(1, 161) <= input(42);
output(1, 162) <= input(39);
output(1, 163) <= input(38);
output(1, 164) <= input(35);
output(1, 165) <= input(36);
output(1, 166) <= input(32);
output(1, 167) <= input(0);
output(1, 168) <= input(1);
output(1, 169) <= input(2);
output(1, 170) <= input(3);
output(1, 171) <= input(4);
output(1, 172) <= input(5);
output(1, 173) <= input(6);
output(1, 174) <= input(7);
output(1, 175) <= input(8);
output(1, 176) <= input(45);
output(1, 177) <= input(46);
output(1, 178) <= input(42);
output(1, 179) <= input(39);
output(1, 180) <= input(38);
output(1, 181) <= input(35);
output(1, 182) <= input(36);
output(1, 183) <= input(32);
output(1, 184) <= input(0);
output(1, 185) <= input(1);
output(1, 186) <= input(2);
output(1, 187) <= input(3);
output(1, 188) <= input(4);
output(1, 189) <= input(5);
output(1, 190) <= input(6);
output(1, 191) <= input(7);
output(1, 192) <= input(47);
output(1, 193) <= input(44);
output(1, 194) <= input(43);
output(1, 195) <= input(40);
output(1, 196) <= input(41);
output(1, 197) <= input(37);
output(1, 198) <= input(34);
output(1, 199) <= input(33);
output(1, 200) <= input(16);
output(1, 201) <= input(17);
output(1, 202) <= input(18);
output(1, 203) <= input(19);
output(1, 204) <= input(20);
output(1, 205) <= input(21);
output(1, 206) <= input(22);
output(1, 207) <= input(23);
output(1, 208) <= input(49);
output(1, 209) <= input(47);
output(1, 210) <= input(44);
output(1, 211) <= input(43);
output(1, 212) <= input(40);
output(1, 213) <= input(41);
output(1, 214) <= input(37);
output(1, 215) <= input(34);
output(1, 216) <= input(33);
output(1, 217) <= input(16);
output(1, 218) <= input(17);
output(1, 219) <= input(18);
output(1, 220) <= input(19);
output(1, 221) <= input(20);
output(1, 222) <= input(21);
output(1, 223) <= input(22);
output(1, 224) <= input(50);
output(1, 225) <= input(48);
output(1, 226) <= input(45);
output(1, 227) <= input(46);
output(1, 228) <= input(42);
output(1, 229) <= input(39);
output(1, 230) <= input(38);
output(1, 231) <= input(35);
output(1, 232) <= input(36);
output(1, 233) <= input(32);
output(1, 234) <= input(0);
output(1, 235) <= input(1);
output(1, 236) <= input(2);
output(1, 237) <= input(3);
output(1, 238) <= input(4);
output(1, 239) <= input(5);
output(1, 240) <= input(51);
output(1, 241) <= input(49);
output(1, 242) <= input(47);
output(1, 243) <= input(44);
output(1, 244) <= input(43);
output(1, 245) <= input(40);
output(1, 246) <= input(41);
output(1, 247) <= input(37);
output(1, 248) <= input(34);
output(1, 249) <= input(33);
output(1, 250) <= input(16);
output(1, 251) <= input(17);
output(1, 252) <= input(18);
output(1, 253) <= input(19);
output(1, 254) <= input(20);
output(1, 255) <= input(21);
output(2, 0) <= input(0);
output(2, 1) <= input(1);
output(2, 2) <= input(2);
output(2, 3) <= input(3);
output(2, 4) <= input(4);
output(2, 5) <= input(5);
output(2, 6) <= input(6);
output(2, 7) <= input(7);
output(2, 8) <= input(8);
output(2, 9) <= input(9);
output(2, 10) <= input(10);
output(2, 11) <= input(11);
output(2, 12) <= input(12);
output(2, 13) <= input(13);
output(2, 14) <= input(14);
output(2, 15) <= input(15);
output(2, 16) <= input(32);
output(2, 17) <= input(0);
output(2, 18) <= input(1);
output(2, 19) <= input(2);
output(2, 20) <= input(3);
output(2, 21) <= input(4);
output(2, 22) <= input(5);
output(2, 23) <= input(6);
output(2, 24) <= input(7);
output(2, 25) <= input(8);
output(2, 26) <= input(9);
output(2, 27) <= input(10);
output(2, 28) <= input(11);
output(2, 29) <= input(12);
output(2, 30) <= input(13);
output(2, 31) <= input(14);
output(2, 32) <= input(33);
output(2, 33) <= input(16);
output(2, 34) <= input(17);
output(2, 35) <= input(18);
output(2, 36) <= input(19);
output(2, 37) <= input(20);
output(2, 38) <= input(21);
output(2, 39) <= input(22);
output(2, 40) <= input(23);
output(2, 41) <= input(24);
output(2, 42) <= input(25);
output(2, 43) <= input(26);
output(2, 44) <= input(27);
output(2, 45) <= input(28);
output(2, 46) <= input(29);
output(2, 47) <= input(30);
output(2, 48) <= input(34);
output(2, 49) <= input(33);
output(2, 50) <= input(16);
output(2, 51) <= input(17);
output(2, 52) <= input(18);
output(2, 53) <= input(19);
output(2, 54) <= input(20);
output(2, 55) <= input(21);
output(2, 56) <= input(22);
output(2, 57) <= input(23);
output(2, 58) <= input(24);
output(2, 59) <= input(25);
output(2, 60) <= input(26);
output(2, 61) <= input(27);
output(2, 62) <= input(28);
output(2, 63) <= input(29);
output(2, 64) <= input(37);
output(2, 65) <= input(34);
output(2, 66) <= input(33);
output(2, 67) <= input(16);
output(2, 68) <= input(17);
output(2, 69) <= input(18);
output(2, 70) <= input(19);
output(2, 71) <= input(20);
output(2, 72) <= input(21);
output(2, 73) <= input(22);
output(2, 74) <= input(23);
output(2, 75) <= input(24);
output(2, 76) <= input(25);
output(2, 77) <= input(26);
output(2, 78) <= input(27);
output(2, 79) <= input(28);
output(2, 80) <= input(38);
output(2, 81) <= input(35);
output(2, 82) <= input(36);
output(2, 83) <= input(32);
output(2, 84) <= input(0);
output(2, 85) <= input(1);
output(2, 86) <= input(2);
output(2, 87) <= input(3);
output(2, 88) <= input(4);
output(2, 89) <= input(5);
output(2, 90) <= input(6);
output(2, 91) <= input(7);
output(2, 92) <= input(8);
output(2, 93) <= input(9);
output(2, 94) <= input(10);
output(2, 95) <= input(11);
output(2, 96) <= input(39);
output(2, 97) <= input(38);
output(2, 98) <= input(35);
output(2, 99) <= input(36);
output(2, 100) <= input(32);
output(2, 101) <= input(0);
output(2, 102) <= input(1);
output(2, 103) <= input(2);
output(2, 104) <= input(3);
output(2, 105) <= input(4);
output(2, 106) <= input(5);
output(2, 107) <= input(6);
output(2, 108) <= input(7);
output(2, 109) <= input(8);
output(2, 110) <= input(9);
output(2, 111) <= input(10);
output(2, 112) <= input(40);
output(2, 113) <= input(41);
output(2, 114) <= input(37);
output(2, 115) <= input(34);
output(2, 116) <= input(33);
output(2, 117) <= input(16);
output(2, 118) <= input(17);
output(2, 119) <= input(18);
output(2, 120) <= input(19);
output(2, 121) <= input(20);
output(2, 122) <= input(21);
output(2, 123) <= input(22);
output(2, 124) <= input(23);
output(2, 125) <= input(24);
output(2, 126) <= input(25);
output(2, 127) <= input(26);
output(2, 128) <= input(43);
output(2, 129) <= input(40);
output(2, 130) <= input(41);
output(2, 131) <= input(37);
output(2, 132) <= input(34);
output(2, 133) <= input(33);
output(2, 134) <= input(16);
output(2, 135) <= input(17);
output(2, 136) <= input(18);
output(2, 137) <= input(19);
output(2, 138) <= input(20);
output(2, 139) <= input(21);
output(2, 140) <= input(22);
output(2, 141) <= input(23);
output(2, 142) <= input(24);
output(2, 143) <= input(25);
output(2, 144) <= input(44);
output(2, 145) <= input(43);
output(2, 146) <= input(40);
output(2, 147) <= input(41);
output(2, 148) <= input(37);
output(2, 149) <= input(34);
output(2, 150) <= input(33);
output(2, 151) <= input(16);
output(2, 152) <= input(17);
output(2, 153) <= input(18);
output(2, 154) <= input(19);
output(2, 155) <= input(20);
output(2, 156) <= input(21);
output(2, 157) <= input(22);
output(2, 158) <= input(23);
output(2, 159) <= input(24);
output(2, 160) <= input(45);
output(2, 161) <= input(46);
output(2, 162) <= input(42);
output(2, 163) <= input(39);
output(2, 164) <= input(38);
output(2, 165) <= input(35);
output(2, 166) <= input(36);
output(2, 167) <= input(32);
output(2, 168) <= input(0);
output(2, 169) <= input(1);
output(2, 170) <= input(2);
output(2, 171) <= input(3);
output(2, 172) <= input(4);
output(2, 173) <= input(5);
output(2, 174) <= input(6);
output(2, 175) <= input(7);
output(2, 176) <= input(48);
output(2, 177) <= input(45);
output(2, 178) <= input(46);
output(2, 179) <= input(42);
output(2, 180) <= input(39);
output(2, 181) <= input(38);
output(2, 182) <= input(35);
output(2, 183) <= input(36);
output(2, 184) <= input(32);
output(2, 185) <= input(0);
output(2, 186) <= input(1);
output(2, 187) <= input(2);
output(2, 188) <= input(3);
output(2, 189) <= input(4);
output(2, 190) <= input(5);
output(2, 191) <= input(6);
output(2, 192) <= input(50);
output(2, 193) <= input(48);
output(2, 194) <= input(45);
output(2, 195) <= input(46);
output(2, 196) <= input(42);
output(2, 197) <= input(39);
output(2, 198) <= input(38);
output(2, 199) <= input(35);
output(2, 200) <= input(36);
output(2, 201) <= input(32);
output(2, 202) <= input(0);
output(2, 203) <= input(1);
output(2, 204) <= input(2);
output(2, 205) <= input(3);
output(2, 206) <= input(4);
output(2, 207) <= input(5);
output(2, 208) <= input(51);
output(2, 209) <= input(49);
output(2, 210) <= input(47);
output(2, 211) <= input(44);
output(2, 212) <= input(43);
output(2, 213) <= input(40);
output(2, 214) <= input(41);
output(2, 215) <= input(37);
output(2, 216) <= input(34);
output(2, 217) <= input(33);
output(2, 218) <= input(16);
output(2, 219) <= input(17);
output(2, 220) <= input(18);
output(2, 221) <= input(19);
output(2, 222) <= input(20);
output(2, 223) <= input(21);
output(2, 224) <= input(52);
output(2, 225) <= input(51);
output(2, 226) <= input(49);
output(2, 227) <= input(47);
output(2, 228) <= input(44);
output(2, 229) <= input(43);
output(2, 230) <= input(40);
output(2, 231) <= input(41);
output(2, 232) <= input(37);
output(2, 233) <= input(34);
output(2, 234) <= input(33);
output(2, 235) <= input(16);
output(2, 236) <= input(17);
output(2, 237) <= input(18);
output(2, 238) <= input(19);
output(2, 239) <= input(20);
output(2, 240) <= input(53);
output(2, 241) <= input(54);
output(2, 242) <= input(50);
output(2, 243) <= input(48);
output(2, 244) <= input(45);
output(2, 245) <= input(46);
output(2, 246) <= input(42);
output(2, 247) <= input(39);
output(2, 248) <= input(38);
output(2, 249) <= input(35);
output(2, 250) <= input(36);
output(2, 251) <= input(32);
output(2, 252) <= input(0);
output(2, 253) <= input(1);
output(2, 254) <= input(2);
output(2, 255) <= input(3);
when "0111" =>
output(0, 0) <= input(0);
output(0, 1) <= input(1);
output(0, 2) <= input(2);
output(0, 3) <= input(3);
output(0, 4) <= input(4);
output(0, 5) <= input(5);
output(0, 6) <= input(6);
output(0, 7) <= input(7);
output(0, 8) <= input(8);
output(0, 9) <= input(9);
output(0, 10) <= input(10);
output(0, 11) <= input(11);
output(0, 12) <= input(12);
output(0, 13) <= input(13);
output(0, 14) <= input(14);
output(0, 15) <= input(15);
output(0, 16) <= input(16);
output(0, 17) <= input(0);
output(0, 18) <= input(1);
output(0, 19) <= input(2);
output(0, 20) <= input(3);
output(0, 21) <= input(4);
output(0, 22) <= input(5);
output(0, 23) <= input(6);
output(0, 24) <= input(7);
output(0, 25) <= input(8);
output(0, 26) <= input(9);
output(0, 27) <= input(10);
output(0, 28) <= input(11);
output(0, 29) <= input(12);
output(0, 30) <= input(13);
output(0, 31) <= input(14);
output(0, 32) <= input(17);
output(0, 33) <= input(16);
output(0, 34) <= input(0);
output(0, 35) <= input(1);
output(0, 36) <= input(2);
output(0, 37) <= input(3);
output(0, 38) <= input(4);
output(0, 39) <= input(5);
output(0, 40) <= input(6);
output(0, 41) <= input(7);
output(0, 42) <= input(8);
output(0, 43) <= input(9);
output(0, 44) <= input(10);
output(0, 45) <= input(11);
output(0, 46) <= input(12);
output(0, 47) <= input(13);
output(0, 48) <= input(18);
output(0, 49) <= input(17);
output(0, 50) <= input(16);
output(0, 51) <= input(0);
output(0, 52) <= input(1);
output(0, 53) <= input(2);
output(0, 54) <= input(3);
output(0, 55) <= input(4);
output(0, 56) <= input(5);
output(0, 57) <= input(6);
output(0, 58) <= input(7);
output(0, 59) <= input(8);
output(0, 60) <= input(9);
output(0, 61) <= input(10);
output(0, 62) <= input(11);
output(0, 63) <= input(12);
output(0, 64) <= input(19);
output(0, 65) <= input(18);
output(0, 66) <= input(17);
output(0, 67) <= input(16);
output(0, 68) <= input(0);
output(0, 69) <= input(1);
output(0, 70) <= input(2);
output(0, 71) <= input(3);
output(0, 72) <= input(4);
output(0, 73) <= input(5);
output(0, 74) <= input(6);
output(0, 75) <= input(7);
output(0, 76) <= input(8);
output(0, 77) <= input(9);
output(0, 78) <= input(10);
output(0, 79) <= input(11);
output(0, 80) <= input(20);
output(0, 81) <= input(21);
output(0, 82) <= input(22);
output(0, 83) <= input(23);
output(0, 84) <= input(24);
output(0, 85) <= input(25);
output(0, 86) <= input(26);
output(0, 87) <= input(27);
output(0, 88) <= input(28);
output(0, 89) <= input(29);
output(0, 90) <= input(30);
output(0, 91) <= input(31);
output(0, 92) <= input(32);
output(0, 93) <= input(33);
output(0, 94) <= input(34);
output(0, 95) <= input(35);
output(0, 96) <= input(36);
output(0, 97) <= input(20);
output(0, 98) <= input(21);
output(0, 99) <= input(22);
output(0, 100) <= input(23);
output(0, 101) <= input(24);
output(0, 102) <= input(25);
output(0, 103) <= input(26);
output(0, 104) <= input(27);
output(0, 105) <= input(28);
output(0, 106) <= input(29);
output(0, 107) <= input(30);
output(0, 108) <= input(31);
output(0, 109) <= input(32);
output(0, 110) <= input(33);
output(0, 111) <= input(34);
output(0, 112) <= input(37);
output(0, 113) <= input(36);
output(0, 114) <= input(20);
output(0, 115) <= input(21);
output(0, 116) <= input(22);
output(0, 117) <= input(23);
output(0, 118) <= input(24);
output(0, 119) <= input(25);
output(0, 120) <= input(26);
output(0, 121) <= input(27);
output(0, 122) <= input(28);
output(0, 123) <= input(29);
output(0, 124) <= input(30);
output(0, 125) <= input(31);
output(0, 126) <= input(32);
output(0, 127) <= input(33);
output(0, 128) <= input(38);
output(0, 129) <= input(37);
output(0, 130) <= input(36);
output(0, 131) <= input(20);
output(0, 132) <= input(21);
output(0, 133) <= input(22);
output(0, 134) <= input(23);
output(0, 135) <= input(24);
output(0, 136) <= input(25);
output(0, 137) <= input(26);
output(0, 138) <= input(27);
output(0, 139) <= input(28);
output(0, 140) <= input(29);
output(0, 141) <= input(30);
output(0, 142) <= input(31);
output(0, 143) <= input(32);
output(0, 144) <= input(39);
output(0, 145) <= input(38);
output(0, 146) <= input(37);
output(0, 147) <= input(36);
output(0, 148) <= input(20);
output(0, 149) <= input(21);
output(0, 150) <= input(22);
output(0, 151) <= input(23);
output(0, 152) <= input(24);
output(0, 153) <= input(25);
output(0, 154) <= input(26);
output(0, 155) <= input(27);
output(0, 156) <= input(28);
output(0, 157) <= input(29);
output(0, 158) <= input(30);
output(0, 159) <= input(31);
output(0, 160) <= input(40);
output(0, 161) <= input(41);
output(0, 162) <= input(42);
output(0, 163) <= input(43);
output(0, 164) <= input(44);
output(0, 165) <= input(19);
output(0, 166) <= input(18);
output(0, 167) <= input(17);
output(0, 168) <= input(16);
output(0, 169) <= input(0);
output(0, 170) <= input(1);
output(0, 171) <= input(2);
output(0, 172) <= input(3);
output(0, 173) <= input(4);
output(0, 174) <= input(5);
output(0, 175) <= input(6);
output(0, 176) <= input(45);
output(0, 177) <= input(40);
output(0, 178) <= input(41);
output(0, 179) <= input(42);
output(0, 180) <= input(43);
output(0, 181) <= input(44);
output(0, 182) <= input(19);
output(0, 183) <= input(18);
output(0, 184) <= input(17);
output(0, 185) <= input(16);
output(0, 186) <= input(0);
output(0, 187) <= input(1);
output(0, 188) <= input(2);
output(0, 189) <= input(3);
output(0, 190) <= input(4);
output(0, 191) <= input(5);
output(0, 192) <= input(46);
output(0, 193) <= input(45);
output(0, 194) <= input(40);
output(0, 195) <= input(41);
output(0, 196) <= input(42);
output(0, 197) <= input(43);
output(0, 198) <= input(44);
output(0, 199) <= input(19);
output(0, 200) <= input(18);
output(0, 201) <= input(17);
output(0, 202) <= input(16);
output(0, 203) <= input(0);
output(0, 204) <= input(1);
output(0, 205) <= input(2);
output(0, 206) <= input(3);
output(0, 207) <= input(4);
output(0, 208) <= input(47);
output(0, 209) <= input(46);
output(0, 210) <= input(45);
output(0, 211) <= input(40);
output(0, 212) <= input(41);
output(0, 213) <= input(42);
output(0, 214) <= input(43);
output(0, 215) <= input(44);
output(0, 216) <= input(19);
output(0, 217) <= input(18);
output(0, 218) <= input(17);
output(0, 219) <= input(16);
output(0, 220) <= input(0);
output(0, 221) <= input(1);
output(0, 222) <= input(2);
output(0, 223) <= input(3);
output(0, 224) <= input(48);
output(0, 225) <= input(47);
output(0, 226) <= input(46);
output(0, 227) <= input(45);
output(0, 228) <= input(40);
output(0, 229) <= input(41);
output(0, 230) <= input(42);
output(0, 231) <= input(43);
output(0, 232) <= input(44);
output(0, 233) <= input(19);
output(0, 234) <= input(18);
output(0, 235) <= input(17);
output(0, 236) <= input(16);
output(0, 237) <= input(0);
output(0, 238) <= input(1);
output(0, 239) <= input(2);
output(0, 240) <= input(49);
output(0, 241) <= input(50);
output(0, 242) <= input(51);
output(0, 243) <= input(52);
output(0, 244) <= input(53);
output(0, 245) <= input(39);
output(0, 246) <= input(38);
output(0, 247) <= input(37);
output(0, 248) <= input(36);
output(0, 249) <= input(20);
output(0, 250) <= input(21);
output(0, 251) <= input(22);
output(0, 252) <= input(23);
output(0, 253) <= input(24);
output(0, 254) <= input(25);
output(0, 255) <= input(26);
output(1, 0) <= input(54);
output(1, 1) <= input(55);
output(1, 2) <= input(56);
output(1, 3) <= input(57);
output(1, 4) <= input(58);
output(1, 5) <= input(59);
output(1, 6) <= input(60);
output(1, 7) <= input(61);
output(1, 8) <= input(62);
output(1, 9) <= input(63);
output(1, 10) <= input(64);
output(1, 11) <= input(65);
output(1, 12) <= input(66);
output(1, 13) <= input(67);
output(1, 14) <= input(68);
output(1, 15) <= input(69);
output(1, 16) <= input(70);
output(1, 17) <= input(54);
output(1, 18) <= input(55);
output(1, 19) <= input(56);
output(1, 20) <= input(57);
output(1, 21) <= input(58);
output(1, 22) <= input(59);
output(1, 23) <= input(60);
output(1, 24) <= input(61);
output(1, 25) <= input(62);
output(1, 26) <= input(63);
output(1, 27) <= input(64);
output(1, 28) <= input(65);
output(1, 29) <= input(66);
output(1, 30) <= input(67);
output(1, 31) <= input(68);
output(1, 32) <= input(71);
output(1, 33) <= input(70);
output(1, 34) <= input(54);
output(1, 35) <= input(55);
output(1, 36) <= input(56);
output(1, 37) <= input(57);
output(1, 38) <= input(58);
output(1, 39) <= input(59);
output(1, 40) <= input(60);
output(1, 41) <= input(61);
output(1, 42) <= input(62);
output(1, 43) <= input(63);
output(1, 44) <= input(64);
output(1, 45) <= input(65);
output(1, 46) <= input(66);
output(1, 47) <= input(67);
output(1, 48) <= input(72);
output(1, 49) <= input(71);
output(1, 50) <= input(70);
output(1, 51) <= input(54);
output(1, 52) <= input(55);
output(1, 53) <= input(56);
output(1, 54) <= input(57);
output(1, 55) <= input(58);
output(1, 56) <= input(59);
output(1, 57) <= input(60);
output(1, 58) <= input(61);
output(1, 59) <= input(62);
output(1, 60) <= input(63);
output(1, 61) <= input(64);
output(1, 62) <= input(65);
output(1, 63) <= input(66);
output(1, 64) <= input(73);
output(1, 65) <= input(72);
output(1, 66) <= input(71);
output(1, 67) <= input(70);
output(1, 68) <= input(54);
output(1, 69) <= input(55);
output(1, 70) <= input(56);
output(1, 71) <= input(57);
output(1, 72) <= input(58);
output(1, 73) <= input(59);
output(1, 74) <= input(60);
output(1, 75) <= input(61);
output(1, 76) <= input(62);
output(1, 77) <= input(63);
output(1, 78) <= input(64);
output(1, 79) <= input(65);
output(1, 80) <= input(74);
output(1, 81) <= input(73);
output(1, 82) <= input(72);
output(1, 83) <= input(71);
output(1, 84) <= input(70);
output(1, 85) <= input(54);
output(1, 86) <= input(55);
output(1, 87) <= input(56);
output(1, 88) <= input(57);
output(1, 89) <= input(58);
output(1, 90) <= input(59);
output(1, 91) <= input(60);
output(1, 92) <= input(61);
output(1, 93) <= input(62);
output(1, 94) <= input(63);
output(1, 95) <= input(64);
output(1, 96) <= input(75);
output(1, 97) <= input(74);
output(1, 98) <= input(73);
output(1, 99) <= input(72);
output(1, 100) <= input(71);
output(1, 101) <= input(70);
output(1, 102) <= input(54);
output(1, 103) <= input(55);
output(1, 104) <= input(56);
output(1, 105) <= input(57);
output(1, 106) <= input(58);
output(1, 107) <= input(59);
output(1, 108) <= input(60);
output(1, 109) <= input(61);
output(1, 110) <= input(62);
output(1, 111) <= input(63);
output(1, 112) <= input(76);
output(1, 113) <= input(75);
output(1, 114) <= input(74);
output(1, 115) <= input(73);
output(1, 116) <= input(72);
output(1, 117) <= input(71);
output(1, 118) <= input(70);
output(1, 119) <= input(54);
output(1, 120) <= input(55);
output(1, 121) <= input(56);
output(1, 122) <= input(57);
output(1, 123) <= input(58);
output(1, 124) <= input(59);
output(1, 125) <= input(60);
output(1, 126) <= input(61);
output(1, 127) <= input(62);
output(1, 128) <= input(77);
output(1, 129) <= input(76);
output(1, 130) <= input(75);
output(1, 131) <= input(74);
output(1, 132) <= input(73);
output(1, 133) <= input(72);
output(1, 134) <= input(71);
output(1, 135) <= input(70);
output(1, 136) <= input(54);
output(1, 137) <= input(55);
output(1, 138) <= input(56);
output(1, 139) <= input(57);
output(1, 140) <= input(58);
output(1, 141) <= input(59);
output(1, 142) <= input(60);
output(1, 143) <= input(61);
output(1, 144) <= input(78);
output(1, 145) <= input(77);
output(1, 146) <= input(76);
output(1, 147) <= input(75);
output(1, 148) <= input(74);
output(1, 149) <= input(73);
output(1, 150) <= input(72);
output(1, 151) <= input(71);
output(1, 152) <= input(70);
output(1, 153) <= input(54);
output(1, 154) <= input(55);
output(1, 155) <= input(56);
output(1, 156) <= input(57);
output(1, 157) <= input(58);
output(1, 158) <= input(59);
output(1, 159) <= input(60);
output(1, 160) <= input(79);
output(1, 161) <= input(78);
output(1, 162) <= input(77);
output(1, 163) <= input(76);
output(1, 164) <= input(75);
output(1, 165) <= input(74);
output(1, 166) <= input(73);
output(1, 167) <= input(72);
output(1, 168) <= input(71);
output(1, 169) <= input(70);
output(1, 170) <= input(54);
output(1, 171) <= input(55);
output(1, 172) <= input(56);
output(1, 173) <= input(57);
output(1, 174) <= input(58);
output(1, 175) <= input(59);
output(1, 176) <= input(80);
output(1, 177) <= input(79);
output(1, 178) <= input(78);
output(1, 179) <= input(77);
output(1, 180) <= input(76);
output(1, 181) <= input(75);
output(1, 182) <= input(74);
output(1, 183) <= input(73);
output(1, 184) <= input(72);
output(1, 185) <= input(71);
output(1, 186) <= input(70);
output(1, 187) <= input(54);
output(1, 188) <= input(55);
output(1, 189) <= input(56);
output(1, 190) <= input(57);
output(1, 191) <= input(58);
output(1, 192) <= input(81);
output(1, 193) <= input(80);
output(1, 194) <= input(79);
output(1, 195) <= input(78);
output(1, 196) <= input(77);
output(1, 197) <= input(76);
output(1, 198) <= input(75);
output(1, 199) <= input(74);
output(1, 200) <= input(73);
output(1, 201) <= input(72);
output(1, 202) <= input(71);
output(1, 203) <= input(70);
output(1, 204) <= input(54);
output(1, 205) <= input(55);
output(1, 206) <= input(56);
output(1, 207) <= input(57);
output(1, 208) <= input(82);
output(1, 209) <= input(81);
output(1, 210) <= input(80);
output(1, 211) <= input(79);
output(1, 212) <= input(78);
output(1, 213) <= input(77);
output(1, 214) <= input(76);
output(1, 215) <= input(75);
output(1, 216) <= input(74);
output(1, 217) <= input(73);
output(1, 218) <= input(72);
output(1, 219) <= input(71);
output(1, 220) <= input(70);
output(1, 221) <= input(54);
output(1, 222) <= input(55);
output(1, 223) <= input(56);
output(1, 224) <= input(83);
output(1, 225) <= input(82);
output(1, 226) <= input(81);
output(1, 227) <= input(80);
output(1, 228) <= input(79);
output(1, 229) <= input(78);
output(1, 230) <= input(77);
output(1, 231) <= input(76);
output(1, 232) <= input(75);
output(1, 233) <= input(74);
output(1, 234) <= input(73);
output(1, 235) <= input(72);
output(1, 236) <= input(71);
output(1, 237) <= input(70);
output(1, 238) <= input(54);
output(1, 239) <= input(55);
output(1, 240) <= input(84);
output(1, 241) <= input(83);
output(1, 242) <= input(82);
output(1, 243) <= input(81);
output(1, 244) <= input(80);
output(1, 245) <= input(79);
output(1, 246) <= input(78);
output(1, 247) <= input(77);
output(1, 248) <= input(76);
output(1, 249) <= input(75);
output(1, 250) <= input(74);
output(1, 251) <= input(73);
output(1, 252) <= input(72);
output(1, 253) <= input(71);
output(1, 254) <= input(70);
output(1, 255) <= input(54);
when "1000" =>
output(0, 0) <= input(0);
output(0, 1) <= input(1);
output(0, 2) <= input(2);
output(0, 3) <= input(3);
output(0, 4) <= input(4);
output(0, 5) <= input(5);
output(0, 6) <= input(6);
output(0, 7) <= input(7);
output(0, 8) <= input(8);
output(0, 9) <= input(9);
output(0, 10) <= input(10);
output(0, 11) <= input(11);
output(0, 12) <= input(12);
output(0, 13) <= input(13);
output(0, 14) <= input(14);
output(0, 15) <= input(15);
output(0, 16) <= input(16);
output(0, 17) <= input(0);
output(0, 18) <= input(1);
output(0, 19) <= input(2);
output(0, 20) <= input(3);
output(0, 21) <= input(4);
output(0, 22) <= input(5);
output(0, 23) <= input(6);
output(0, 24) <= input(7);
output(0, 25) <= input(8);
output(0, 26) <= input(9);
output(0, 27) <= input(10);
output(0, 28) <= input(11);
output(0, 29) <= input(12);
output(0, 30) <= input(13);
output(0, 31) <= input(14);
output(0, 32) <= input(17);
output(0, 33) <= input(16);
output(0, 34) <= input(0);
output(0, 35) <= input(1);
output(0, 36) <= input(2);
output(0, 37) <= input(3);
output(0, 38) <= input(4);
output(0, 39) <= input(5);
output(0, 40) <= input(6);
output(0, 41) <= input(7);
output(0, 42) <= input(8);
output(0, 43) <= input(9);
output(0, 44) <= input(10);
output(0, 45) <= input(11);
output(0, 46) <= input(12);
output(0, 47) <= input(13);
output(0, 48) <= input(18);
output(0, 49) <= input(17);
output(0, 50) <= input(16);
output(0, 51) <= input(0);
output(0, 52) <= input(1);
output(0, 53) <= input(2);
output(0, 54) <= input(3);
output(0, 55) <= input(4);
output(0, 56) <= input(5);
output(0, 57) <= input(6);
output(0, 58) <= input(7);
output(0, 59) <= input(8);
output(0, 60) <= input(9);
output(0, 61) <= input(10);
output(0, 62) <= input(11);
output(0, 63) <= input(12);
output(0, 64) <= input(19);
output(0, 65) <= input(18);
output(0, 66) <= input(17);
output(0, 67) <= input(16);
output(0, 68) <= input(0);
output(0, 69) <= input(1);
output(0, 70) <= input(2);
output(0, 71) <= input(3);
output(0, 72) <= input(4);
output(0, 73) <= input(5);
output(0, 74) <= input(6);
output(0, 75) <= input(7);
output(0, 76) <= input(8);
output(0, 77) <= input(9);
output(0, 78) <= input(10);
output(0, 79) <= input(11);
output(0, 80) <= input(20);
output(0, 81) <= input(21);
output(0, 82) <= input(22);
output(0, 83) <= input(23);
output(0, 84) <= input(24);
output(0, 85) <= input(25);
output(0, 86) <= input(26);
output(0, 87) <= input(27);
output(0, 88) <= input(28);
output(0, 89) <= input(29);
output(0, 90) <= input(30);
output(0, 91) <= input(31);
output(0, 92) <= input(32);
output(0, 93) <= input(33);
output(0, 94) <= input(34);
output(0, 95) <= input(35);
output(0, 96) <= input(36);
output(0, 97) <= input(20);
output(0, 98) <= input(21);
output(0, 99) <= input(22);
output(0, 100) <= input(23);
output(0, 101) <= input(24);
output(0, 102) <= input(25);
output(0, 103) <= input(26);
output(0, 104) <= input(27);
output(0, 105) <= input(28);
output(0, 106) <= input(29);
output(0, 107) <= input(30);
output(0, 108) <= input(31);
output(0, 109) <= input(32);
output(0, 110) <= input(33);
output(0, 111) <= input(34);
output(0, 112) <= input(37);
output(0, 113) <= input(36);
output(0, 114) <= input(20);
output(0, 115) <= input(21);
output(0, 116) <= input(22);
output(0, 117) <= input(23);
output(0, 118) <= input(24);
output(0, 119) <= input(25);
output(0, 120) <= input(26);
output(0, 121) <= input(27);
output(0, 122) <= input(28);
output(0, 123) <= input(29);
output(0, 124) <= input(30);
output(0, 125) <= input(31);
output(0, 126) <= input(32);
output(0, 127) <= input(33);
output(0, 128) <= input(38);
output(0, 129) <= input(37);
output(0, 130) <= input(36);
output(0, 131) <= input(20);
output(0, 132) <= input(21);
output(0, 133) <= input(22);
output(0, 134) <= input(23);
output(0, 135) <= input(24);
output(0, 136) <= input(25);
output(0, 137) <= input(26);
output(0, 138) <= input(27);
output(0, 139) <= input(28);
output(0, 140) <= input(29);
output(0, 141) <= input(30);
output(0, 142) <= input(31);
output(0, 143) <= input(32);
output(0, 144) <= input(39);
output(0, 145) <= input(38);
output(0, 146) <= input(37);
output(0, 147) <= input(36);
output(0, 148) <= input(20);
output(0, 149) <= input(21);
output(0, 150) <= input(22);
output(0, 151) <= input(23);
output(0, 152) <= input(24);
output(0, 153) <= input(25);
output(0, 154) <= input(26);
output(0, 155) <= input(27);
output(0, 156) <= input(28);
output(0, 157) <= input(29);
output(0, 158) <= input(30);
output(0, 159) <= input(31);
output(0, 160) <= input(40);
output(0, 161) <= input(41);
output(0, 162) <= input(42);
output(0, 163) <= input(43);
output(0, 164) <= input(44);
output(0, 165) <= input(19);
output(0, 166) <= input(18);
output(0, 167) <= input(17);
output(0, 168) <= input(16);
output(0, 169) <= input(0);
output(0, 170) <= input(1);
output(0, 171) <= input(2);
output(0, 172) <= input(3);
output(0, 173) <= input(4);
output(0, 174) <= input(5);
output(0, 175) <= input(6);
output(0, 176) <= input(45);
output(0, 177) <= input(40);
output(0, 178) <= input(41);
output(0, 179) <= input(42);
output(0, 180) <= input(43);
output(0, 181) <= input(44);
output(0, 182) <= input(19);
output(0, 183) <= input(18);
output(0, 184) <= input(17);
output(0, 185) <= input(16);
output(0, 186) <= input(0);
output(0, 187) <= input(1);
output(0, 188) <= input(2);
output(0, 189) <= input(3);
output(0, 190) <= input(4);
output(0, 191) <= input(5);
output(0, 192) <= input(46);
output(0, 193) <= input(45);
output(0, 194) <= input(40);
output(0, 195) <= input(41);
output(0, 196) <= input(42);
output(0, 197) <= input(43);
output(0, 198) <= input(44);
output(0, 199) <= input(19);
output(0, 200) <= input(18);
output(0, 201) <= input(17);
output(0, 202) <= input(16);
output(0, 203) <= input(0);
output(0, 204) <= input(1);
output(0, 205) <= input(2);
output(0, 206) <= input(3);
output(0, 207) <= input(4);
output(0, 208) <= input(47);
output(0, 209) <= input(46);
output(0, 210) <= input(45);
output(0, 211) <= input(40);
output(0, 212) <= input(41);
output(0, 213) <= input(42);
output(0, 214) <= input(43);
output(0, 215) <= input(44);
output(0, 216) <= input(19);
output(0, 217) <= input(18);
output(0, 218) <= input(17);
output(0, 219) <= input(16);
output(0, 220) <= input(0);
output(0, 221) <= input(1);
output(0, 222) <= input(2);
output(0, 223) <= input(3);
output(0, 224) <= input(48);
output(0, 225) <= input(47);
output(0, 226) <= input(46);
output(0, 227) <= input(45);
output(0, 228) <= input(40);
output(0, 229) <= input(41);
output(0, 230) <= input(42);
output(0, 231) <= input(43);
output(0, 232) <= input(44);
output(0, 233) <= input(19);
output(0, 234) <= input(18);
output(0, 235) <= input(17);
output(0, 236) <= input(16);
output(0, 237) <= input(0);
output(0, 238) <= input(1);
output(0, 239) <= input(2);
output(0, 240) <= input(49);
output(0, 241) <= input(50);
output(0, 242) <= input(51);
output(0, 243) <= input(52);
output(0, 244) <= input(53);
output(0, 245) <= input(39);
output(0, 246) <= input(38);
output(0, 247) <= input(37);
output(0, 248) <= input(36);
output(0, 249) <= input(20);
output(0, 250) <= input(21);
output(0, 251) <= input(22);
output(0, 252) <= input(23);
output(0, 253) <= input(24);
output(0, 254) <= input(25);
output(0, 255) <= input(26);
when "1001" =>
output(0, 0) <= input(0);
output(0, 1) <= input(1);
output(0, 2) <= input(2);
output(0, 3) <= input(3);
output(0, 4) <= input(4);
output(0, 5) <= input(5);
output(0, 6) <= input(6);
output(0, 7) <= input(7);
output(0, 8) <= input(8);
output(0, 9) <= input(9);
output(0, 10) <= input(10);
output(0, 11) <= input(11);
output(0, 12) <= input(12);
output(0, 13) <= input(13);
output(0, 14) <= input(14);
output(0, 15) <= input(15);
output(0, 16) <= input(16);
output(0, 17) <= input(0);
output(0, 18) <= input(1);
output(0, 19) <= input(2);
output(0, 20) <= input(3);
output(0, 21) <= input(4);
output(0, 22) <= input(5);
output(0, 23) <= input(6);
output(0, 24) <= input(7);
output(0, 25) <= input(8);
output(0, 26) <= input(9);
output(0, 27) <= input(10);
output(0, 28) <= input(11);
output(0, 29) <= input(12);
output(0, 30) <= input(13);
output(0, 31) <= input(14);
output(0, 32) <= input(17);
output(0, 33) <= input(18);
output(0, 34) <= input(19);
output(0, 35) <= input(20);
output(0, 36) <= input(21);
output(0, 37) <= input(22);
output(0, 38) <= input(23);
output(0, 39) <= input(24);
output(0, 40) <= input(25);
output(0, 41) <= input(26);
output(0, 42) <= input(27);
output(0, 43) <= input(28);
output(0, 44) <= input(29);
output(0, 45) <= input(30);
output(0, 46) <= input(31);
output(0, 47) <= input(32);
output(0, 48) <= input(33);
output(0, 49) <= input(17);
output(0, 50) <= input(18);
output(0, 51) <= input(19);
output(0, 52) <= input(20);
output(0, 53) <= input(21);
output(0, 54) <= input(22);
output(0, 55) <= input(23);
output(0, 56) <= input(24);
output(0, 57) <= input(25);
output(0, 58) <= input(26);
output(0, 59) <= input(27);
output(0, 60) <= input(28);
output(0, 61) <= input(29);
output(0, 62) <= input(30);
output(0, 63) <= input(31);
output(0, 64) <= input(34);
output(0, 65) <= input(33);
output(0, 66) <= input(17);
output(0, 67) <= input(18);
output(0, 68) <= input(19);
output(0, 69) <= input(20);
output(0, 70) <= input(21);
output(0, 71) <= input(22);
output(0, 72) <= input(23);
output(0, 73) <= input(24);
output(0, 74) <= input(25);
output(0, 75) <= input(26);
output(0, 76) <= input(27);
output(0, 77) <= input(28);
output(0, 78) <= input(29);
output(0, 79) <= input(30);
output(0, 80) <= input(35);
output(0, 81) <= input(36);
output(0, 82) <= input(37);
output(0, 83) <= input(16);
output(0, 84) <= input(0);
output(0, 85) <= input(1);
output(0, 86) <= input(2);
output(0, 87) <= input(3);
output(0, 88) <= input(4);
output(0, 89) <= input(5);
output(0, 90) <= input(6);
output(0, 91) <= input(7);
output(0, 92) <= input(8);
output(0, 93) <= input(9);
output(0, 94) <= input(10);
output(0, 95) <= input(11);
output(0, 96) <= input(38);
output(0, 97) <= input(35);
output(0, 98) <= input(36);
output(0, 99) <= input(37);
output(0, 100) <= input(16);
output(0, 101) <= input(0);
output(0, 102) <= input(1);
output(0, 103) <= input(2);
output(0, 104) <= input(3);
output(0, 105) <= input(4);
output(0, 106) <= input(5);
output(0, 107) <= input(6);
output(0, 108) <= input(7);
output(0, 109) <= input(8);
output(0, 110) <= input(9);
output(0, 111) <= input(10);
output(0, 112) <= input(39);
output(0, 113) <= input(40);
output(0, 114) <= input(34);
output(0, 115) <= input(33);
output(0, 116) <= input(17);
output(0, 117) <= input(18);
output(0, 118) <= input(19);
output(0, 119) <= input(20);
output(0, 120) <= input(21);
output(0, 121) <= input(22);
output(0, 122) <= input(23);
output(0, 123) <= input(24);
output(0, 124) <= input(25);
output(0, 125) <= input(26);
output(0, 126) <= input(27);
output(0, 127) <= input(28);
output(0, 128) <= input(41);
output(0, 129) <= input(39);
output(0, 130) <= input(40);
output(0, 131) <= input(34);
output(0, 132) <= input(33);
output(0, 133) <= input(17);
output(0, 134) <= input(18);
output(0, 135) <= input(19);
output(0, 136) <= input(20);
output(0, 137) <= input(21);
output(0, 138) <= input(22);
output(0, 139) <= input(23);
output(0, 140) <= input(24);
output(0, 141) <= input(25);
output(0, 142) <= input(26);
output(0, 143) <= input(27);
output(0, 144) <= input(42);
output(0, 145) <= input(41);
output(0, 146) <= input(39);
output(0, 147) <= input(40);
output(0, 148) <= input(34);
output(0, 149) <= input(33);
output(0, 150) <= input(17);
output(0, 151) <= input(18);
output(0, 152) <= input(19);
output(0, 153) <= input(20);
output(0, 154) <= input(21);
output(0, 155) <= input(22);
output(0, 156) <= input(23);
output(0, 157) <= input(24);
output(0, 158) <= input(25);
output(0, 159) <= input(26);
output(0, 160) <= input(43);
output(0, 161) <= input(44);
output(0, 162) <= input(45);
output(0, 163) <= input(38);
output(0, 164) <= input(35);
output(0, 165) <= input(36);
output(0, 166) <= input(37);
output(0, 167) <= input(16);
output(0, 168) <= input(0);
output(0, 169) <= input(1);
output(0, 170) <= input(2);
output(0, 171) <= input(3);
output(0, 172) <= input(4);
output(0, 173) <= input(5);
output(0, 174) <= input(6);
output(0, 175) <= input(7);
output(0, 176) <= input(46);
output(0, 177) <= input(43);
output(0, 178) <= input(44);
output(0, 179) <= input(45);
output(0, 180) <= input(38);
output(0, 181) <= input(35);
output(0, 182) <= input(36);
output(0, 183) <= input(37);
output(0, 184) <= input(16);
output(0, 185) <= input(0);
output(0, 186) <= input(1);
output(0, 187) <= input(2);
output(0, 188) <= input(3);
output(0, 189) <= input(4);
output(0, 190) <= input(5);
output(0, 191) <= input(6);
output(0, 192) <= input(47);
output(0, 193) <= input(46);
output(0, 194) <= input(43);
output(0, 195) <= input(44);
output(0, 196) <= input(45);
output(0, 197) <= input(38);
output(0, 198) <= input(35);
output(0, 199) <= input(36);
output(0, 200) <= input(37);
output(0, 201) <= input(16);
output(0, 202) <= input(0);
output(0, 203) <= input(1);
output(0, 204) <= input(2);
output(0, 205) <= input(3);
output(0, 206) <= input(4);
output(0, 207) <= input(5);
output(0, 208) <= input(48);
output(0, 209) <= input(49);
output(0, 210) <= input(50);
output(0, 211) <= input(42);
output(0, 212) <= input(41);
output(0, 213) <= input(39);
output(0, 214) <= input(40);
output(0, 215) <= input(34);
output(0, 216) <= input(33);
output(0, 217) <= input(17);
output(0, 218) <= input(18);
output(0, 219) <= input(19);
output(0, 220) <= input(20);
output(0, 221) <= input(21);
output(0, 222) <= input(22);
output(0, 223) <= input(23);
output(0, 224) <= input(51);
output(0, 225) <= input(48);
output(0, 226) <= input(49);
output(0, 227) <= input(50);
output(0, 228) <= input(42);
output(0, 229) <= input(41);
output(0, 230) <= input(39);
output(0, 231) <= input(40);
output(0, 232) <= input(34);
output(0, 233) <= input(33);
output(0, 234) <= input(17);
output(0, 235) <= input(18);
output(0, 236) <= input(19);
output(0, 237) <= input(20);
output(0, 238) <= input(21);
output(0, 239) <= input(22);
output(0, 240) <= input(52);
output(0, 241) <= input(53);
output(0, 242) <= input(47);
output(0, 243) <= input(46);
output(0, 244) <= input(43);
output(0, 245) <= input(44);
output(0, 246) <= input(45);
output(0, 247) <= input(38);
output(0, 248) <= input(35);
output(0, 249) <= input(36);
output(0, 250) <= input(37);
output(0, 251) <= input(16);
output(0, 252) <= input(0);
output(0, 253) <= input(1);
output(0, 254) <= input(2);
output(0, 255) <= input(3);
output(1, 0) <= input(0);
output(1, 1) <= input(1);
output(1, 2) <= input(2);
output(1, 3) <= input(3);
output(1, 4) <= input(4);
output(1, 5) <= input(5);
output(1, 6) <= input(6);
output(1, 7) <= input(7);
output(1, 8) <= input(8);
output(1, 9) <= input(9);
output(1, 10) <= input(10);
output(1, 11) <= input(11);
output(1, 12) <= input(12);
output(1, 13) <= input(13);
output(1, 14) <= input(14);
output(1, 15) <= input(15);
output(1, 16) <= input(18);
output(1, 17) <= input(19);
output(1, 18) <= input(20);
output(1, 19) <= input(21);
output(1, 20) <= input(22);
output(1, 21) <= input(23);
output(1, 22) <= input(24);
output(1, 23) <= input(25);
output(1, 24) <= input(26);
output(1, 25) <= input(27);
output(1, 26) <= input(28);
output(1, 27) <= input(29);
output(1, 28) <= input(30);
output(1, 29) <= input(31);
output(1, 30) <= input(32);
output(1, 31) <= input(54);
output(1, 32) <= input(17);
output(1, 33) <= input(18);
output(1, 34) <= input(19);
output(1, 35) <= input(20);
output(1, 36) <= input(21);
output(1, 37) <= input(22);
output(1, 38) <= input(23);
output(1, 39) <= input(24);
output(1, 40) <= input(25);
output(1, 41) <= input(26);
output(1, 42) <= input(27);
output(1, 43) <= input(28);
output(1, 44) <= input(29);
output(1, 45) <= input(30);
output(1, 46) <= input(31);
output(1, 47) <= input(32);
output(1, 48) <= input(37);
output(1, 49) <= input(16);
output(1, 50) <= input(0);
output(1, 51) <= input(1);
output(1, 52) <= input(2);
output(1, 53) <= input(3);
output(1, 54) <= input(4);
output(1, 55) <= input(5);
output(1, 56) <= input(6);
output(1, 57) <= input(7);
output(1, 58) <= input(8);
output(1, 59) <= input(9);
output(1, 60) <= input(10);
output(1, 61) <= input(11);
output(1, 62) <= input(12);
output(1, 63) <= input(13);
output(1, 64) <= input(36);
output(1, 65) <= input(37);
output(1, 66) <= input(16);
output(1, 67) <= input(0);
output(1, 68) <= input(1);
output(1, 69) <= input(2);
output(1, 70) <= input(3);
output(1, 71) <= input(4);
output(1, 72) <= input(5);
output(1, 73) <= input(6);
output(1, 74) <= input(7);
output(1, 75) <= input(8);
output(1, 76) <= input(9);
output(1, 77) <= input(10);
output(1, 78) <= input(11);
output(1, 79) <= input(12);
output(1, 80) <= input(34);
output(1, 81) <= input(33);
output(1, 82) <= input(17);
output(1, 83) <= input(18);
output(1, 84) <= input(19);
output(1, 85) <= input(20);
output(1, 86) <= input(21);
output(1, 87) <= input(22);
output(1, 88) <= input(23);
output(1, 89) <= input(24);
output(1, 90) <= input(25);
output(1, 91) <= input(26);
output(1, 92) <= input(27);
output(1, 93) <= input(28);
output(1, 94) <= input(29);
output(1, 95) <= input(30);
output(1, 96) <= input(40);
output(1, 97) <= input(34);
output(1, 98) <= input(33);
output(1, 99) <= input(17);
output(1, 100) <= input(18);
output(1, 101) <= input(19);
output(1, 102) <= input(20);
output(1, 103) <= input(21);
output(1, 104) <= input(22);
output(1, 105) <= input(23);
output(1, 106) <= input(24);
output(1, 107) <= input(25);
output(1, 108) <= input(26);
output(1, 109) <= input(27);
output(1, 110) <= input(28);
output(1, 111) <= input(29);
output(1, 112) <= input(38);
output(1, 113) <= input(35);
output(1, 114) <= input(36);
output(1, 115) <= input(37);
output(1, 116) <= input(16);
output(1, 117) <= input(0);
output(1, 118) <= input(1);
output(1, 119) <= input(2);
output(1, 120) <= input(3);
output(1, 121) <= input(4);
output(1, 122) <= input(5);
output(1, 123) <= input(6);
output(1, 124) <= input(7);
output(1, 125) <= input(8);
output(1, 126) <= input(9);
output(1, 127) <= input(10);
output(1, 128) <= input(39);
output(1, 129) <= input(40);
output(1, 130) <= input(34);
output(1, 131) <= input(33);
output(1, 132) <= input(17);
output(1, 133) <= input(18);
output(1, 134) <= input(19);
output(1, 135) <= input(20);
output(1, 136) <= input(21);
output(1, 137) <= input(22);
output(1, 138) <= input(23);
output(1, 139) <= input(24);
output(1, 140) <= input(25);
output(1, 141) <= input(26);
output(1, 142) <= input(27);
output(1, 143) <= input(28);
output(1, 144) <= input(41);
output(1, 145) <= input(39);
output(1, 146) <= input(40);
output(1, 147) <= input(34);
output(1, 148) <= input(33);
output(1, 149) <= input(17);
output(1, 150) <= input(18);
output(1, 151) <= input(19);
output(1, 152) <= input(20);
output(1, 153) <= input(21);
output(1, 154) <= input(22);
output(1, 155) <= input(23);
output(1, 156) <= input(24);
output(1, 157) <= input(25);
output(1, 158) <= input(26);
output(1, 159) <= input(27);
output(1, 160) <= input(44);
output(1, 161) <= input(45);
output(1, 162) <= input(38);
output(1, 163) <= input(35);
output(1, 164) <= input(36);
output(1, 165) <= input(37);
output(1, 166) <= input(16);
output(1, 167) <= input(0);
output(1, 168) <= input(1);
output(1, 169) <= input(2);
output(1, 170) <= input(3);
output(1, 171) <= input(4);
output(1, 172) <= input(5);
output(1, 173) <= input(6);
output(1, 174) <= input(7);
output(1, 175) <= input(8);
output(1, 176) <= input(43);
output(1, 177) <= input(44);
output(1, 178) <= input(45);
output(1, 179) <= input(38);
output(1, 180) <= input(35);
output(1, 181) <= input(36);
output(1, 182) <= input(37);
output(1, 183) <= input(16);
output(1, 184) <= input(0);
output(1, 185) <= input(1);
output(1, 186) <= input(2);
output(1, 187) <= input(3);
output(1, 188) <= input(4);
output(1, 189) <= input(5);
output(1, 190) <= input(6);
output(1, 191) <= input(7);
output(1, 192) <= input(50);
output(1, 193) <= input(42);
output(1, 194) <= input(41);
output(1, 195) <= input(39);
output(1, 196) <= input(40);
output(1, 197) <= input(34);
output(1, 198) <= input(33);
output(1, 199) <= input(17);
output(1, 200) <= input(18);
output(1, 201) <= input(19);
output(1, 202) <= input(20);
output(1, 203) <= input(21);
output(1, 204) <= input(22);
output(1, 205) <= input(23);
output(1, 206) <= input(24);
output(1, 207) <= input(25);
output(1, 208) <= input(49);
output(1, 209) <= input(50);
output(1, 210) <= input(42);
output(1, 211) <= input(41);
output(1, 212) <= input(39);
output(1, 213) <= input(40);
output(1, 214) <= input(34);
output(1, 215) <= input(33);
output(1, 216) <= input(17);
output(1, 217) <= input(18);
output(1, 218) <= input(19);
output(1, 219) <= input(20);
output(1, 220) <= input(21);
output(1, 221) <= input(22);
output(1, 222) <= input(23);
output(1, 223) <= input(24);
output(1, 224) <= input(47);
output(1, 225) <= input(46);
output(1, 226) <= input(43);
output(1, 227) <= input(44);
output(1, 228) <= input(45);
output(1, 229) <= input(38);
output(1, 230) <= input(35);
output(1, 231) <= input(36);
output(1, 232) <= input(37);
output(1, 233) <= input(16);
output(1, 234) <= input(0);
output(1, 235) <= input(1);
output(1, 236) <= input(2);
output(1, 237) <= input(3);
output(1, 238) <= input(4);
output(1, 239) <= input(5);
output(1, 240) <= input(48);
output(1, 241) <= input(49);
output(1, 242) <= input(50);
output(1, 243) <= input(42);
output(1, 244) <= input(41);
output(1, 245) <= input(39);
output(1, 246) <= input(40);
output(1, 247) <= input(34);
output(1, 248) <= input(33);
output(1, 249) <= input(17);
output(1, 250) <= input(18);
output(1, 251) <= input(19);
output(1, 252) <= input(20);
output(1, 253) <= input(21);
output(1, 254) <= input(22);
output(1, 255) <= input(23);
output(2, 0) <= input(0);
output(2, 1) <= input(1);
output(2, 2) <= input(2);
output(2, 3) <= input(3);
output(2, 4) <= input(4);
output(2, 5) <= input(5);
output(2, 6) <= input(6);
output(2, 7) <= input(7);
output(2, 8) <= input(8);
output(2, 9) <= input(9);
output(2, 10) <= input(10);
output(2, 11) <= input(11);
output(2, 12) <= input(12);
output(2, 13) <= input(13);
output(2, 14) <= input(14);
output(2, 15) <= input(15);
output(2, 16) <= input(18);
output(2, 17) <= input(19);
output(2, 18) <= input(20);
output(2, 19) <= input(21);
output(2, 20) <= input(22);
output(2, 21) <= input(23);
output(2, 22) <= input(24);
output(2, 23) <= input(25);
output(2, 24) <= input(26);
output(2, 25) <= input(27);
output(2, 26) <= input(28);
output(2, 27) <= input(29);
output(2, 28) <= input(30);
output(2, 29) <= input(31);
output(2, 30) <= input(32);
output(2, 31) <= input(54);
output(2, 32) <= input(16);
output(2, 33) <= input(0);
output(2, 34) <= input(1);
output(2, 35) <= input(2);
output(2, 36) <= input(3);
output(2, 37) <= input(4);
output(2, 38) <= input(5);
output(2, 39) <= input(6);
output(2, 40) <= input(7);
output(2, 41) <= input(8);
output(2, 42) <= input(9);
output(2, 43) <= input(10);
output(2, 44) <= input(11);
output(2, 45) <= input(12);
output(2, 46) <= input(13);
output(2, 47) <= input(14);
output(2, 48) <= input(17);
output(2, 49) <= input(18);
output(2, 50) <= input(19);
output(2, 51) <= input(20);
output(2, 52) <= input(21);
output(2, 53) <= input(22);
output(2, 54) <= input(23);
output(2, 55) <= input(24);
output(2, 56) <= input(25);
output(2, 57) <= input(26);
output(2, 58) <= input(27);
output(2, 59) <= input(28);
output(2, 60) <= input(29);
output(2, 61) <= input(30);
output(2, 62) <= input(31);
output(2, 63) <= input(32);
output(2, 64) <= input(33);
output(2, 65) <= input(17);
output(2, 66) <= input(18);
output(2, 67) <= input(19);
output(2, 68) <= input(20);
output(2, 69) <= input(21);
output(2, 70) <= input(22);
output(2, 71) <= input(23);
output(2, 72) <= input(24);
output(2, 73) <= input(25);
output(2, 74) <= input(26);
output(2, 75) <= input(27);
output(2, 76) <= input(28);
output(2, 77) <= input(29);
output(2, 78) <= input(30);
output(2, 79) <= input(31);
output(2, 80) <= input(36);
output(2, 81) <= input(37);
output(2, 82) <= input(16);
output(2, 83) <= input(0);
output(2, 84) <= input(1);
output(2, 85) <= input(2);
output(2, 86) <= input(3);
output(2, 87) <= input(4);
output(2, 88) <= input(5);
output(2, 89) <= input(6);
output(2, 90) <= input(7);
output(2, 91) <= input(8);
output(2, 92) <= input(9);
output(2, 93) <= input(10);
output(2, 94) <= input(11);
output(2, 95) <= input(12);
output(2, 96) <= input(34);
output(2, 97) <= input(33);
output(2, 98) <= input(17);
output(2, 99) <= input(18);
output(2, 100) <= input(19);
output(2, 101) <= input(20);
output(2, 102) <= input(21);
output(2, 103) <= input(22);
output(2, 104) <= input(23);
output(2, 105) <= input(24);
output(2, 106) <= input(25);
output(2, 107) <= input(26);
output(2, 108) <= input(27);
output(2, 109) <= input(28);
output(2, 110) <= input(29);
output(2, 111) <= input(30);
output(2, 112) <= input(35);
output(2, 113) <= input(36);
output(2, 114) <= input(37);
output(2, 115) <= input(16);
output(2, 116) <= input(0);
output(2, 117) <= input(1);
output(2, 118) <= input(2);
output(2, 119) <= input(3);
output(2, 120) <= input(4);
output(2, 121) <= input(5);
output(2, 122) <= input(6);
output(2, 123) <= input(7);
output(2, 124) <= input(8);
output(2, 125) <= input(9);
output(2, 126) <= input(10);
output(2, 127) <= input(11);
output(2, 128) <= input(38);
output(2, 129) <= input(35);
output(2, 130) <= input(36);
output(2, 131) <= input(37);
output(2, 132) <= input(16);
output(2, 133) <= input(0);
output(2, 134) <= input(1);
output(2, 135) <= input(2);
output(2, 136) <= input(3);
output(2, 137) <= input(4);
output(2, 138) <= input(5);
output(2, 139) <= input(6);
output(2, 140) <= input(7);
output(2, 141) <= input(8);
output(2, 142) <= input(9);
output(2, 143) <= input(10);
output(2, 144) <= input(39);
output(2, 145) <= input(40);
output(2, 146) <= input(34);
output(2, 147) <= input(33);
output(2, 148) <= input(17);
output(2, 149) <= input(18);
output(2, 150) <= input(19);
output(2, 151) <= input(20);
output(2, 152) <= input(21);
output(2, 153) <= input(22);
output(2, 154) <= input(23);
output(2, 155) <= input(24);
output(2, 156) <= input(25);
output(2, 157) <= input(26);
output(2, 158) <= input(27);
output(2, 159) <= input(28);
output(2, 160) <= input(45);
output(2, 161) <= input(38);
output(2, 162) <= input(35);
output(2, 163) <= input(36);
output(2, 164) <= input(37);
output(2, 165) <= input(16);
output(2, 166) <= input(0);
output(2, 167) <= input(1);
output(2, 168) <= input(2);
output(2, 169) <= input(3);
output(2, 170) <= input(4);
output(2, 171) <= input(5);
output(2, 172) <= input(6);
output(2, 173) <= input(7);
output(2, 174) <= input(8);
output(2, 175) <= input(9);
output(2, 176) <= input(41);
output(2, 177) <= input(39);
output(2, 178) <= input(40);
output(2, 179) <= input(34);
output(2, 180) <= input(33);
output(2, 181) <= input(17);
output(2, 182) <= input(18);
output(2, 183) <= input(19);
output(2, 184) <= input(20);
output(2, 185) <= input(21);
output(2, 186) <= input(22);
output(2, 187) <= input(23);
output(2, 188) <= input(24);
output(2, 189) <= input(25);
output(2, 190) <= input(26);
output(2, 191) <= input(27);
output(2, 192) <= input(42);
output(2, 193) <= input(41);
output(2, 194) <= input(39);
output(2, 195) <= input(40);
output(2, 196) <= input(34);
output(2, 197) <= input(33);
output(2, 198) <= input(17);
output(2, 199) <= input(18);
output(2, 200) <= input(19);
output(2, 201) <= input(20);
output(2, 202) <= input(21);
output(2, 203) <= input(22);
output(2, 204) <= input(23);
output(2, 205) <= input(24);
output(2, 206) <= input(25);
output(2, 207) <= input(26);
output(2, 208) <= input(43);
output(2, 209) <= input(44);
output(2, 210) <= input(45);
output(2, 211) <= input(38);
output(2, 212) <= input(35);
output(2, 213) <= input(36);
output(2, 214) <= input(37);
output(2, 215) <= input(16);
output(2, 216) <= input(0);
output(2, 217) <= input(1);
output(2, 218) <= input(2);
output(2, 219) <= input(3);
output(2, 220) <= input(4);
output(2, 221) <= input(5);
output(2, 222) <= input(6);
output(2, 223) <= input(7);
output(2, 224) <= input(50);
output(2, 225) <= input(42);
output(2, 226) <= input(41);
output(2, 227) <= input(39);
output(2, 228) <= input(40);
output(2, 229) <= input(34);
output(2, 230) <= input(33);
output(2, 231) <= input(17);
output(2, 232) <= input(18);
output(2, 233) <= input(19);
output(2, 234) <= input(20);
output(2, 235) <= input(21);
output(2, 236) <= input(22);
output(2, 237) <= input(23);
output(2, 238) <= input(24);
output(2, 239) <= input(25);
output(2, 240) <= input(46);
output(2, 241) <= input(43);
output(2, 242) <= input(44);
output(2, 243) <= input(45);
output(2, 244) <= input(38);
output(2, 245) <= input(35);
output(2, 246) <= input(36);
output(2, 247) <= input(37);
output(2, 248) <= input(16);
output(2, 249) <= input(0);
output(2, 250) <= input(1);
output(2, 251) <= input(2);
output(2, 252) <= input(3);
output(2, 253) <= input(4);
output(2, 254) <= input(5);
output(2, 255) <= input(6);
when "1010" =>
output(0, 0) <= input(0);
output(0, 1) <= input(1);
output(0, 2) <= input(2);
output(0, 3) <= input(3);
output(0, 4) <= input(4);
output(0, 5) <= input(5);
output(0, 6) <= input(6);
output(0, 7) <= input(7);
output(0, 8) <= input(8);
output(0, 9) <= input(9);
output(0, 10) <= input(10);
output(0, 11) <= input(11);
output(0, 12) <= input(12);
output(0, 13) <= input(13);
output(0, 14) <= input(14);
output(0, 15) <= input(15);
output(0, 16) <= input(16);
output(0, 17) <= input(17);
output(0, 18) <= input(18);
output(0, 19) <= input(19);
output(0, 20) <= input(20);
output(0, 21) <= input(21);
output(0, 22) <= input(22);
output(0, 23) <= input(23);
output(0, 24) <= input(24);
output(0, 25) <= input(25);
output(0, 26) <= input(26);
output(0, 27) <= input(27);
output(0, 28) <= input(28);
output(0, 29) <= input(29);
output(0, 30) <= input(30);
output(0, 31) <= input(31);
output(0, 32) <= input(32);
output(0, 33) <= input(0);
output(0, 34) <= input(1);
output(0, 35) <= input(2);
output(0, 36) <= input(3);
output(0, 37) <= input(4);
output(0, 38) <= input(5);
output(0, 39) <= input(6);
output(0, 40) <= input(7);
output(0, 41) <= input(8);
output(0, 42) <= input(9);
output(0, 43) <= input(10);
output(0, 44) <= input(11);
output(0, 45) <= input(12);
output(0, 46) <= input(13);
output(0, 47) <= input(14);
output(0, 48) <= input(33);
output(0, 49) <= input(16);
output(0, 50) <= input(17);
output(0, 51) <= input(18);
output(0, 52) <= input(19);
output(0, 53) <= input(20);
output(0, 54) <= input(21);
output(0, 55) <= input(22);
output(0, 56) <= input(23);
output(0, 57) <= input(24);
output(0, 58) <= input(25);
output(0, 59) <= input(26);
output(0, 60) <= input(27);
output(0, 61) <= input(28);
output(0, 62) <= input(29);
output(0, 63) <= input(30);
output(0, 64) <= input(34);
output(0, 65) <= input(32);
output(0, 66) <= input(0);
output(0, 67) <= input(1);
output(0, 68) <= input(2);
output(0, 69) <= input(3);
output(0, 70) <= input(4);
output(0, 71) <= input(5);
output(0, 72) <= input(6);
output(0, 73) <= input(7);
output(0, 74) <= input(8);
output(0, 75) <= input(9);
output(0, 76) <= input(10);
output(0, 77) <= input(11);
output(0, 78) <= input(12);
output(0, 79) <= input(13);
output(0, 80) <= input(35);
output(0, 81) <= input(33);
output(0, 82) <= input(16);
output(0, 83) <= input(17);
output(0, 84) <= input(18);
output(0, 85) <= input(19);
output(0, 86) <= input(20);
output(0, 87) <= input(21);
output(0, 88) <= input(22);
output(0, 89) <= input(23);
output(0, 90) <= input(24);
output(0, 91) <= input(25);
output(0, 92) <= input(26);
output(0, 93) <= input(27);
output(0, 94) <= input(28);
output(0, 95) <= input(29);
output(0, 96) <= input(36);
output(0, 97) <= input(34);
output(0, 98) <= input(32);
output(0, 99) <= input(0);
output(0, 100) <= input(1);
output(0, 101) <= input(2);
output(0, 102) <= input(3);
output(0, 103) <= input(4);
output(0, 104) <= input(5);
output(0, 105) <= input(6);
output(0, 106) <= input(7);
output(0, 107) <= input(8);
output(0, 108) <= input(9);
output(0, 109) <= input(10);
output(0, 110) <= input(11);
output(0, 111) <= input(12);
output(0, 112) <= input(37);
output(0, 113) <= input(35);
output(0, 114) <= input(33);
output(0, 115) <= input(16);
output(0, 116) <= input(17);
output(0, 117) <= input(18);
output(0, 118) <= input(19);
output(0, 119) <= input(20);
output(0, 120) <= input(21);
output(0, 121) <= input(22);
output(0, 122) <= input(23);
output(0, 123) <= input(24);
output(0, 124) <= input(25);
output(0, 125) <= input(26);
output(0, 126) <= input(27);
output(0, 127) <= input(28);
output(0, 128) <= input(38);
output(0, 129) <= input(37);
output(0, 130) <= input(35);
output(0, 131) <= input(33);
output(0, 132) <= input(16);
output(0, 133) <= input(17);
output(0, 134) <= input(18);
output(0, 135) <= input(19);
output(0, 136) <= input(20);
output(0, 137) <= input(21);
output(0, 138) <= input(22);
output(0, 139) <= input(23);
output(0, 140) <= input(24);
output(0, 141) <= input(25);
output(0, 142) <= input(26);
output(0, 143) <= input(27);
output(0, 144) <= input(39);
output(0, 145) <= input(40);
output(0, 146) <= input(36);
output(0, 147) <= input(34);
output(0, 148) <= input(32);
output(0, 149) <= input(0);
output(0, 150) <= input(1);
output(0, 151) <= input(2);
output(0, 152) <= input(3);
output(0, 153) <= input(4);
output(0, 154) <= input(5);
output(0, 155) <= input(6);
output(0, 156) <= input(7);
output(0, 157) <= input(8);
output(0, 158) <= input(9);
output(0, 159) <= input(10);
output(0, 160) <= input(41);
output(0, 161) <= input(38);
output(0, 162) <= input(37);
output(0, 163) <= input(35);
output(0, 164) <= input(33);
output(0, 165) <= input(16);
output(0, 166) <= input(17);
output(0, 167) <= input(18);
output(0, 168) <= input(19);
output(0, 169) <= input(20);
output(0, 170) <= input(21);
output(0, 171) <= input(22);
output(0, 172) <= input(23);
output(0, 173) <= input(24);
output(0, 174) <= input(25);
output(0, 175) <= input(26);
output(0, 176) <= input(42);
output(0, 177) <= input(39);
output(0, 178) <= input(40);
output(0, 179) <= input(36);
output(0, 180) <= input(34);
output(0, 181) <= input(32);
output(0, 182) <= input(0);
output(0, 183) <= input(1);
output(0, 184) <= input(2);
output(0, 185) <= input(3);
output(0, 186) <= input(4);
output(0, 187) <= input(5);
output(0, 188) <= input(6);
output(0, 189) <= input(7);
output(0, 190) <= input(8);
output(0, 191) <= input(9);
output(0, 192) <= input(43);
output(0, 193) <= input(41);
output(0, 194) <= input(38);
output(0, 195) <= input(37);
output(0, 196) <= input(35);
output(0, 197) <= input(33);
output(0, 198) <= input(16);
output(0, 199) <= input(17);
output(0, 200) <= input(18);
output(0, 201) <= input(19);
output(0, 202) <= input(20);
output(0, 203) <= input(21);
output(0, 204) <= input(22);
output(0, 205) <= input(23);
output(0, 206) <= input(24);
output(0, 207) <= input(25);
output(0, 208) <= input(44);
output(0, 209) <= input(42);
output(0, 210) <= input(39);
output(0, 211) <= input(40);
output(0, 212) <= input(36);
output(0, 213) <= input(34);
output(0, 214) <= input(32);
output(0, 215) <= input(0);
output(0, 216) <= input(1);
output(0, 217) <= input(2);
output(0, 218) <= input(3);
output(0, 219) <= input(4);
output(0, 220) <= input(5);
output(0, 221) <= input(6);
output(0, 222) <= input(7);
output(0, 223) <= input(8);
output(0, 224) <= input(45);
output(0, 225) <= input(43);
output(0, 226) <= input(41);
output(0, 227) <= input(38);
output(0, 228) <= input(37);
output(0, 229) <= input(35);
output(0, 230) <= input(33);
output(0, 231) <= input(16);
output(0, 232) <= input(17);
output(0, 233) <= input(18);
output(0, 234) <= input(19);
output(0, 235) <= input(20);
output(0, 236) <= input(21);
output(0, 237) <= input(22);
output(0, 238) <= input(23);
output(0, 239) <= input(24);
output(0, 240) <= input(46);
output(0, 241) <= input(44);
output(0, 242) <= input(42);
output(0, 243) <= input(39);
output(0, 244) <= input(40);
output(0, 245) <= input(36);
output(0, 246) <= input(34);
output(0, 247) <= input(32);
output(0, 248) <= input(0);
output(0, 249) <= input(1);
output(0, 250) <= input(2);
output(0, 251) <= input(3);
output(0, 252) <= input(4);
output(0, 253) <= input(5);
output(0, 254) <= input(6);
output(0, 255) <= input(7);
output(1, 0) <= input(17);
output(1, 1) <= input(18);
output(1, 2) <= input(19);
output(1, 3) <= input(20);
output(1, 4) <= input(21);
output(1, 5) <= input(22);
output(1, 6) <= input(23);
output(1, 7) <= input(24);
output(1, 8) <= input(25);
output(1, 9) <= input(26);
output(1, 10) <= input(27);
output(1, 11) <= input(28);
output(1, 12) <= input(29);
output(1, 13) <= input(30);
output(1, 14) <= input(31);
output(1, 15) <= input(47);
output(1, 16) <= input(0);
output(1, 17) <= input(1);
output(1, 18) <= input(2);
output(1, 19) <= input(3);
output(1, 20) <= input(4);
output(1, 21) <= input(5);
output(1, 22) <= input(6);
output(1, 23) <= input(7);
output(1, 24) <= input(8);
output(1, 25) <= input(9);
output(1, 26) <= input(10);
output(1, 27) <= input(11);
output(1, 28) <= input(12);
output(1, 29) <= input(13);
output(1, 30) <= input(14);
output(1, 31) <= input(15);
output(1, 32) <= input(16);
output(1, 33) <= input(17);
output(1, 34) <= input(18);
output(1, 35) <= input(19);
output(1, 36) <= input(20);
output(1, 37) <= input(21);
output(1, 38) <= input(22);
output(1, 39) <= input(23);
output(1, 40) <= input(24);
output(1, 41) <= input(25);
output(1, 42) <= input(26);
output(1, 43) <= input(27);
output(1, 44) <= input(28);
output(1, 45) <= input(29);
output(1, 46) <= input(30);
output(1, 47) <= input(31);
output(1, 48) <= input(32);
output(1, 49) <= input(0);
output(1, 50) <= input(1);
output(1, 51) <= input(2);
output(1, 52) <= input(3);
output(1, 53) <= input(4);
output(1, 54) <= input(5);
output(1, 55) <= input(6);
output(1, 56) <= input(7);
output(1, 57) <= input(8);
output(1, 58) <= input(9);
output(1, 59) <= input(10);
output(1, 60) <= input(11);
output(1, 61) <= input(12);
output(1, 62) <= input(13);
output(1, 63) <= input(14);
output(1, 64) <= input(33);
output(1, 65) <= input(16);
output(1, 66) <= input(17);
output(1, 67) <= input(18);
output(1, 68) <= input(19);
output(1, 69) <= input(20);
output(1, 70) <= input(21);
output(1, 71) <= input(22);
output(1, 72) <= input(23);
output(1, 73) <= input(24);
output(1, 74) <= input(25);
output(1, 75) <= input(26);
output(1, 76) <= input(27);
output(1, 77) <= input(28);
output(1, 78) <= input(29);
output(1, 79) <= input(30);
output(1, 80) <= input(34);
output(1, 81) <= input(32);
output(1, 82) <= input(0);
output(1, 83) <= input(1);
output(1, 84) <= input(2);
output(1, 85) <= input(3);
output(1, 86) <= input(4);
output(1, 87) <= input(5);
output(1, 88) <= input(6);
output(1, 89) <= input(7);
output(1, 90) <= input(8);
output(1, 91) <= input(9);
output(1, 92) <= input(10);
output(1, 93) <= input(11);
output(1, 94) <= input(12);
output(1, 95) <= input(13);
output(1, 96) <= input(35);
output(1, 97) <= input(33);
output(1, 98) <= input(16);
output(1, 99) <= input(17);
output(1, 100) <= input(18);
output(1, 101) <= input(19);
output(1, 102) <= input(20);
output(1, 103) <= input(21);
output(1, 104) <= input(22);
output(1, 105) <= input(23);
output(1, 106) <= input(24);
output(1, 107) <= input(25);
output(1, 108) <= input(26);
output(1, 109) <= input(27);
output(1, 110) <= input(28);
output(1, 111) <= input(29);
output(1, 112) <= input(36);
output(1, 113) <= input(34);
output(1, 114) <= input(32);
output(1, 115) <= input(0);
output(1, 116) <= input(1);
output(1, 117) <= input(2);
output(1, 118) <= input(3);
output(1, 119) <= input(4);
output(1, 120) <= input(5);
output(1, 121) <= input(6);
output(1, 122) <= input(7);
output(1, 123) <= input(8);
output(1, 124) <= input(9);
output(1, 125) <= input(10);
output(1, 126) <= input(11);
output(1, 127) <= input(12);
output(1, 128) <= input(37);
output(1, 129) <= input(35);
output(1, 130) <= input(33);
output(1, 131) <= input(16);
output(1, 132) <= input(17);
output(1, 133) <= input(18);
output(1, 134) <= input(19);
output(1, 135) <= input(20);
output(1, 136) <= input(21);
output(1, 137) <= input(22);
output(1, 138) <= input(23);
output(1, 139) <= input(24);
output(1, 140) <= input(25);
output(1, 141) <= input(26);
output(1, 142) <= input(27);
output(1, 143) <= input(28);
output(1, 144) <= input(40);
output(1, 145) <= input(36);
output(1, 146) <= input(34);
output(1, 147) <= input(32);
output(1, 148) <= input(0);
output(1, 149) <= input(1);
output(1, 150) <= input(2);
output(1, 151) <= input(3);
output(1, 152) <= input(4);
output(1, 153) <= input(5);
output(1, 154) <= input(6);
output(1, 155) <= input(7);
output(1, 156) <= input(8);
output(1, 157) <= input(9);
output(1, 158) <= input(10);
output(1, 159) <= input(11);
output(1, 160) <= input(38);
output(1, 161) <= input(37);
output(1, 162) <= input(35);
output(1, 163) <= input(33);
output(1, 164) <= input(16);
output(1, 165) <= input(17);
output(1, 166) <= input(18);
output(1, 167) <= input(19);
output(1, 168) <= input(20);
output(1, 169) <= input(21);
output(1, 170) <= input(22);
output(1, 171) <= input(23);
output(1, 172) <= input(24);
output(1, 173) <= input(25);
output(1, 174) <= input(26);
output(1, 175) <= input(27);
output(1, 176) <= input(39);
output(1, 177) <= input(40);
output(1, 178) <= input(36);
output(1, 179) <= input(34);
output(1, 180) <= input(32);
output(1, 181) <= input(0);
output(1, 182) <= input(1);
output(1, 183) <= input(2);
output(1, 184) <= input(3);
output(1, 185) <= input(4);
output(1, 186) <= input(5);
output(1, 187) <= input(6);
output(1, 188) <= input(7);
output(1, 189) <= input(8);
output(1, 190) <= input(9);
output(1, 191) <= input(10);
output(1, 192) <= input(41);
output(1, 193) <= input(38);
output(1, 194) <= input(37);
output(1, 195) <= input(35);
output(1, 196) <= input(33);
output(1, 197) <= input(16);
output(1, 198) <= input(17);
output(1, 199) <= input(18);
output(1, 200) <= input(19);
output(1, 201) <= input(20);
output(1, 202) <= input(21);
output(1, 203) <= input(22);
output(1, 204) <= input(23);
output(1, 205) <= input(24);
output(1, 206) <= input(25);
output(1, 207) <= input(26);
output(1, 208) <= input(42);
output(1, 209) <= input(39);
output(1, 210) <= input(40);
output(1, 211) <= input(36);
output(1, 212) <= input(34);
output(1, 213) <= input(32);
output(1, 214) <= input(0);
output(1, 215) <= input(1);
output(1, 216) <= input(2);
output(1, 217) <= input(3);
output(1, 218) <= input(4);
output(1, 219) <= input(5);
output(1, 220) <= input(6);
output(1, 221) <= input(7);
output(1, 222) <= input(8);
output(1, 223) <= input(9);
output(1, 224) <= input(43);
output(1, 225) <= input(41);
output(1, 226) <= input(38);
output(1, 227) <= input(37);
output(1, 228) <= input(35);
output(1, 229) <= input(33);
output(1, 230) <= input(16);
output(1, 231) <= input(17);
output(1, 232) <= input(18);
output(1, 233) <= input(19);
output(1, 234) <= input(20);
output(1, 235) <= input(21);
output(1, 236) <= input(22);
output(1, 237) <= input(23);
output(1, 238) <= input(24);
output(1, 239) <= input(25);
output(1, 240) <= input(44);
output(1, 241) <= input(42);
output(1, 242) <= input(39);
output(1, 243) <= input(40);
output(1, 244) <= input(36);
output(1, 245) <= input(34);
output(1, 246) <= input(32);
output(1, 247) <= input(0);
output(1, 248) <= input(1);
output(1, 249) <= input(2);
output(1, 250) <= input(3);
output(1, 251) <= input(4);
output(1, 252) <= input(5);
output(1, 253) <= input(6);
output(1, 254) <= input(7);
output(1, 255) <= input(8);
when "1011" =>
output(0, 0) <= input(0);
output(0, 1) <= input(1);
output(0, 2) <= input(2);
output(0, 3) <= input(3);
output(0, 4) <= input(4);
output(0, 5) <= input(5);
output(0, 6) <= input(6);
output(0, 7) <= input(7);
output(0, 8) <= input(8);
output(0, 9) <= input(9);
output(0, 10) <= input(10);
output(0, 11) <= input(11);
output(0, 12) <= input(12);
output(0, 13) <= input(13);
output(0, 14) <= input(14);
output(0, 15) <= input(15);
output(0, 16) <= input(16);
output(0, 17) <= input(17);
output(0, 18) <= input(18);
output(0, 19) <= input(19);
output(0, 20) <= input(20);
output(0, 21) <= input(21);
output(0, 22) <= input(22);
output(0, 23) <= input(23);
output(0, 24) <= input(24);
output(0, 25) <= input(25);
output(0, 26) <= input(26);
output(0, 27) <= input(27);
output(0, 28) <= input(28);
output(0, 29) <= input(29);
output(0, 30) <= input(30);
output(0, 31) <= input(31);
output(0, 32) <= input(32);
output(0, 33) <= input(0);
output(0, 34) <= input(1);
output(0, 35) <= input(2);
output(0, 36) <= input(3);
output(0, 37) <= input(4);
output(0, 38) <= input(5);
output(0, 39) <= input(6);
output(0, 40) <= input(7);
output(0, 41) <= input(8);
output(0, 42) <= input(9);
output(0, 43) <= input(10);
output(0, 44) <= input(11);
output(0, 45) <= input(12);
output(0, 46) <= input(13);
output(0, 47) <= input(14);
output(0, 48) <= input(33);
output(0, 49) <= input(16);
output(0, 50) <= input(17);
output(0, 51) <= input(18);
output(0, 52) <= input(19);
output(0, 53) <= input(20);
output(0, 54) <= input(21);
output(0, 55) <= input(22);
output(0, 56) <= input(23);
output(0, 57) <= input(24);
output(0, 58) <= input(25);
output(0, 59) <= input(26);
output(0, 60) <= input(27);
output(0, 61) <= input(28);
output(0, 62) <= input(29);
output(0, 63) <= input(30);
output(0, 64) <= input(34);
output(0, 65) <= input(32);
output(0, 66) <= input(0);
output(0, 67) <= input(1);
output(0, 68) <= input(2);
output(0, 69) <= input(3);
output(0, 70) <= input(4);
output(0, 71) <= input(5);
output(0, 72) <= input(6);
output(0, 73) <= input(7);
output(0, 74) <= input(8);
output(0, 75) <= input(9);
output(0, 76) <= input(10);
output(0, 77) <= input(11);
output(0, 78) <= input(12);
output(0, 79) <= input(13);
output(0, 80) <= input(35);
output(0, 81) <= input(33);
output(0, 82) <= input(16);
output(0, 83) <= input(17);
output(0, 84) <= input(18);
output(0, 85) <= input(19);
output(0, 86) <= input(20);
output(0, 87) <= input(21);
output(0, 88) <= input(22);
output(0, 89) <= input(23);
output(0, 90) <= input(24);
output(0, 91) <= input(25);
output(0, 92) <= input(26);
output(0, 93) <= input(27);
output(0, 94) <= input(28);
output(0, 95) <= input(29);
output(0, 96) <= input(36);
output(0, 97) <= input(34);
output(0, 98) <= input(32);
output(0, 99) <= input(0);
output(0, 100) <= input(1);
output(0, 101) <= input(2);
output(0, 102) <= input(3);
output(0, 103) <= input(4);
output(0, 104) <= input(5);
output(0, 105) <= input(6);
output(0, 106) <= input(7);
output(0, 107) <= input(8);
output(0, 108) <= input(9);
output(0, 109) <= input(10);
output(0, 110) <= input(11);
output(0, 111) <= input(12);
output(0, 112) <= input(36);
output(0, 113) <= input(34);
output(0, 114) <= input(32);
output(0, 115) <= input(0);
output(0, 116) <= input(1);
output(0, 117) <= input(2);
output(0, 118) <= input(3);
output(0, 119) <= input(4);
output(0, 120) <= input(5);
output(0, 121) <= input(6);
output(0, 122) <= input(7);
output(0, 123) <= input(8);
output(0, 124) <= input(9);
output(0, 125) <= input(10);
output(0, 126) <= input(11);
output(0, 127) <= input(12);
output(0, 128) <= input(37);
output(0, 129) <= input(35);
output(0, 130) <= input(33);
output(0, 131) <= input(16);
output(0, 132) <= input(17);
output(0, 133) <= input(18);
output(0, 134) <= input(19);
output(0, 135) <= input(20);
output(0, 136) <= input(21);
output(0, 137) <= input(22);
output(0, 138) <= input(23);
output(0, 139) <= input(24);
output(0, 140) <= input(25);
output(0, 141) <= input(26);
output(0, 142) <= input(27);
output(0, 143) <= input(28);
output(0, 144) <= input(38);
output(0, 145) <= input(36);
output(0, 146) <= input(34);
output(0, 147) <= input(32);
output(0, 148) <= input(0);
output(0, 149) <= input(1);
output(0, 150) <= input(2);
output(0, 151) <= input(3);
output(0, 152) <= input(4);
output(0, 153) <= input(5);
output(0, 154) <= input(6);
output(0, 155) <= input(7);
output(0, 156) <= input(8);
output(0, 157) <= input(9);
output(0, 158) <= input(10);
output(0, 159) <= input(11);
output(0, 160) <= input(39);
output(0, 161) <= input(37);
output(0, 162) <= input(35);
output(0, 163) <= input(33);
output(0, 164) <= input(16);
output(0, 165) <= input(17);
output(0, 166) <= input(18);
output(0, 167) <= input(19);
output(0, 168) <= input(20);
output(0, 169) <= input(21);
output(0, 170) <= input(22);
output(0, 171) <= input(23);
output(0, 172) <= input(24);
output(0, 173) <= input(25);
output(0, 174) <= input(26);
output(0, 175) <= input(27);
output(0, 176) <= input(40);
output(0, 177) <= input(38);
output(0, 178) <= input(36);
output(0, 179) <= input(34);
output(0, 180) <= input(32);
output(0, 181) <= input(0);
output(0, 182) <= input(1);
output(0, 183) <= input(2);
output(0, 184) <= input(3);
output(0, 185) <= input(4);
output(0, 186) <= input(5);
output(0, 187) <= input(6);
output(0, 188) <= input(7);
output(0, 189) <= input(8);
output(0, 190) <= input(9);
output(0, 191) <= input(10);
output(0, 192) <= input(41);
output(0, 193) <= input(39);
output(0, 194) <= input(37);
output(0, 195) <= input(35);
output(0, 196) <= input(33);
output(0, 197) <= input(16);
output(0, 198) <= input(17);
output(0, 199) <= input(18);
output(0, 200) <= input(19);
output(0, 201) <= input(20);
output(0, 202) <= input(21);
output(0, 203) <= input(22);
output(0, 204) <= input(23);
output(0, 205) <= input(24);
output(0, 206) <= input(25);
output(0, 207) <= input(26);
output(0, 208) <= input(42);
output(0, 209) <= input(40);
output(0, 210) <= input(38);
output(0, 211) <= input(36);
output(0, 212) <= input(34);
output(0, 213) <= input(32);
output(0, 214) <= input(0);
output(0, 215) <= input(1);
output(0, 216) <= input(2);
output(0, 217) <= input(3);
output(0, 218) <= input(4);
output(0, 219) <= input(5);
output(0, 220) <= input(6);
output(0, 221) <= input(7);
output(0, 222) <= input(8);
output(0, 223) <= input(9);
output(0, 224) <= input(43);
output(0, 225) <= input(41);
output(0, 226) <= input(39);
output(0, 227) <= input(37);
output(0, 228) <= input(35);
output(0, 229) <= input(33);
output(0, 230) <= input(16);
output(0, 231) <= input(17);
output(0, 232) <= input(18);
output(0, 233) <= input(19);
output(0, 234) <= input(20);
output(0, 235) <= input(21);
output(0, 236) <= input(22);
output(0, 237) <= input(23);
output(0, 238) <= input(24);
output(0, 239) <= input(25);
output(0, 240) <= input(43);
output(0, 241) <= input(41);
output(0, 242) <= input(39);
output(0, 243) <= input(37);
output(0, 244) <= input(35);
output(0, 245) <= input(33);
output(0, 246) <= input(16);
output(0, 247) <= input(17);
output(0, 248) <= input(18);
output(0, 249) <= input(19);
output(0, 250) <= input(20);
output(0, 251) <= input(21);
output(0, 252) <= input(22);
output(0, 253) <= input(23);
output(0, 254) <= input(24);
output(0, 255) <= input(25);
output(1, 0) <= input(0);
output(1, 1) <= input(1);
output(1, 2) <= input(2);
output(1, 3) <= input(3);
output(1, 4) <= input(4);
output(1, 5) <= input(5);
output(1, 6) <= input(6);
output(1, 7) <= input(7);
output(1, 8) <= input(8);
output(1, 9) <= input(9);
output(1, 10) <= input(10);
output(1, 11) <= input(11);
output(1, 12) <= input(12);
output(1, 13) <= input(13);
output(1, 14) <= input(14);
output(1, 15) <= input(15);
output(1, 16) <= input(16);
output(1, 17) <= input(17);
output(1, 18) <= input(18);
output(1, 19) <= input(19);
output(1, 20) <= input(20);
output(1, 21) <= input(21);
output(1, 22) <= input(22);
output(1, 23) <= input(23);
output(1, 24) <= input(24);
output(1, 25) <= input(25);
output(1, 26) <= input(26);
output(1, 27) <= input(27);
output(1, 28) <= input(28);
output(1, 29) <= input(29);
output(1, 30) <= input(30);
output(1, 31) <= input(31);
output(1, 32) <= input(32);
output(1, 33) <= input(0);
output(1, 34) <= input(1);
output(1, 35) <= input(2);
output(1, 36) <= input(3);
output(1, 37) <= input(4);
output(1, 38) <= input(5);
output(1, 39) <= input(6);
output(1, 40) <= input(7);
output(1, 41) <= input(8);
output(1, 42) <= input(9);
output(1, 43) <= input(10);
output(1, 44) <= input(11);
output(1, 45) <= input(12);
output(1, 46) <= input(13);
output(1, 47) <= input(14);
output(1, 48) <= input(32);
output(1, 49) <= input(0);
output(1, 50) <= input(1);
output(1, 51) <= input(2);
output(1, 52) <= input(3);
output(1, 53) <= input(4);
output(1, 54) <= input(5);
output(1, 55) <= input(6);
output(1, 56) <= input(7);
output(1, 57) <= input(8);
output(1, 58) <= input(9);
output(1, 59) <= input(10);
output(1, 60) <= input(11);
output(1, 61) <= input(12);
output(1, 62) <= input(13);
output(1, 63) <= input(14);
output(1, 64) <= input(33);
output(1, 65) <= input(16);
output(1, 66) <= input(17);
output(1, 67) <= input(18);
output(1, 68) <= input(19);
output(1, 69) <= input(20);
output(1, 70) <= input(21);
output(1, 71) <= input(22);
output(1, 72) <= input(23);
output(1, 73) <= input(24);
output(1, 74) <= input(25);
output(1, 75) <= input(26);
output(1, 76) <= input(27);
output(1, 77) <= input(28);
output(1, 78) <= input(29);
output(1, 79) <= input(30);
output(1, 80) <= input(34);
output(1, 81) <= input(32);
output(1, 82) <= input(0);
output(1, 83) <= input(1);
output(1, 84) <= input(2);
output(1, 85) <= input(3);
output(1, 86) <= input(4);
output(1, 87) <= input(5);
output(1, 88) <= input(6);
output(1, 89) <= input(7);
output(1, 90) <= input(8);
output(1, 91) <= input(9);
output(1, 92) <= input(10);
output(1, 93) <= input(11);
output(1, 94) <= input(12);
output(1, 95) <= input(13);
output(1, 96) <= input(35);
output(1, 97) <= input(33);
output(1, 98) <= input(16);
output(1, 99) <= input(17);
output(1, 100) <= input(18);
output(1, 101) <= input(19);
output(1, 102) <= input(20);
output(1, 103) <= input(21);
output(1, 104) <= input(22);
output(1, 105) <= input(23);
output(1, 106) <= input(24);
output(1, 107) <= input(25);
output(1, 108) <= input(26);
output(1, 109) <= input(27);
output(1, 110) <= input(28);
output(1, 111) <= input(29);
output(1, 112) <= input(35);
output(1, 113) <= input(33);
output(1, 114) <= input(16);
output(1, 115) <= input(17);
output(1, 116) <= input(18);
output(1, 117) <= input(19);
output(1, 118) <= input(20);
output(1, 119) <= input(21);
output(1, 120) <= input(22);
output(1, 121) <= input(23);
output(1, 122) <= input(24);
output(1, 123) <= input(25);
output(1, 124) <= input(26);
output(1, 125) <= input(27);
output(1, 126) <= input(28);
output(1, 127) <= input(29);
output(1, 128) <= input(36);
output(1, 129) <= input(34);
output(1, 130) <= input(32);
output(1, 131) <= input(0);
output(1, 132) <= input(1);
output(1, 133) <= input(2);
output(1, 134) <= input(3);
output(1, 135) <= input(4);
output(1, 136) <= input(5);
output(1, 137) <= input(6);
output(1, 138) <= input(7);
output(1, 139) <= input(8);
output(1, 140) <= input(9);
output(1, 141) <= input(10);
output(1, 142) <= input(11);
output(1, 143) <= input(12);
output(1, 144) <= input(37);
output(1, 145) <= input(35);
output(1, 146) <= input(33);
output(1, 147) <= input(16);
output(1, 148) <= input(17);
output(1, 149) <= input(18);
output(1, 150) <= input(19);
output(1, 151) <= input(20);
output(1, 152) <= input(21);
output(1, 153) <= input(22);
output(1, 154) <= input(23);
output(1, 155) <= input(24);
output(1, 156) <= input(25);
output(1, 157) <= input(26);
output(1, 158) <= input(27);
output(1, 159) <= input(28);
output(1, 160) <= input(38);
output(1, 161) <= input(36);
output(1, 162) <= input(34);
output(1, 163) <= input(32);
output(1, 164) <= input(0);
output(1, 165) <= input(1);
output(1, 166) <= input(2);
output(1, 167) <= input(3);
output(1, 168) <= input(4);
output(1, 169) <= input(5);
output(1, 170) <= input(6);
output(1, 171) <= input(7);
output(1, 172) <= input(8);
output(1, 173) <= input(9);
output(1, 174) <= input(10);
output(1, 175) <= input(11);
output(1, 176) <= input(38);
output(1, 177) <= input(36);
output(1, 178) <= input(34);
output(1, 179) <= input(32);
output(1, 180) <= input(0);
output(1, 181) <= input(1);
output(1, 182) <= input(2);
output(1, 183) <= input(3);
output(1, 184) <= input(4);
output(1, 185) <= input(5);
output(1, 186) <= input(6);
output(1, 187) <= input(7);
output(1, 188) <= input(8);
output(1, 189) <= input(9);
output(1, 190) <= input(10);
output(1, 191) <= input(11);
output(1, 192) <= input(39);
output(1, 193) <= input(37);
output(1, 194) <= input(35);
output(1, 195) <= input(33);
output(1, 196) <= input(16);
output(1, 197) <= input(17);
output(1, 198) <= input(18);
output(1, 199) <= input(19);
output(1, 200) <= input(20);
output(1, 201) <= input(21);
output(1, 202) <= input(22);
output(1, 203) <= input(23);
output(1, 204) <= input(24);
output(1, 205) <= input(25);
output(1, 206) <= input(26);
output(1, 207) <= input(27);
output(1, 208) <= input(40);
output(1, 209) <= input(38);
output(1, 210) <= input(36);
output(1, 211) <= input(34);
output(1, 212) <= input(32);
output(1, 213) <= input(0);
output(1, 214) <= input(1);
output(1, 215) <= input(2);
output(1, 216) <= input(3);
output(1, 217) <= input(4);
output(1, 218) <= input(5);
output(1, 219) <= input(6);
output(1, 220) <= input(7);
output(1, 221) <= input(8);
output(1, 222) <= input(9);
output(1, 223) <= input(10);
output(1, 224) <= input(41);
output(1, 225) <= input(39);
output(1, 226) <= input(37);
output(1, 227) <= input(35);
output(1, 228) <= input(33);
output(1, 229) <= input(16);
output(1, 230) <= input(17);
output(1, 231) <= input(18);
output(1, 232) <= input(19);
output(1, 233) <= input(20);
output(1, 234) <= input(21);
output(1, 235) <= input(22);
output(1, 236) <= input(23);
output(1, 237) <= input(24);
output(1, 238) <= input(25);
output(1, 239) <= input(26);
output(1, 240) <= input(41);
output(1, 241) <= input(39);
output(1, 242) <= input(37);
output(1, 243) <= input(35);
output(1, 244) <= input(33);
output(1, 245) <= input(16);
output(1, 246) <= input(17);
output(1, 247) <= input(18);
output(1, 248) <= input(19);
output(1, 249) <= input(20);
output(1, 250) <= input(21);
output(1, 251) <= input(22);
output(1, 252) <= input(23);
output(1, 253) <= input(24);
output(1, 254) <= input(25);
output(1, 255) <= input(26);
output(2, 0) <= input(0);
output(2, 1) <= input(1);
output(2, 2) <= input(2);
output(2, 3) <= input(3);
output(2, 4) <= input(4);
output(2, 5) <= input(5);
output(2, 6) <= input(6);
output(2, 7) <= input(7);
output(2, 8) <= input(8);
output(2, 9) <= input(9);
output(2, 10) <= input(10);
output(2, 11) <= input(11);
output(2, 12) <= input(12);
output(2, 13) <= input(13);
output(2, 14) <= input(14);
output(2, 15) <= input(15);
output(2, 16) <= input(16);
output(2, 17) <= input(17);
output(2, 18) <= input(18);
output(2, 19) <= input(19);
output(2, 20) <= input(20);
output(2, 21) <= input(21);
output(2, 22) <= input(22);
output(2, 23) <= input(23);
output(2, 24) <= input(24);
output(2, 25) <= input(25);
output(2, 26) <= input(26);
output(2, 27) <= input(27);
output(2, 28) <= input(28);
output(2, 29) <= input(29);
output(2, 30) <= input(30);
output(2, 31) <= input(31);
output(2, 32) <= input(16);
output(2, 33) <= input(17);
output(2, 34) <= input(18);
output(2, 35) <= input(19);
output(2, 36) <= input(20);
output(2, 37) <= input(21);
output(2, 38) <= input(22);
output(2, 39) <= input(23);
output(2, 40) <= input(24);
output(2, 41) <= input(25);
output(2, 42) <= input(26);
output(2, 43) <= input(27);
output(2, 44) <= input(28);
output(2, 45) <= input(29);
output(2, 46) <= input(30);
output(2, 47) <= input(31);
output(2, 48) <= input(32);
output(2, 49) <= input(0);
output(2, 50) <= input(1);
output(2, 51) <= input(2);
output(2, 52) <= input(3);
output(2, 53) <= input(4);
output(2, 54) <= input(5);
output(2, 55) <= input(6);
output(2, 56) <= input(7);
output(2, 57) <= input(8);
output(2, 58) <= input(9);
output(2, 59) <= input(10);
output(2, 60) <= input(11);
output(2, 61) <= input(12);
output(2, 62) <= input(13);
output(2, 63) <= input(14);
output(2, 64) <= input(33);
output(2, 65) <= input(16);
output(2, 66) <= input(17);
output(2, 67) <= input(18);
output(2, 68) <= input(19);
output(2, 69) <= input(20);
output(2, 70) <= input(21);
output(2, 71) <= input(22);
output(2, 72) <= input(23);
output(2, 73) <= input(24);
output(2, 74) <= input(25);
output(2, 75) <= input(26);
output(2, 76) <= input(27);
output(2, 77) <= input(28);
output(2, 78) <= input(29);
output(2, 79) <= input(30);
output(2, 80) <= input(33);
output(2, 81) <= input(16);
output(2, 82) <= input(17);
output(2, 83) <= input(18);
output(2, 84) <= input(19);
output(2, 85) <= input(20);
output(2, 86) <= input(21);
output(2, 87) <= input(22);
output(2, 88) <= input(23);
output(2, 89) <= input(24);
output(2, 90) <= input(25);
output(2, 91) <= input(26);
output(2, 92) <= input(27);
output(2, 93) <= input(28);
output(2, 94) <= input(29);
output(2, 95) <= input(30);
output(2, 96) <= input(34);
output(2, 97) <= input(32);
output(2, 98) <= input(0);
output(2, 99) <= input(1);
output(2, 100) <= input(2);
output(2, 101) <= input(3);
output(2, 102) <= input(4);
output(2, 103) <= input(5);
output(2, 104) <= input(6);
output(2, 105) <= input(7);
output(2, 106) <= input(8);
output(2, 107) <= input(9);
output(2, 108) <= input(10);
output(2, 109) <= input(11);
output(2, 110) <= input(12);
output(2, 111) <= input(13);
output(2, 112) <= input(34);
output(2, 113) <= input(32);
output(2, 114) <= input(0);
output(2, 115) <= input(1);
output(2, 116) <= input(2);
output(2, 117) <= input(3);
output(2, 118) <= input(4);
output(2, 119) <= input(5);
output(2, 120) <= input(6);
output(2, 121) <= input(7);
output(2, 122) <= input(8);
output(2, 123) <= input(9);
output(2, 124) <= input(10);
output(2, 125) <= input(11);
output(2, 126) <= input(12);
output(2, 127) <= input(13);
output(2, 128) <= input(35);
output(2, 129) <= input(33);
output(2, 130) <= input(16);
output(2, 131) <= input(17);
output(2, 132) <= input(18);
output(2, 133) <= input(19);
output(2, 134) <= input(20);
output(2, 135) <= input(21);
output(2, 136) <= input(22);
output(2, 137) <= input(23);
output(2, 138) <= input(24);
output(2, 139) <= input(25);
output(2, 140) <= input(26);
output(2, 141) <= input(27);
output(2, 142) <= input(28);
output(2, 143) <= input(29);
output(2, 144) <= input(36);
output(2, 145) <= input(34);
output(2, 146) <= input(32);
output(2, 147) <= input(0);
output(2, 148) <= input(1);
output(2, 149) <= input(2);
output(2, 150) <= input(3);
output(2, 151) <= input(4);
output(2, 152) <= input(5);
output(2, 153) <= input(6);
output(2, 154) <= input(7);
output(2, 155) <= input(8);
output(2, 156) <= input(9);
output(2, 157) <= input(10);
output(2, 158) <= input(11);
output(2, 159) <= input(12);
output(2, 160) <= input(36);
output(2, 161) <= input(34);
output(2, 162) <= input(32);
output(2, 163) <= input(0);
output(2, 164) <= input(1);
output(2, 165) <= input(2);
output(2, 166) <= input(3);
output(2, 167) <= input(4);
output(2, 168) <= input(5);
output(2, 169) <= input(6);
output(2, 170) <= input(7);
output(2, 171) <= input(8);
output(2, 172) <= input(9);
output(2, 173) <= input(10);
output(2, 174) <= input(11);
output(2, 175) <= input(12);
output(2, 176) <= input(37);
output(2, 177) <= input(35);
output(2, 178) <= input(33);
output(2, 179) <= input(16);
output(2, 180) <= input(17);
output(2, 181) <= input(18);
output(2, 182) <= input(19);
output(2, 183) <= input(20);
output(2, 184) <= input(21);
output(2, 185) <= input(22);
output(2, 186) <= input(23);
output(2, 187) <= input(24);
output(2, 188) <= input(25);
output(2, 189) <= input(26);
output(2, 190) <= input(27);
output(2, 191) <= input(28);
output(2, 192) <= input(38);
output(2, 193) <= input(36);
output(2, 194) <= input(34);
output(2, 195) <= input(32);
output(2, 196) <= input(0);
output(2, 197) <= input(1);
output(2, 198) <= input(2);
output(2, 199) <= input(3);
output(2, 200) <= input(4);
output(2, 201) <= input(5);
output(2, 202) <= input(6);
output(2, 203) <= input(7);
output(2, 204) <= input(8);
output(2, 205) <= input(9);
output(2, 206) <= input(10);
output(2, 207) <= input(11);
output(2, 208) <= input(38);
output(2, 209) <= input(36);
output(2, 210) <= input(34);
output(2, 211) <= input(32);
output(2, 212) <= input(0);
output(2, 213) <= input(1);
output(2, 214) <= input(2);
output(2, 215) <= input(3);
output(2, 216) <= input(4);
output(2, 217) <= input(5);
output(2, 218) <= input(6);
output(2, 219) <= input(7);
output(2, 220) <= input(8);
output(2, 221) <= input(9);
output(2, 222) <= input(10);
output(2, 223) <= input(11);
output(2, 224) <= input(39);
output(2, 225) <= input(37);
output(2, 226) <= input(35);
output(2, 227) <= input(33);
output(2, 228) <= input(16);
output(2, 229) <= input(17);
output(2, 230) <= input(18);
output(2, 231) <= input(19);
output(2, 232) <= input(20);
output(2, 233) <= input(21);
output(2, 234) <= input(22);
output(2, 235) <= input(23);
output(2, 236) <= input(24);
output(2, 237) <= input(25);
output(2, 238) <= input(26);
output(2, 239) <= input(27);
output(2, 240) <= input(39);
output(2, 241) <= input(37);
output(2, 242) <= input(35);
output(2, 243) <= input(33);
output(2, 244) <= input(16);
output(2, 245) <= input(17);
output(2, 246) <= input(18);
output(2, 247) <= input(19);
output(2, 248) <= input(20);
output(2, 249) <= input(21);
output(2, 250) <= input(22);
output(2, 251) <= input(23);
output(2, 252) <= input(24);
output(2, 253) <= input(25);
output(2, 254) <= input(26);
output(2, 255) <= input(27);
when "1100" =>
output(0, 0) <= input(0);
output(0, 1) <= input(1);
output(0, 2) <= input(2);
output(0, 3) <= input(3);
output(0, 4) <= input(4);
output(0, 5) <= input(5);
output(0, 6) <= input(6);
output(0, 7) <= input(7);
output(0, 8) <= input(8);
output(0, 9) <= input(9);
output(0, 10) <= input(10);
output(0, 11) <= input(11);
output(0, 12) <= input(12);
output(0, 13) <= input(13);
output(0, 14) <= input(14);
output(0, 15) <= input(15);
output(0, 16) <= input(0);
output(0, 17) <= input(1);
output(0, 18) <= input(2);
output(0, 19) <= input(3);
output(0, 20) <= input(4);
output(0, 21) <= input(5);
output(0, 22) <= input(6);
output(0, 23) <= input(7);
output(0, 24) <= input(8);
output(0, 25) <= input(9);
output(0, 26) <= input(10);
output(0, 27) <= input(11);
output(0, 28) <= input(12);
output(0, 29) <= input(13);
output(0, 30) <= input(14);
output(0, 31) <= input(15);
output(0, 32) <= input(16);
output(0, 33) <= input(17);
output(0, 34) <= input(18);
output(0, 35) <= input(19);
output(0, 36) <= input(20);
output(0, 37) <= input(21);
output(0, 38) <= input(22);
output(0, 39) <= input(23);
output(0, 40) <= input(24);
output(0, 41) <= input(25);
output(0, 42) <= input(26);
output(0, 43) <= input(27);
output(0, 44) <= input(28);
output(0, 45) <= input(29);
output(0, 46) <= input(30);
output(0, 47) <= input(31);
output(0, 48) <= input(16);
output(0, 49) <= input(17);
output(0, 50) <= input(18);
output(0, 51) <= input(19);
output(0, 52) <= input(20);
output(0, 53) <= input(21);
output(0, 54) <= input(22);
output(0, 55) <= input(23);
output(0, 56) <= input(24);
output(0, 57) <= input(25);
output(0, 58) <= input(26);
output(0, 59) <= input(27);
output(0, 60) <= input(28);
output(0, 61) <= input(29);
output(0, 62) <= input(30);
output(0, 63) <= input(31);
output(0, 64) <= input(32);
output(0, 65) <= input(0);
output(0, 66) <= input(1);
output(0, 67) <= input(2);
output(0, 68) <= input(3);
output(0, 69) <= input(4);
output(0, 70) <= input(5);
output(0, 71) <= input(6);
output(0, 72) <= input(7);
output(0, 73) <= input(8);
output(0, 74) <= input(9);
output(0, 75) <= input(10);
output(0, 76) <= input(11);
output(0, 77) <= input(12);
output(0, 78) <= input(13);
output(0, 79) <= input(14);
output(0, 80) <= input(32);
output(0, 81) <= input(0);
output(0, 82) <= input(1);
output(0, 83) <= input(2);
output(0, 84) <= input(3);
output(0, 85) <= input(4);
output(0, 86) <= input(5);
output(0, 87) <= input(6);
output(0, 88) <= input(7);
output(0, 89) <= input(8);
output(0, 90) <= input(9);
output(0, 91) <= input(10);
output(0, 92) <= input(11);
output(0, 93) <= input(12);
output(0, 94) <= input(13);
output(0, 95) <= input(14);
output(0, 96) <= input(33);
output(0, 97) <= input(16);
output(0, 98) <= input(17);
output(0, 99) <= input(18);
output(0, 100) <= input(19);
output(0, 101) <= input(20);
output(0, 102) <= input(21);
output(0, 103) <= input(22);
output(0, 104) <= input(23);
output(0, 105) <= input(24);
output(0, 106) <= input(25);
output(0, 107) <= input(26);
output(0, 108) <= input(27);
output(0, 109) <= input(28);
output(0, 110) <= input(29);
output(0, 111) <= input(30);
output(0, 112) <= input(33);
output(0, 113) <= input(16);
output(0, 114) <= input(17);
output(0, 115) <= input(18);
output(0, 116) <= input(19);
output(0, 117) <= input(20);
output(0, 118) <= input(21);
output(0, 119) <= input(22);
output(0, 120) <= input(23);
output(0, 121) <= input(24);
output(0, 122) <= input(25);
output(0, 123) <= input(26);
output(0, 124) <= input(27);
output(0, 125) <= input(28);
output(0, 126) <= input(29);
output(0, 127) <= input(30);
output(0, 128) <= input(34);
output(0, 129) <= input(32);
output(0, 130) <= input(0);
output(0, 131) <= input(1);
output(0, 132) <= input(2);
output(0, 133) <= input(3);
output(0, 134) <= input(4);
output(0, 135) <= input(5);
output(0, 136) <= input(6);
output(0, 137) <= input(7);
output(0, 138) <= input(8);
output(0, 139) <= input(9);
output(0, 140) <= input(10);
output(0, 141) <= input(11);
output(0, 142) <= input(12);
output(0, 143) <= input(13);
output(0, 144) <= input(34);
output(0, 145) <= input(32);
output(0, 146) <= input(0);
output(0, 147) <= input(1);
output(0, 148) <= input(2);
output(0, 149) <= input(3);
output(0, 150) <= input(4);
output(0, 151) <= input(5);
output(0, 152) <= input(6);
output(0, 153) <= input(7);
output(0, 154) <= input(8);
output(0, 155) <= input(9);
output(0, 156) <= input(10);
output(0, 157) <= input(11);
output(0, 158) <= input(12);
output(0, 159) <= input(13);
output(0, 160) <= input(35);
output(0, 161) <= input(33);
output(0, 162) <= input(16);
output(0, 163) <= input(17);
output(0, 164) <= input(18);
output(0, 165) <= input(19);
output(0, 166) <= input(20);
output(0, 167) <= input(21);
output(0, 168) <= input(22);
output(0, 169) <= input(23);
output(0, 170) <= input(24);
output(0, 171) <= input(25);
output(0, 172) <= input(26);
output(0, 173) <= input(27);
output(0, 174) <= input(28);
output(0, 175) <= input(29);
output(0, 176) <= input(35);
output(0, 177) <= input(33);
output(0, 178) <= input(16);
output(0, 179) <= input(17);
output(0, 180) <= input(18);
output(0, 181) <= input(19);
output(0, 182) <= input(20);
output(0, 183) <= input(21);
output(0, 184) <= input(22);
output(0, 185) <= input(23);
output(0, 186) <= input(24);
output(0, 187) <= input(25);
output(0, 188) <= input(26);
output(0, 189) <= input(27);
output(0, 190) <= input(28);
output(0, 191) <= input(29);
output(0, 192) <= input(36);
output(0, 193) <= input(34);
output(0, 194) <= input(32);
output(0, 195) <= input(0);
output(0, 196) <= input(1);
output(0, 197) <= input(2);
output(0, 198) <= input(3);
output(0, 199) <= input(4);
output(0, 200) <= input(5);
output(0, 201) <= input(6);
output(0, 202) <= input(7);
output(0, 203) <= input(8);
output(0, 204) <= input(9);
output(0, 205) <= input(10);
output(0, 206) <= input(11);
output(0, 207) <= input(12);
output(0, 208) <= input(36);
output(0, 209) <= input(34);
output(0, 210) <= input(32);
output(0, 211) <= input(0);
output(0, 212) <= input(1);
output(0, 213) <= input(2);
output(0, 214) <= input(3);
output(0, 215) <= input(4);
output(0, 216) <= input(5);
output(0, 217) <= input(6);
output(0, 218) <= input(7);
output(0, 219) <= input(8);
output(0, 220) <= input(9);
output(0, 221) <= input(10);
output(0, 222) <= input(11);
output(0, 223) <= input(12);
output(0, 224) <= input(37);
output(0, 225) <= input(35);
output(0, 226) <= input(33);
output(0, 227) <= input(16);
output(0, 228) <= input(17);
output(0, 229) <= input(18);
output(0, 230) <= input(19);
output(0, 231) <= input(20);
output(0, 232) <= input(21);
output(0, 233) <= input(22);
output(0, 234) <= input(23);
output(0, 235) <= input(24);
output(0, 236) <= input(25);
output(0, 237) <= input(26);
output(0, 238) <= input(27);
output(0, 239) <= input(28);
output(0, 240) <= input(37);
output(0, 241) <= input(35);
output(0, 242) <= input(33);
output(0, 243) <= input(16);
output(0, 244) <= input(17);
output(0, 245) <= input(18);
output(0, 246) <= input(19);
output(0, 247) <= input(20);
output(0, 248) <= input(21);
output(0, 249) <= input(22);
output(0, 250) <= input(23);
output(0, 251) <= input(24);
output(0, 252) <= input(25);
output(0, 253) <= input(26);
output(0, 254) <= input(27);
output(0, 255) <= input(28);
output(1, 0) <= input(0);
output(1, 1) <= input(1);
output(1, 2) <= input(2);
output(1, 3) <= input(3);
output(1, 4) <= input(4);
output(1, 5) <= input(5);
output(1, 6) <= input(6);
output(1, 7) <= input(7);
output(1, 8) <= input(8);
output(1, 9) <= input(9);
output(1, 10) <= input(10);
output(1, 11) <= input(11);
output(1, 12) <= input(12);
output(1, 13) <= input(13);
output(1, 14) <= input(14);
output(1, 15) <= input(15);
output(1, 16) <= input(0);
output(1, 17) <= input(1);
output(1, 18) <= input(2);
output(1, 19) <= input(3);
output(1, 20) <= input(4);
output(1, 21) <= input(5);
output(1, 22) <= input(6);
output(1, 23) <= input(7);
output(1, 24) <= input(8);
output(1, 25) <= input(9);
output(1, 26) <= input(10);
output(1, 27) <= input(11);
output(1, 28) <= input(12);
output(1, 29) <= input(13);
output(1, 30) <= input(14);
output(1, 31) <= input(15);
output(1, 32) <= input(16);
output(1, 33) <= input(17);
output(1, 34) <= input(18);
output(1, 35) <= input(19);
output(1, 36) <= input(20);
output(1, 37) <= input(21);
output(1, 38) <= input(22);
output(1, 39) <= input(23);
output(1, 40) <= input(24);
output(1, 41) <= input(25);
output(1, 42) <= input(26);
output(1, 43) <= input(27);
output(1, 44) <= input(28);
output(1, 45) <= input(29);
output(1, 46) <= input(30);
output(1, 47) <= input(31);
output(1, 48) <= input(16);
output(1, 49) <= input(17);
output(1, 50) <= input(18);
output(1, 51) <= input(19);
output(1, 52) <= input(20);
output(1, 53) <= input(21);
output(1, 54) <= input(22);
output(1, 55) <= input(23);
output(1, 56) <= input(24);
output(1, 57) <= input(25);
output(1, 58) <= input(26);
output(1, 59) <= input(27);
output(1, 60) <= input(28);
output(1, 61) <= input(29);
output(1, 62) <= input(30);
output(1, 63) <= input(31);
output(1, 64) <= input(16);
output(1, 65) <= input(17);
output(1, 66) <= input(18);
output(1, 67) <= input(19);
output(1, 68) <= input(20);
output(1, 69) <= input(21);
output(1, 70) <= input(22);
output(1, 71) <= input(23);
output(1, 72) <= input(24);
output(1, 73) <= input(25);
output(1, 74) <= input(26);
output(1, 75) <= input(27);
output(1, 76) <= input(28);
output(1, 77) <= input(29);
output(1, 78) <= input(30);
output(1, 79) <= input(31);
output(1, 80) <= input(32);
output(1, 81) <= input(0);
output(1, 82) <= input(1);
output(1, 83) <= input(2);
output(1, 84) <= input(3);
output(1, 85) <= input(4);
output(1, 86) <= input(5);
output(1, 87) <= input(6);
output(1, 88) <= input(7);
output(1, 89) <= input(8);
output(1, 90) <= input(9);
output(1, 91) <= input(10);
output(1, 92) <= input(11);
output(1, 93) <= input(12);
output(1, 94) <= input(13);
output(1, 95) <= input(14);
output(1, 96) <= input(32);
output(1, 97) <= input(0);
output(1, 98) <= input(1);
output(1, 99) <= input(2);
output(1, 100) <= input(3);
output(1, 101) <= input(4);
output(1, 102) <= input(5);
output(1, 103) <= input(6);
output(1, 104) <= input(7);
output(1, 105) <= input(8);
output(1, 106) <= input(9);
output(1, 107) <= input(10);
output(1, 108) <= input(11);
output(1, 109) <= input(12);
output(1, 110) <= input(13);
output(1, 111) <= input(14);
output(1, 112) <= input(32);
output(1, 113) <= input(0);
output(1, 114) <= input(1);
output(1, 115) <= input(2);
output(1, 116) <= input(3);
output(1, 117) <= input(4);
output(1, 118) <= input(5);
output(1, 119) <= input(6);
output(1, 120) <= input(7);
output(1, 121) <= input(8);
output(1, 122) <= input(9);
output(1, 123) <= input(10);
output(1, 124) <= input(11);
output(1, 125) <= input(12);
output(1, 126) <= input(13);
output(1, 127) <= input(14);
output(1, 128) <= input(33);
output(1, 129) <= input(16);
output(1, 130) <= input(17);
output(1, 131) <= input(18);
output(1, 132) <= input(19);
output(1, 133) <= input(20);
output(1, 134) <= input(21);
output(1, 135) <= input(22);
output(1, 136) <= input(23);
output(1, 137) <= input(24);
output(1, 138) <= input(25);
output(1, 139) <= input(26);
output(1, 140) <= input(27);
output(1, 141) <= input(28);
output(1, 142) <= input(29);
output(1, 143) <= input(30);
output(1, 144) <= input(33);
output(1, 145) <= input(16);
output(1, 146) <= input(17);
output(1, 147) <= input(18);
output(1, 148) <= input(19);
output(1, 149) <= input(20);
output(1, 150) <= input(21);
output(1, 151) <= input(22);
output(1, 152) <= input(23);
output(1, 153) <= input(24);
output(1, 154) <= input(25);
output(1, 155) <= input(26);
output(1, 156) <= input(27);
output(1, 157) <= input(28);
output(1, 158) <= input(29);
output(1, 159) <= input(30);
output(1, 160) <= input(34);
output(1, 161) <= input(32);
output(1, 162) <= input(0);
output(1, 163) <= input(1);
output(1, 164) <= input(2);
output(1, 165) <= input(3);
output(1, 166) <= input(4);
output(1, 167) <= input(5);
output(1, 168) <= input(6);
output(1, 169) <= input(7);
output(1, 170) <= input(8);
output(1, 171) <= input(9);
output(1, 172) <= input(10);
output(1, 173) <= input(11);
output(1, 174) <= input(12);
output(1, 175) <= input(13);
output(1, 176) <= input(34);
output(1, 177) <= input(32);
output(1, 178) <= input(0);
output(1, 179) <= input(1);
output(1, 180) <= input(2);
output(1, 181) <= input(3);
output(1, 182) <= input(4);
output(1, 183) <= input(5);
output(1, 184) <= input(6);
output(1, 185) <= input(7);
output(1, 186) <= input(8);
output(1, 187) <= input(9);
output(1, 188) <= input(10);
output(1, 189) <= input(11);
output(1, 190) <= input(12);
output(1, 191) <= input(13);
output(1, 192) <= input(34);
output(1, 193) <= input(32);
output(1, 194) <= input(0);
output(1, 195) <= input(1);
output(1, 196) <= input(2);
output(1, 197) <= input(3);
output(1, 198) <= input(4);
output(1, 199) <= input(5);
output(1, 200) <= input(6);
output(1, 201) <= input(7);
output(1, 202) <= input(8);
output(1, 203) <= input(9);
output(1, 204) <= input(10);
output(1, 205) <= input(11);
output(1, 206) <= input(12);
output(1, 207) <= input(13);
output(1, 208) <= input(35);
output(1, 209) <= input(33);
output(1, 210) <= input(16);
output(1, 211) <= input(17);
output(1, 212) <= input(18);
output(1, 213) <= input(19);
output(1, 214) <= input(20);
output(1, 215) <= input(21);
output(1, 216) <= input(22);
output(1, 217) <= input(23);
output(1, 218) <= input(24);
output(1, 219) <= input(25);
output(1, 220) <= input(26);
output(1, 221) <= input(27);
output(1, 222) <= input(28);
output(1, 223) <= input(29);
output(1, 224) <= input(35);
output(1, 225) <= input(33);
output(1, 226) <= input(16);
output(1, 227) <= input(17);
output(1, 228) <= input(18);
output(1, 229) <= input(19);
output(1, 230) <= input(20);
output(1, 231) <= input(21);
output(1, 232) <= input(22);
output(1, 233) <= input(23);
output(1, 234) <= input(24);
output(1, 235) <= input(25);
output(1, 236) <= input(26);
output(1, 237) <= input(27);
output(1, 238) <= input(28);
output(1, 239) <= input(29);
output(1, 240) <= input(35);
output(1, 241) <= input(33);
output(1, 242) <= input(16);
output(1, 243) <= input(17);
output(1, 244) <= input(18);
output(1, 245) <= input(19);
output(1, 246) <= input(20);
output(1, 247) <= input(21);
output(1, 248) <= input(22);
output(1, 249) <= input(23);
output(1, 250) <= input(24);
output(1, 251) <= input(25);
output(1, 252) <= input(26);
output(1, 253) <= input(27);
output(1, 254) <= input(28);
output(1, 255) <= input(29);
output(2, 0) <= input(0);
output(2, 1) <= input(1);
output(2, 2) <= input(2);
output(2, 3) <= input(3);
output(2, 4) <= input(4);
output(2, 5) <= input(5);
output(2, 6) <= input(6);
output(2, 7) <= input(7);
output(2, 8) <= input(8);
output(2, 9) <= input(9);
output(2, 10) <= input(10);
output(2, 11) <= input(11);
output(2, 12) <= input(12);
output(2, 13) <= input(13);
output(2, 14) <= input(14);
output(2, 15) <= input(15);
output(2, 16) <= input(0);
output(2, 17) <= input(1);
output(2, 18) <= input(2);
output(2, 19) <= input(3);
output(2, 20) <= input(4);
output(2, 21) <= input(5);
output(2, 22) <= input(6);
output(2, 23) <= input(7);
output(2, 24) <= input(8);
output(2, 25) <= input(9);
output(2, 26) <= input(10);
output(2, 27) <= input(11);
output(2, 28) <= input(12);
output(2, 29) <= input(13);
output(2, 30) <= input(14);
output(2, 31) <= input(15);
output(2, 32) <= input(0);
output(2, 33) <= input(1);
output(2, 34) <= input(2);
output(2, 35) <= input(3);
output(2, 36) <= input(4);
output(2, 37) <= input(5);
output(2, 38) <= input(6);
output(2, 39) <= input(7);
output(2, 40) <= input(8);
output(2, 41) <= input(9);
output(2, 42) <= input(10);
output(2, 43) <= input(11);
output(2, 44) <= input(12);
output(2, 45) <= input(13);
output(2, 46) <= input(14);
output(2, 47) <= input(15);
output(2, 48) <= input(0);
output(2, 49) <= input(1);
output(2, 50) <= input(2);
output(2, 51) <= input(3);
output(2, 52) <= input(4);
output(2, 53) <= input(5);
output(2, 54) <= input(6);
output(2, 55) <= input(7);
output(2, 56) <= input(8);
output(2, 57) <= input(9);
output(2, 58) <= input(10);
output(2, 59) <= input(11);
output(2, 60) <= input(12);
output(2, 61) <= input(13);
output(2, 62) <= input(14);
output(2, 63) <= input(15);
output(2, 64) <= input(16);
output(2, 65) <= input(17);
output(2, 66) <= input(18);
output(2, 67) <= input(19);
output(2, 68) <= input(20);
output(2, 69) <= input(21);
output(2, 70) <= input(22);
output(2, 71) <= input(23);
output(2, 72) <= input(24);
output(2, 73) <= input(25);
output(2, 74) <= input(26);
output(2, 75) <= input(27);
output(2, 76) <= input(28);
output(2, 77) <= input(29);
output(2, 78) <= input(30);
output(2, 79) <= input(31);
output(2, 80) <= input(16);
output(2, 81) <= input(17);
output(2, 82) <= input(18);
output(2, 83) <= input(19);
output(2, 84) <= input(20);
output(2, 85) <= input(21);
output(2, 86) <= input(22);
output(2, 87) <= input(23);
output(2, 88) <= input(24);
output(2, 89) <= input(25);
output(2, 90) <= input(26);
output(2, 91) <= input(27);
output(2, 92) <= input(28);
output(2, 93) <= input(29);
output(2, 94) <= input(30);
output(2, 95) <= input(31);
output(2, 96) <= input(16);
output(2, 97) <= input(17);
output(2, 98) <= input(18);
output(2, 99) <= input(19);
output(2, 100) <= input(20);
output(2, 101) <= input(21);
output(2, 102) <= input(22);
output(2, 103) <= input(23);
output(2, 104) <= input(24);
output(2, 105) <= input(25);
output(2, 106) <= input(26);
output(2, 107) <= input(27);
output(2, 108) <= input(28);
output(2, 109) <= input(29);
output(2, 110) <= input(30);
output(2, 111) <= input(31);
output(2, 112) <= input(16);
output(2, 113) <= input(17);
output(2, 114) <= input(18);
output(2, 115) <= input(19);
output(2, 116) <= input(20);
output(2, 117) <= input(21);
output(2, 118) <= input(22);
output(2, 119) <= input(23);
output(2, 120) <= input(24);
output(2, 121) <= input(25);
output(2, 122) <= input(26);
output(2, 123) <= input(27);
output(2, 124) <= input(28);
output(2, 125) <= input(29);
output(2, 126) <= input(30);
output(2, 127) <= input(31);
output(2, 128) <= input(32);
output(2, 129) <= input(0);
output(2, 130) <= input(1);
output(2, 131) <= input(2);
output(2, 132) <= input(3);
output(2, 133) <= input(4);
output(2, 134) <= input(5);
output(2, 135) <= input(6);
output(2, 136) <= input(7);
output(2, 137) <= input(8);
output(2, 138) <= input(9);
output(2, 139) <= input(10);
output(2, 140) <= input(11);
output(2, 141) <= input(12);
output(2, 142) <= input(13);
output(2, 143) <= input(14);
output(2, 144) <= input(32);
output(2, 145) <= input(0);
output(2, 146) <= input(1);
output(2, 147) <= input(2);
output(2, 148) <= input(3);
output(2, 149) <= input(4);
output(2, 150) <= input(5);
output(2, 151) <= input(6);
output(2, 152) <= input(7);
output(2, 153) <= input(8);
output(2, 154) <= input(9);
output(2, 155) <= input(10);
output(2, 156) <= input(11);
output(2, 157) <= input(12);
output(2, 158) <= input(13);
output(2, 159) <= input(14);
output(2, 160) <= input(32);
output(2, 161) <= input(0);
output(2, 162) <= input(1);
output(2, 163) <= input(2);
output(2, 164) <= input(3);
output(2, 165) <= input(4);
output(2, 166) <= input(5);
output(2, 167) <= input(6);
output(2, 168) <= input(7);
output(2, 169) <= input(8);
output(2, 170) <= input(9);
output(2, 171) <= input(10);
output(2, 172) <= input(11);
output(2, 173) <= input(12);
output(2, 174) <= input(13);
output(2, 175) <= input(14);
output(2, 176) <= input(32);
output(2, 177) <= input(0);
output(2, 178) <= input(1);
output(2, 179) <= input(2);
output(2, 180) <= input(3);
output(2, 181) <= input(4);
output(2, 182) <= input(5);
output(2, 183) <= input(6);
output(2, 184) <= input(7);
output(2, 185) <= input(8);
output(2, 186) <= input(9);
output(2, 187) <= input(10);
output(2, 188) <= input(11);
output(2, 189) <= input(12);
output(2, 190) <= input(13);
output(2, 191) <= input(14);
output(2, 192) <= input(33);
output(2, 193) <= input(16);
output(2, 194) <= input(17);
output(2, 195) <= input(18);
output(2, 196) <= input(19);
output(2, 197) <= input(20);
output(2, 198) <= input(21);
output(2, 199) <= input(22);
output(2, 200) <= input(23);
output(2, 201) <= input(24);
output(2, 202) <= input(25);
output(2, 203) <= input(26);
output(2, 204) <= input(27);
output(2, 205) <= input(28);
output(2, 206) <= input(29);
output(2, 207) <= input(30);
output(2, 208) <= input(33);
output(2, 209) <= input(16);
output(2, 210) <= input(17);
output(2, 211) <= input(18);
output(2, 212) <= input(19);
output(2, 213) <= input(20);
output(2, 214) <= input(21);
output(2, 215) <= input(22);
output(2, 216) <= input(23);
output(2, 217) <= input(24);
output(2, 218) <= input(25);
output(2, 219) <= input(26);
output(2, 220) <= input(27);
output(2, 221) <= input(28);
output(2, 222) <= input(29);
output(2, 223) <= input(30);
output(2, 224) <= input(33);
output(2, 225) <= input(16);
output(2, 226) <= input(17);
output(2, 227) <= input(18);
output(2, 228) <= input(19);
output(2, 229) <= input(20);
output(2, 230) <= input(21);
output(2, 231) <= input(22);
output(2, 232) <= input(23);
output(2, 233) <= input(24);
output(2, 234) <= input(25);
output(2, 235) <= input(26);
output(2, 236) <= input(27);
output(2, 237) <= input(28);
output(2, 238) <= input(29);
output(2, 239) <= input(30);
output(2, 240) <= input(33);
output(2, 241) <= input(16);
output(2, 242) <= input(17);
output(2, 243) <= input(18);
output(2, 244) <= input(19);
output(2, 245) <= input(20);
output(2, 246) <= input(21);
output(2, 247) <= input(22);
output(2, 248) <= input(23);
output(2, 249) <= input(24);
output(2, 250) <= input(25);
output(2, 251) <= input(26);
output(2, 252) <= input(27);
output(2, 253) <= input(28);
output(2, 254) <= input(29);
output(2, 255) <= input(30);
when "1101" =>
output(0, 0) <= input(0);
output(0, 1) <= input(1);
output(0, 2) <= input(2);
output(0, 3) <= input(3);
output(0, 4) <= input(4);
output(0, 5) <= input(5);
output(0, 6) <= input(6);
output(0, 7) <= input(7);
output(0, 8) <= input(8);
output(0, 9) <= input(9);
output(0, 10) <= input(10);
output(0, 11) <= input(11);
output(0, 12) <= input(12);
output(0, 13) <= input(13);
output(0, 14) <= input(14);
output(0, 15) <= input(15);
output(0, 16) <= input(0);
output(0, 17) <= input(1);
output(0, 18) <= input(2);
output(0, 19) <= input(3);
output(0, 20) <= input(4);
output(0, 21) <= input(5);
output(0, 22) <= input(6);
output(0, 23) <= input(7);
output(0, 24) <= input(8);
output(0, 25) <= input(9);
output(0, 26) <= input(10);
output(0, 27) <= input(11);
output(0, 28) <= input(12);
output(0, 29) <= input(13);
output(0, 30) <= input(14);
output(0, 31) <= input(15);
output(0, 32) <= input(0);
output(0, 33) <= input(1);
output(0, 34) <= input(2);
output(0, 35) <= input(3);
output(0, 36) <= input(4);
output(0, 37) <= input(5);
output(0, 38) <= input(6);
output(0, 39) <= input(7);
output(0, 40) <= input(8);
output(0, 41) <= input(9);
output(0, 42) <= input(10);
output(0, 43) <= input(11);
output(0, 44) <= input(12);
output(0, 45) <= input(13);
output(0, 46) <= input(14);
output(0, 47) <= input(15);
output(0, 48) <= input(0);
output(0, 49) <= input(1);
output(0, 50) <= input(2);
output(0, 51) <= input(3);
output(0, 52) <= input(4);
output(0, 53) <= input(5);
output(0, 54) <= input(6);
output(0, 55) <= input(7);
output(0, 56) <= input(8);
output(0, 57) <= input(9);
output(0, 58) <= input(10);
output(0, 59) <= input(11);
output(0, 60) <= input(12);
output(0, 61) <= input(13);
output(0, 62) <= input(14);
output(0, 63) <= input(15);
output(0, 64) <= input(0);
output(0, 65) <= input(1);
output(0, 66) <= input(2);
output(0, 67) <= input(3);
output(0, 68) <= input(4);
output(0, 69) <= input(5);
output(0, 70) <= input(6);
output(0, 71) <= input(7);
output(0, 72) <= input(8);
output(0, 73) <= input(9);
output(0, 74) <= input(10);
output(0, 75) <= input(11);
output(0, 76) <= input(12);
output(0, 77) <= input(13);
output(0, 78) <= input(14);
output(0, 79) <= input(15);
output(0, 80) <= input(16);
output(0, 81) <= input(17);
output(0, 82) <= input(18);
output(0, 83) <= input(19);
output(0, 84) <= input(20);
output(0, 85) <= input(21);
output(0, 86) <= input(22);
output(0, 87) <= input(23);
output(0, 88) <= input(24);
output(0, 89) <= input(25);
output(0, 90) <= input(26);
output(0, 91) <= input(27);
output(0, 92) <= input(28);
output(0, 93) <= input(29);
output(0, 94) <= input(30);
output(0, 95) <= input(31);
output(0, 96) <= input(16);
output(0, 97) <= input(17);
output(0, 98) <= input(18);
output(0, 99) <= input(19);
output(0, 100) <= input(20);
output(0, 101) <= input(21);
output(0, 102) <= input(22);
output(0, 103) <= input(23);
output(0, 104) <= input(24);
output(0, 105) <= input(25);
output(0, 106) <= input(26);
output(0, 107) <= input(27);
output(0, 108) <= input(28);
output(0, 109) <= input(29);
output(0, 110) <= input(30);
output(0, 111) <= input(31);
output(0, 112) <= input(16);
output(0, 113) <= input(17);
output(0, 114) <= input(18);
output(0, 115) <= input(19);
output(0, 116) <= input(20);
output(0, 117) <= input(21);
output(0, 118) <= input(22);
output(0, 119) <= input(23);
output(0, 120) <= input(24);
output(0, 121) <= input(25);
output(0, 122) <= input(26);
output(0, 123) <= input(27);
output(0, 124) <= input(28);
output(0, 125) <= input(29);
output(0, 126) <= input(30);
output(0, 127) <= input(31);
output(0, 128) <= input(16);
output(0, 129) <= input(17);
output(0, 130) <= input(18);
output(0, 131) <= input(19);
output(0, 132) <= input(20);
output(0, 133) <= input(21);
output(0, 134) <= input(22);
output(0, 135) <= input(23);
output(0, 136) <= input(24);
output(0, 137) <= input(25);
output(0, 138) <= input(26);
output(0, 139) <= input(27);
output(0, 140) <= input(28);
output(0, 141) <= input(29);
output(0, 142) <= input(30);
output(0, 143) <= input(31);
output(0, 144) <= input(16);
output(0, 145) <= input(17);
output(0, 146) <= input(18);
output(0, 147) <= input(19);
output(0, 148) <= input(20);
output(0, 149) <= input(21);
output(0, 150) <= input(22);
output(0, 151) <= input(23);
output(0, 152) <= input(24);
output(0, 153) <= input(25);
output(0, 154) <= input(26);
output(0, 155) <= input(27);
output(0, 156) <= input(28);
output(0, 157) <= input(29);
output(0, 158) <= input(30);
output(0, 159) <= input(31);
output(0, 160) <= input(32);
output(0, 161) <= input(0);
output(0, 162) <= input(1);
output(0, 163) <= input(2);
output(0, 164) <= input(3);
output(0, 165) <= input(4);
output(0, 166) <= input(5);
output(0, 167) <= input(6);
output(0, 168) <= input(7);
output(0, 169) <= input(8);
output(0, 170) <= input(9);
output(0, 171) <= input(10);
output(0, 172) <= input(11);
output(0, 173) <= input(12);
output(0, 174) <= input(13);
output(0, 175) <= input(14);
output(0, 176) <= input(32);
output(0, 177) <= input(0);
output(0, 178) <= input(1);
output(0, 179) <= input(2);
output(0, 180) <= input(3);
output(0, 181) <= input(4);
output(0, 182) <= input(5);
output(0, 183) <= input(6);
output(0, 184) <= input(7);
output(0, 185) <= input(8);
output(0, 186) <= input(9);
output(0, 187) <= input(10);
output(0, 188) <= input(11);
output(0, 189) <= input(12);
output(0, 190) <= input(13);
output(0, 191) <= input(14);
output(0, 192) <= input(32);
output(0, 193) <= input(0);
output(0, 194) <= input(1);
output(0, 195) <= input(2);
output(0, 196) <= input(3);
output(0, 197) <= input(4);
output(0, 198) <= input(5);
output(0, 199) <= input(6);
output(0, 200) <= input(7);
output(0, 201) <= input(8);
output(0, 202) <= input(9);
output(0, 203) <= input(10);
output(0, 204) <= input(11);
output(0, 205) <= input(12);
output(0, 206) <= input(13);
output(0, 207) <= input(14);
output(0, 208) <= input(32);
output(0, 209) <= input(0);
output(0, 210) <= input(1);
output(0, 211) <= input(2);
output(0, 212) <= input(3);
output(0, 213) <= input(4);
output(0, 214) <= input(5);
output(0, 215) <= input(6);
output(0, 216) <= input(7);
output(0, 217) <= input(8);
output(0, 218) <= input(9);
output(0, 219) <= input(10);
output(0, 220) <= input(11);
output(0, 221) <= input(12);
output(0, 222) <= input(13);
output(0, 223) <= input(14);
output(0, 224) <= input(32);
output(0, 225) <= input(0);
output(0, 226) <= input(1);
output(0, 227) <= input(2);
output(0, 228) <= input(3);
output(0, 229) <= input(4);
output(0, 230) <= input(5);
output(0, 231) <= input(6);
output(0, 232) <= input(7);
output(0, 233) <= input(8);
output(0, 234) <= input(9);
output(0, 235) <= input(10);
output(0, 236) <= input(11);
output(0, 237) <= input(12);
output(0, 238) <= input(13);
output(0, 239) <= input(14);
output(0, 240) <= input(32);
output(0, 241) <= input(0);
output(0, 242) <= input(1);
output(0, 243) <= input(2);
output(0, 244) <= input(3);
output(0, 245) <= input(4);
output(0, 246) <= input(5);
output(0, 247) <= input(6);
output(0, 248) <= input(7);
output(0, 249) <= input(8);
output(0, 250) <= input(9);
output(0, 251) <= input(10);
output(0, 252) <= input(11);
output(0, 253) <= input(12);
output(0, 254) <= input(13);
output(0, 255) <= input(14);
output(1, 0) <= input(0);
output(1, 1) <= input(1);
output(1, 2) <= input(2);
output(1, 3) <= input(3);
output(1, 4) <= input(4);
output(1, 5) <= input(5);
output(1, 6) <= input(6);
output(1, 7) <= input(7);
output(1, 8) <= input(8);
output(1, 9) <= input(9);
output(1, 10) <= input(10);
output(1, 11) <= input(11);
output(1, 12) <= input(12);
output(1, 13) <= input(13);
output(1, 14) <= input(14);
output(1, 15) <= input(15);
output(1, 16) <= input(0);
output(1, 17) <= input(1);
output(1, 18) <= input(2);
output(1, 19) <= input(3);
output(1, 20) <= input(4);
output(1, 21) <= input(5);
output(1, 22) <= input(6);
output(1, 23) <= input(7);
output(1, 24) <= input(8);
output(1, 25) <= input(9);
output(1, 26) <= input(10);
output(1, 27) <= input(11);
output(1, 28) <= input(12);
output(1, 29) <= input(13);
output(1, 30) <= input(14);
output(1, 31) <= input(15);
output(1, 32) <= input(0);
output(1, 33) <= input(1);
output(1, 34) <= input(2);
output(1, 35) <= input(3);
output(1, 36) <= input(4);
output(1, 37) <= input(5);
output(1, 38) <= input(6);
output(1, 39) <= input(7);
output(1, 40) <= input(8);
output(1, 41) <= input(9);
output(1, 42) <= input(10);
output(1, 43) <= input(11);
output(1, 44) <= input(12);
output(1, 45) <= input(13);
output(1, 46) <= input(14);
output(1, 47) <= input(15);
output(1, 48) <= input(0);
output(1, 49) <= input(1);
output(1, 50) <= input(2);
output(1, 51) <= input(3);
output(1, 52) <= input(4);
output(1, 53) <= input(5);
output(1, 54) <= input(6);
output(1, 55) <= input(7);
output(1, 56) <= input(8);
output(1, 57) <= input(9);
output(1, 58) <= input(10);
output(1, 59) <= input(11);
output(1, 60) <= input(12);
output(1, 61) <= input(13);
output(1, 62) <= input(14);
output(1, 63) <= input(15);
output(1, 64) <= input(0);
output(1, 65) <= input(1);
output(1, 66) <= input(2);
output(1, 67) <= input(3);
output(1, 68) <= input(4);
output(1, 69) <= input(5);
output(1, 70) <= input(6);
output(1, 71) <= input(7);
output(1, 72) <= input(8);
output(1, 73) <= input(9);
output(1, 74) <= input(10);
output(1, 75) <= input(11);
output(1, 76) <= input(12);
output(1, 77) <= input(13);
output(1, 78) <= input(14);
output(1, 79) <= input(15);
output(1, 80) <= input(0);
output(1, 81) <= input(1);
output(1, 82) <= input(2);
output(1, 83) <= input(3);
output(1, 84) <= input(4);
output(1, 85) <= input(5);
output(1, 86) <= input(6);
output(1, 87) <= input(7);
output(1, 88) <= input(8);
output(1, 89) <= input(9);
output(1, 90) <= input(10);
output(1, 91) <= input(11);
output(1, 92) <= input(12);
output(1, 93) <= input(13);
output(1, 94) <= input(14);
output(1, 95) <= input(15);
output(1, 96) <= input(0);
output(1, 97) <= input(1);
output(1, 98) <= input(2);
output(1, 99) <= input(3);
output(1, 100) <= input(4);
output(1, 101) <= input(5);
output(1, 102) <= input(6);
output(1, 103) <= input(7);
output(1, 104) <= input(8);
output(1, 105) <= input(9);
output(1, 106) <= input(10);
output(1, 107) <= input(11);
output(1, 108) <= input(12);
output(1, 109) <= input(13);
output(1, 110) <= input(14);
output(1, 111) <= input(15);
output(1, 112) <= input(0);
output(1, 113) <= input(1);
output(1, 114) <= input(2);
output(1, 115) <= input(3);
output(1, 116) <= input(4);
output(1, 117) <= input(5);
output(1, 118) <= input(6);
output(1, 119) <= input(7);
output(1, 120) <= input(8);
output(1, 121) <= input(9);
output(1, 122) <= input(10);
output(1, 123) <= input(11);
output(1, 124) <= input(12);
output(1, 125) <= input(13);
output(1, 126) <= input(14);
output(1, 127) <= input(15);
output(1, 128) <= input(16);
output(1, 129) <= input(17);
output(1, 130) <= input(18);
output(1, 131) <= input(19);
output(1, 132) <= input(20);
output(1, 133) <= input(21);
output(1, 134) <= input(22);
output(1, 135) <= input(23);
output(1, 136) <= input(24);
output(1, 137) <= input(25);
output(1, 138) <= input(26);
output(1, 139) <= input(27);
output(1, 140) <= input(28);
output(1, 141) <= input(29);
output(1, 142) <= input(30);
output(1, 143) <= input(31);
output(1, 144) <= input(16);
output(1, 145) <= input(17);
output(1, 146) <= input(18);
output(1, 147) <= input(19);
output(1, 148) <= input(20);
output(1, 149) <= input(21);
output(1, 150) <= input(22);
output(1, 151) <= input(23);
output(1, 152) <= input(24);
output(1, 153) <= input(25);
output(1, 154) <= input(26);
output(1, 155) <= input(27);
output(1, 156) <= input(28);
output(1, 157) <= input(29);
output(1, 158) <= input(30);
output(1, 159) <= input(31);
output(1, 160) <= input(16);
output(1, 161) <= input(17);
output(1, 162) <= input(18);
output(1, 163) <= input(19);
output(1, 164) <= input(20);
output(1, 165) <= input(21);
output(1, 166) <= input(22);
output(1, 167) <= input(23);
output(1, 168) <= input(24);
output(1, 169) <= input(25);
output(1, 170) <= input(26);
output(1, 171) <= input(27);
output(1, 172) <= input(28);
output(1, 173) <= input(29);
output(1, 174) <= input(30);
output(1, 175) <= input(31);
output(1, 176) <= input(16);
output(1, 177) <= input(17);
output(1, 178) <= input(18);
output(1, 179) <= input(19);
output(1, 180) <= input(20);
output(1, 181) <= input(21);
output(1, 182) <= input(22);
output(1, 183) <= input(23);
output(1, 184) <= input(24);
output(1, 185) <= input(25);
output(1, 186) <= input(26);
output(1, 187) <= input(27);
output(1, 188) <= input(28);
output(1, 189) <= input(29);
output(1, 190) <= input(30);
output(1, 191) <= input(31);
output(1, 192) <= input(16);
output(1, 193) <= input(17);
output(1, 194) <= input(18);
output(1, 195) <= input(19);
output(1, 196) <= input(20);
output(1, 197) <= input(21);
output(1, 198) <= input(22);
output(1, 199) <= input(23);
output(1, 200) <= input(24);
output(1, 201) <= input(25);
output(1, 202) <= input(26);
output(1, 203) <= input(27);
output(1, 204) <= input(28);
output(1, 205) <= input(29);
output(1, 206) <= input(30);
output(1, 207) <= input(31);
output(1, 208) <= input(16);
output(1, 209) <= input(17);
output(1, 210) <= input(18);
output(1, 211) <= input(19);
output(1, 212) <= input(20);
output(1, 213) <= input(21);
output(1, 214) <= input(22);
output(1, 215) <= input(23);
output(1, 216) <= input(24);
output(1, 217) <= input(25);
output(1, 218) <= input(26);
output(1, 219) <= input(27);
output(1, 220) <= input(28);
output(1, 221) <= input(29);
output(1, 222) <= input(30);
output(1, 223) <= input(31);
output(1, 224) <= input(16);
output(1, 225) <= input(17);
output(1, 226) <= input(18);
output(1, 227) <= input(19);
output(1, 228) <= input(20);
output(1, 229) <= input(21);
output(1, 230) <= input(22);
output(1, 231) <= input(23);
output(1, 232) <= input(24);
output(1, 233) <= input(25);
output(1, 234) <= input(26);
output(1, 235) <= input(27);
output(1, 236) <= input(28);
output(1, 237) <= input(29);
output(1, 238) <= input(30);
output(1, 239) <= input(31);
output(1, 240) <= input(16);
output(1, 241) <= input(17);
output(1, 242) <= input(18);
output(1, 243) <= input(19);
output(1, 244) <= input(20);
output(1, 245) <= input(21);
output(1, 246) <= input(22);
output(1, 247) <= input(23);
output(1, 248) <= input(24);
output(1, 249) <= input(25);
output(1, 250) <= input(26);
output(1, 251) <= input(27);
output(1, 252) <= input(28);
output(1, 253) <= input(29);
output(1, 254) <= input(30);
output(1, 255) <= input(31);
output(2, 0) <= input(0);
output(2, 1) <= input(1);
output(2, 2) <= input(2);
output(2, 3) <= input(3);
output(2, 4) <= input(4);
output(2, 5) <= input(5);
output(2, 6) <= input(6);
output(2, 7) <= input(7);
output(2, 8) <= input(8);
output(2, 9) <= input(9);
output(2, 10) <= input(10);
output(2, 11) <= input(11);
output(2, 12) <= input(12);
output(2, 13) <= input(13);
output(2, 14) <= input(14);
output(2, 15) <= input(15);
output(2, 16) <= input(0);
output(2, 17) <= input(1);
output(2, 18) <= input(2);
output(2, 19) <= input(3);
output(2, 20) <= input(4);
output(2, 21) <= input(5);
output(2, 22) <= input(6);
output(2, 23) <= input(7);
output(2, 24) <= input(8);
output(2, 25) <= input(9);
output(2, 26) <= input(10);
output(2, 27) <= input(11);
output(2, 28) <= input(12);
output(2, 29) <= input(13);
output(2, 30) <= input(14);
output(2, 31) <= input(15);
output(2, 32) <= input(0);
output(2, 33) <= input(1);
output(2, 34) <= input(2);
output(2, 35) <= input(3);
output(2, 36) <= input(4);
output(2, 37) <= input(5);
output(2, 38) <= input(6);
output(2, 39) <= input(7);
output(2, 40) <= input(8);
output(2, 41) <= input(9);
output(2, 42) <= input(10);
output(2, 43) <= input(11);
output(2, 44) <= input(12);
output(2, 45) <= input(13);
output(2, 46) <= input(14);
output(2, 47) <= input(15);
output(2, 48) <= input(0);
output(2, 49) <= input(1);
output(2, 50) <= input(2);
output(2, 51) <= input(3);
output(2, 52) <= input(4);
output(2, 53) <= input(5);
output(2, 54) <= input(6);
output(2, 55) <= input(7);
output(2, 56) <= input(8);
output(2, 57) <= input(9);
output(2, 58) <= input(10);
output(2, 59) <= input(11);
output(2, 60) <= input(12);
output(2, 61) <= input(13);
output(2, 62) <= input(14);
output(2, 63) <= input(15);
output(2, 64) <= input(0);
output(2, 65) <= input(1);
output(2, 66) <= input(2);
output(2, 67) <= input(3);
output(2, 68) <= input(4);
output(2, 69) <= input(5);
output(2, 70) <= input(6);
output(2, 71) <= input(7);
output(2, 72) <= input(8);
output(2, 73) <= input(9);
output(2, 74) <= input(10);
output(2, 75) <= input(11);
output(2, 76) <= input(12);
output(2, 77) <= input(13);
output(2, 78) <= input(14);
output(2, 79) <= input(15);
output(2, 80) <= input(0);
output(2, 81) <= input(1);
output(2, 82) <= input(2);
output(2, 83) <= input(3);
output(2, 84) <= input(4);
output(2, 85) <= input(5);
output(2, 86) <= input(6);
output(2, 87) <= input(7);
output(2, 88) <= input(8);
output(2, 89) <= input(9);
output(2, 90) <= input(10);
output(2, 91) <= input(11);
output(2, 92) <= input(12);
output(2, 93) <= input(13);
output(2, 94) <= input(14);
output(2, 95) <= input(15);
output(2, 96) <= input(0);
output(2, 97) <= input(1);
output(2, 98) <= input(2);
output(2, 99) <= input(3);
output(2, 100) <= input(4);
output(2, 101) <= input(5);
output(2, 102) <= input(6);
output(2, 103) <= input(7);
output(2, 104) <= input(8);
output(2, 105) <= input(9);
output(2, 106) <= input(10);
output(2, 107) <= input(11);
output(2, 108) <= input(12);
output(2, 109) <= input(13);
output(2, 110) <= input(14);
output(2, 111) <= input(15);
output(2, 112) <= input(0);
output(2, 113) <= input(1);
output(2, 114) <= input(2);
output(2, 115) <= input(3);
output(2, 116) <= input(4);
output(2, 117) <= input(5);
output(2, 118) <= input(6);
output(2, 119) <= input(7);
output(2, 120) <= input(8);
output(2, 121) <= input(9);
output(2, 122) <= input(10);
output(2, 123) <= input(11);
output(2, 124) <= input(12);
output(2, 125) <= input(13);
output(2, 126) <= input(14);
output(2, 127) <= input(15);
output(2, 128) <= input(0);
output(2, 129) <= input(1);
output(2, 130) <= input(2);
output(2, 131) <= input(3);
output(2, 132) <= input(4);
output(2, 133) <= input(5);
output(2, 134) <= input(6);
output(2, 135) <= input(7);
output(2, 136) <= input(8);
output(2, 137) <= input(9);
output(2, 138) <= input(10);
output(2, 139) <= input(11);
output(2, 140) <= input(12);
output(2, 141) <= input(13);
output(2, 142) <= input(14);
output(2, 143) <= input(15);
output(2, 144) <= input(0);
output(2, 145) <= input(1);
output(2, 146) <= input(2);
output(2, 147) <= input(3);
output(2, 148) <= input(4);
output(2, 149) <= input(5);
output(2, 150) <= input(6);
output(2, 151) <= input(7);
output(2, 152) <= input(8);
output(2, 153) <= input(9);
output(2, 154) <= input(10);
output(2, 155) <= input(11);
output(2, 156) <= input(12);
output(2, 157) <= input(13);
output(2, 158) <= input(14);
output(2, 159) <= input(15);
output(2, 160) <= input(0);
output(2, 161) <= input(1);
output(2, 162) <= input(2);
output(2, 163) <= input(3);
output(2, 164) <= input(4);
output(2, 165) <= input(5);
output(2, 166) <= input(6);
output(2, 167) <= input(7);
output(2, 168) <= input(8);
output(2, 169) <= input(9);
output(2, 170) <= input(10);
output(2, 171) <= input(11);
output(2, 172) <= input(12);
output(2, 173) <= input(13);
output(2, 174) <= input(14);
output(2, 175) <= input(15);
output(2, 176) <= input(0);
output(2, 177) <= input(1);
output(2, 178) <= input(2);
output(2, 179) <= input(3);
output(2, 180) <= input(4);
output(2, 181) <= input(5);
output(2, 182) <= input(6);
output(2, 183) <= input(7);
output(2, 184) <= input(8);
output(2, 185) <= input(9);
output(2, 186) <= input(10);
output(2, 187) <= input(11);
output(2, 188) <= input(12);
output(2, 189) <= input(13);
output(2, 190) <= input(14);
output(2, 191) <= input(15);
output(2, 192) <= input(0);
output(2, 193) <= input(1);
output(2, 194) <= input(2);
output(2, 195) <= input(3);
output(2, 196) <= input(4);
output(2, 197) <= input(5);
output(2, 198) <= input(6);
output(2, 199) <= input(7);
output(2, 200) <= input(8);
output(2, 201) <= input(9);
output(2, 202) <= input(10);
output(2, 203) <= input(11);
output(2, 204) <= input(12);
output(2, 205) <= input(13);
output(2, 206) <= input(14);
output(2, 207) <= input(15);
output(2, 208) <= input(0);
output(2, 209) <= input(1);
output(2, 210) <= input(2);
output(2, 211) <= input(3);
output(2, 212) <= input(4);
output(2, 213) <= input(5);
output(2, 214) <= input(6);
output(2, 215) <= input(7);
output(2, 216) <= input(8);
output(2, 217) <= input(9);
output(2, 218) <= input(10);
output(2, 219) <= input(11);
output(2, 220) <= input(12);
output(2, 221) <= input(13);
output(2, 222) <= input(14);
output(2, 223) <= input(15);
output(2, 224) <= input(0);
output(2, 225) <= input(1);
output(2, 226) <= input(2);
output(2, 227) <= input(3);
output(2, 228) <= input(4);
output(2, 229) <= input(5);
output(2, 230) <= input(6);
output(2, 231) <= input(7);
output(2, 232) <= input(8);
output(2, 233) <= input(9);
output(2, 234) <= input(10);
output(2, 235) <= input(11);
output(2, 236) <= input(12);
output(2, 237) <= input(13);
output(2, 238) <= input(14);
output(2, 239) <= input(15);
output(2, 240) <= input(0);
output(2, 241) <= input(1);
output(2, 242) <= input(2);
output(2, 243) <= input(3);
output(2, 244) <= input(4);
output(2, 245) <= input(5);
output(2, 246) <= input(6);
output(2, 247) <= input(7);
output(2, 248) <= input(8);
output(2, 249) <= input(9);
output(2, 250) <= input(10);
output(2, 251) <= input(11);
output(2, 252) <= input(12);
output(2, 253) <= input(13);
output(2, 254) <= input(14);
output(2, 255) <= input(15);
output(3, 0) <= input(17);
output(3, 1) <= input(18);
output(3, 2) <= input(19);
output(3, 3) <= input(20);
output(3, 4) <= input(21);
output(3, 5) <= input(22);
output(3, 6) <= input(23);
output(3, 7) <= input(24);
output(3, 8) <= input(25);
output(3, 9) <= input(26);
output(3, 10) <= input(27);
output(3, 11) <= input(28);
output(3, 12) <= input(29);
output(3, 13) <= input(30);
output(3, 14) <= input(31);
output(3, 15) <= input(33);
output(3, 16) <= input(17);
output(3, 17) <= input(18);
output(3, 18) <= input(19);
output(3, 19) <= input(20);
output(3, 20) <= input(21);
output(3, 21) <= input(22);
output(3, 22) <= input(23);
output(3, 23) <= input(24);
output(3, 24) <= input(25);
output(3, 25) <= input(26);
output(3, 26) <= input(27);
output(3, 27) <= input(28);
output(3, 28) <= input(29);
output(3, 29) <= input(30);
output(3, 30) <= input(31);
output(3, 31) <= input(33);
output(3, 32) <= input(17);
output(3, 33) <= input(18);
output(3, 34) <= input(19);
output(3, 35) <= input(20);
output(3, 36) <= input(21);
output(3, 37) <= input(22);
output(3, 38) <= input(23);
output(3, 39) <= input(24);
output(3, 40) <= input(25);
output(3, 41) <= input(26);
output(3, 42) <= input(27);
output(3, 43) <= input(28);
output(3, 44) <= input(29);
output(3, 45) <= input(30);
output(3, 46) <= input(31);
output(3, 47) <= input(33);
output(3, 48) <= input(17);
output(3, 49) <= input(18);
output(3, 50) <= input(19);
output(3, 51) <= input(20);
output(3, 52) <= input(21);
output(3, 53) <= input(22);
output(3, 54) <= input(23);
output(3, 55) <= input(24);
output(3, 56) <= input(25);
output(3, 57) <= input(26);
output(3, 58) <= input(27);
output(3, 59) <= input(28);
output(3, 60) <= input(29);
output(3, 61) <= input(30);
output(3, 62) <= input(31);
output(3, 63) <= input(33);
output(3, 64) <= input(17);
output(3, 65) <= input(18);
output(3, 66) <= input(19);
output(3, 67) <= input(20);
output(3, 68) <= input(21);
output(3, 69) <= input(22);
output(3, 70) <= input(23);
output(3, 71) <= input(24);
output(3, 72) <= input(25);
output(3, 73) <= input(26);
output(3, 74) <= input(27);
output(3, 75) <= input(28);
output(3, 76) <= input(29);
output(3, 77) <= input(30);
output(3, 78) <= input(31);
output(3, 79) <= input(33);
output(3, 80) <= input(17);
output(3, 81) <= input(18);
output(3, 82) <= input(19);
output(3, 83) <= input(20);
output(3, 84) <= input(21);
output(3, 85) <= input(22);
output(3, 86) <= input(23);
output(3, 87) <= input(24);
output(3, 88) <= input(25);
output(3, 89) <= input(26);
output(3, 90) <= input(27);
output(3, 91) <= input(28);
output(3, 92) <= input(29);
output(3, 93) <= input(30);
output(3, 94) <= input(31);
output(3, 95) <= input(33);
output(3, 96) <= input(17);
output(3, 97) <= input(18);
output(3, 98) <= input(19);
output(3, 99) <= input(20);
output(3, 100) <= input(21);
output(3, 101) <= input(22);
output(3, 102) <= input(23);
output(3, 103) <= input(24);
output(3, 104) <= input(25);
output(3, 105) <= input(26);
output(3, 106) <= input(27);
output(3, 107) <= input(28);
output(3, 108) <= input(29);
output(3, 109) <= input(30);
output(3, 110) <= input(31);
output(3, 111) <= input(33);
output(3, 112) <= input(17);
output(3, 113) <= input(18);
output(3, 114) <= input(19);
output(3, 115) <= input(20);
output(3, 116) <= input(21);
output(3, 117) <= input(22);
output(3, 118) <= input(23);
output(3, 119) <= input(24);
output(3, 120) <= input(25);
output(3, 121) <= input(26);
output(3, 122) <= input(27);
output(3, 123) <= input(28);
output(3, 124) <= input(29);
output(3, 125) <= input(30);
output(3, 126) <= input(31);
output(3, 127) <= input(33);
output(3, 128) <= input(17);
output(3, 129) <= input(18);
output(3, 130) <= input(19);
output(3, 131) <= input(20);
output(3, 132) <= input(21);
output(3, 133) <= input(22);
output(3, 134) <= input(23);
output(3, 135) <= input(24);
output(3, 136) <= input(25);
output(3, 137) <= input(26);
output(3, 138) <= input(27);
output(3, 139) <= input(28);
output(3, 140) <= input(29);
output(3, 141) <= input(30);
output(3, 142) <= input(31);
output(3, 143) <= input(33);
output(3, 144) <= input(17);
output(3, 145) <= input(18);
output(3, 146) <= input(19);
output(3, 147) <= input(20);
output(3, 148) <= input(21);
output(3, 149) <= input(22);
output(3, 150) <= input(23);
output(3, 151) <= input(24);
output(3, 152) <= input(25);
output(3, 153) <= input(26);
output(3, 154) <= input(27);
output(3, 155) <= input(28);
output(3, 156) <= input(29);
output(3, 157) <= input(30);
output(3, 158) <= input(31);
output(3, 159) <= input(33);
output(3, 160) <= input(17);
output(3, 161) <= input(18);
output(3, 162) <= input(19);
output(3, 163) <= input(20);
output(3, 164) <= input(21);
output(3, 165) <= input(22);
output(3, 166) <= input(23);
output(3, 167) <= input(24);
output(3, 168) <= input(25);
output(3, 169) <= input(26);
output(3, 170) <= input(27);
output(3, 171) <= input(28);
output(3, 172) <= input(29);
output(3, 173) <= input(30);
output(3, 174) <= input(31);
output(3, 175) <= input(33);
output(3, 176) <= input(17);
output(3, 177) <= input(18);
output(3, 178) <= input(19);
output(3, 179) <= input(20);
output(3, 180) <= input(21);
output(3, 181) <= input(22);
output(3, 182) <= input(23);
output(3, 183) <= input(24);
output(3, 184) <= input(25);
output(3, 185) <= input(26);
output(3, 186) <= input(27);
output(3, 187) <= input(28);
output(3, 188) <= input(29);
output(3, 189) <= input(30);
output(3, 190) <= input(31);
output(3, 191) <= input(33);
output(3, 192) <= input(17);
output(3, 193) <= input(18);
output(3, 194) <= input(19);
output(3, 195) <= input(20);
output(3, 196) <= input(21);
output(3, 197) <= input(22);
output(3, 198) <= input(23);
output(3, 199) <= input(24);
output(3, 200) <= input(25);
output(3, 201) <= input(26);
output(3, 202) <= input(27);
output(3, 203) <= input(28);
output(3, 204) <= input(29);
output(3, 205) <= input(30);
output(3, 206) <= input(31);
output(3, 207) <= input(33);
output(3, 208) <= input(17);
output(3, 209) <= input(18);
output(3, 210) <= input(19);
output(3, 211) <= input(20);
output(3, 212) <= input(21);
output(3, 213) <= input(22);
output(3, 214) <= input(23);
output(3, 215) <= input(24);
output(3, 216) <= input(25);
output(3, 217) <= input(26);
output(3, 218) <= input(27);
output(3, 219) <= input(28);
output(3, 220) <= input(29);
output(3, 221) <= input(30);
output(3, 222) <= input(31);
output(3, 223) <= input(33);
output(3, 224) <= input(17);
output(3, 225) <= input(18);
output(3, 226) <= input(19);
output(3, 227) <= input(20);
output(3, 228) <= input(21);
output(3, 229) <= input(22);
output(3, 230) <= input(23);
output(3, 231) <= input(24);
output(3, 232) <= input(25);
output(3, 233) <= input(26);
output(3, 234) <= input(27);
output(3, 235) <= input(28);
output(3, 236) <= input(29);
output(3, 237) <= input(30);
output(3, 238) <= input(31);
output(3, 239) <= input(33);
output(3, 240) <= input(17);
output(3, 241) <= input(18);
output(3, 242) <= input(19);
output(3, 243) <= input(20);
output(3, 244) <= input(21);
output(3, 245) <= input(22);
output(3, 246) <= input(23);
output(3, 247) <= input(24);
output(3, 248) <= input(25);
output(3, 249) <= input(26);
output(3, 250) <= input(27);
output(3, 251) <= input(28);
output(3, 252) <= input(29);
output(3, 253) <= input(30);
output(3, 254) <= input(31);
output(3, 255) <= input(33);
output(4, 0) <= input(17);
output(4, 1) <= input(18);
output(4, 2) <= input(19);
output(4, 3) <= input(20);
output(4, 4) <= input(21);
output(4, 5) <= input(22);
output(4, 6) <= input(23);
output(4, 7) <= input(24);
output(4, 8) <= input(25);
output(4, 9) <= input(26);
output(4, 10) <= input(27);
output(4, 11) <= input(28);
output(4, 12) <= input(29);
output(4, 13) <= input(30);
output(4, 14) <= input(31);
output(4, 15) <= input(33);
output(4, 16) <= input(17);
output(4, 17) <= input(18);
output(4, 18) <= input(19);
output(4, 19) <= input(20);
output(4, 20) <= input(21);
output(4, 21) <= input(22);
output(4, 22) <= input(23);
output(4, 23) <= input(24);
output(4, 24) <= input(25);
output(4, 25) <= input(26);
output(4, 26) <= input(27);
output(4, 27) <= input(28);
output(4, 28) <= input(29);
output(4, 29) <= input(30);
output(4, 30) <= input(31);
output(4, 31) <= input(33);
output(4, 32) <= input(17);
output(4, 33) <= input(18);
output(4, 34) <= input(19);
output(4, 35) <= input(20);
output(4, 36) <= input(21);
output(4, 37) <= input(22);
output(4, 38) <= input(23);
output(4, 39) <= input(24);
output(4, 40) <= input(25);
output(4, 41) <= input(26);
output(4, 42) <= input(27);
output(4, 43) <= input(28);
output(4, 44) <= input(29);
output(4, 45) <= input(30);
output(4, 46) <= input(31);
output(4, 47) <= input(33);
output(4, 48) <= input(17);
output(4, 49) <= input(18);
output(4, 50) <= input(19);
output(4, 51) <= input(20);
output(4, 52) <= input(21);
output(4, 53) <= input(22);
output(4, 54) <= input(23);
output(4, 55) <= input(24);
output(4, 56) <= input(25);
output(4, 57) <= input(26);
output(4, 58) <= input(27);
output(4, 59) <= input(28);
output(4, 60) <= input(29);
output(4, 61) <= input(30);
output(4, 62) <= input(31);
output(4, 63) <= input(33);
output(4, 64) <= input(17);
output(4, 65) <= input(18);
output(4, 66) <= input(19);
output(4, 67) <= input(20);
output(4, 68) <= input(21);
output(4, 69) <= input(22);
output(4, 70) <= input(23);
output(4, 71) <= input(24);
output(4, 72) <= input(25);
output(4, 73) <= input(26);
output(4, 74) <= input(27);
output(4, 75) <= input(28);
output(4, 76) <= input(29);
output(4, 77) <= input(30);
output(4, 78) <= input(31);
output(4, 79) <= input(33);
output(4, 80) <= input(17);
output(4, 81) <= input(18);
output(4, 82) <= input(19);
output(4, 83) <= input(20);
output(4, 84) <= input(21);
output(4, 85) <= input(22);
output(4, 86) <= input(23);
output(4, 87) <= input(24);
output(4, 88) <= input(25);
output(4, 89) <= input(26);
output(4, 90) <= input(27);
output(4, 91) <= input(28);
output(4, 92) <= input(29);
output(4, 93) <= input(30);
output(4, 94) <= input(31);
output(4, 95) <= input(33);
output(4, 96) <= input(17);
output(4, 97) <= input(18);
output(4, 98) <= input(19);
output(4, 99) <= input(20);
output(4, 100) <= input(21);
output(4, 101) <= input(22);
output(4, 102) <= input(23);
output(4, 103) <= input(24);
output(4, 104) <= input(25);
output(4, 105) <= input(26);
output(4, 106) <= input(27);
output(4, 107) <= input(28);
output(4, 108) <= input(29);
output(4, 109) <= input(30);
output(4, 110) <= input(31);
output(4, 111) <= input(33);
output(4, 112) <= input(17);
output(4, 113) <= input(18);
output(4, 114) <= input(19);
output(4, 115) <= input(20);
output(4, 116) <= input(21);
output(4, 117) <= input(22);
output(4, 118) <= input(23);
output(4, 119) <= input(24);
output(4, 120) <= input(25);
output(4, 121) <= input(26);
output(4, 122) <= input(27);
output(4, 123) <= input(28);
output(4, 124) <= input(29);
output(4, 125) <= input(30);
output(4, 126) <= input(31);
output(4, 127) <= input(33);
output(4, 128) <= input(17);
output(4, 129) <= input(18);
output(4, 130) <= input(19);
output(4, 131) <= input(20);
output(4, 132) <= input(21);
output(4, 133) <= input(22);
output(4, 134) <= input(23);
output(4, 135) <= input(24);
output(4, 136) <= input(25);
output(4, 137) <= input(26);
output(4, 138) <= input(27);
output(4, 139) <= input(28);
output(4, 140) <= input(29);
output(4, 141) <= input(30);
output(4, 142) <= input(31);
output(4, 143) <= input(33);
output(4, 144) <= input(17);
output(4, 145) <= input(18);
output(4, 146) <= input(19);
output(4, 147) <= input(20);
output(4, 148) <= input(21);
output(4, 149) <= input(22);
output(4, 150) <= input(23);
output(4, 151) <= input(24);
output(4, 152) <= input(25);
output(4, 153) <= input(26);
output(4, 154) <= input(27);
output(4, 155) <= input(28);
output(4, 156) <= input(29);
output(4, 157) <= input(30);
output(4, 158) <= input(31);
output(4, 159) <= input(33);
output(4, 160) <= input(17);
output(4, 161) <= input(18);
output(4, 162) <= input(19);
output(4, 163) <= input(20);
output(4, 164) <= input(21);
output(4, 165) <= input(22);
output(4, 166) <= input(23);
output(4, 167) <= input(24);
output(4, 168) <= input(25);
output(4, 169) <= input(26);
output(4, 170) <= input(27);
output(4, 171) <= input(28);
output(4, 172) <= input(29);
output(4, 173) <= input(30);
output(4, 174) <= input(31);
output(4, 175) <= input(33);
output(4, 176) <= input(17);
output(4, 177) <= input(18);
output(4, 178) <= input(19);
output(4, 179) <= input(20);
output(4, 180) <= input(21);
output(4, 181) <= input(22);
output(4, 182) <= input(23);
output(4, 183) <= input(24);
output(4, 184) <= input(25);
output(4, 185) <= input(26);
output(4, 186) <= input(27);
output(4, 187) <= input(28);
output(4, 188) <= input(29);
output(4, 189) <= input(30);
output(4, 190) <= input(31);
output(4, 191) <= input(33);
output(4, 192) <= input(17);
output(4, 193) <= input(18);
output(4, 194) <= input(19);
output(4, 195) <= input(20);
output(4, 196) <= input(21);
output(4, 197) <= input(22);
output(4, 198) <= input(23);
output(4, 199) <= input(24);
output(4, 200) <= input(25);
output(4, 201) <= input(26);
output(4, 202) <= input(27);
output(4, 203) <= input(28);
output(4, 204) <= input(29);
output(4, 205) <= input(30);
output(4, 206) <= input(31);
output(4, 207) <= input(33);
output(4, 208) <= input(17);
output(4, 209) <= input(18);
output(4, 210) <= input(19);
output(4, 211) <= input(20);
output(4, 212) <= input(21);
output(4, 213) <= input(22);
output(4, 214) <= input(23);
output(4, 215) <= input(24);
output(4, 216) <= input(25);
output(4, 217) <= input(26);
output(4, 218) <= input(27);
output(4, 219) <= input(28);
output(4, 220) <= input(29);
output(4, 221) <= input(30);
output(4, 222) <= input(31);
output(4, 223) <= input(33);
output(4, 224) <= input(17);
output(4, 225) <= input(18);
output(4, 226) <= input(19);
output(4, 227) <= input(20);
output(4, 228) <= input(21);
output(4, 229) <= input(22);
output(4, 230) <= input(23);
output(4, 231) <= input(24);
output(4, 232) <= input(25);
output(4, 233) <= input(26);
output(4, 234) <= input(27);
output(4, 235) <= input(28);
output(4, 236) <= input(29);
output(4, 237) <= input(30);
output(4, 238) <= input(31);
output(4, 239) <= input(33);
output(4, 240) <= input(1);
output(4, 241) <= input(2);
output(4, 242) <= input(3);
output(4, 243) <= input(4);
output(4, 244) <= input(5);
output(4, 245) <= input(6);
output(4, 246) <= input(7);
output(4, 247) <= input(8);
output(4, 248) <= input(9);
output(4, 249) <= input(10);
output(4, 250) <= input(11);
output(4, 251) <= input(12);
output(4, 252) <= input(13);
output(4, 253) <= input(14);
output(4, 254) <= input(15);
output(4, 255) <= input(34);
output(5, 0) <= input(17);
output(5, 1) <= input(18);
output(5, 2) <= input(19);
output(5, 3) <= input(20);
output(5, 4) <= input(21);
output(5, 5) <= input(22);
output(5, 6) <= input(23);
output(5, 7) <= input(24);
output(5, 8) <= input(25);
output(5, 9) <= input(26);
output(5, 10) <= input(27);
output(5, 11) <= input(28);
output(5, 12) <= input(29);
output(5, 13) <= input(30);
output(5, 14) <= input(31);
output(5, 15) <= input(33);
output(5, 16) <= input(17);
output(5, 17) <= input(18);
output(5, 18) <= input(19);
output(5, 19) <= input(20);
output(5, 20) <= input(21);
output(5, 21) <= input(22);
output(5, 22) <= input(23);
output(5, 23) <= input(24);
output(5, 24) <= input(25);
output(5, 25) <= input(26);
output(5, 26) <= input(27);
output(5, 27) <= input(28);
output(5, 28) <= input(29);
output(5, 29) <= input(30);
output(5, 30) <= input(31);
output(5, 31) <= input(33);
output(5, 32) <= input(17);
output(5, 33) <= input(18);
output(5, 34) <= input(19);
output(5, 35) <= input(20);
output(5, 36) <= input(21);
output(5, 37) <= input(22);
output(5, 38) <= input(23);
output(5, 39) <= input(24);
output(5, 40) <= input(25);
output(5, 41) <= input(26);
output(5, 42) <= input(27);
output(5, 43) <= input(28);
output(5, 44) <= input(29);
output(5, 45) <= input(30);
output(5, 46) <= input(31);
output(5, 47) <= input(33);
output(5, 48) <= input(17);
output(5, 49) <= input(18);
output(5, 50) <= input(19);
output(5, 51) <= input(20);
output(5, 52) <= input(21);
output(5, 53) <= input(22);
output(5, 54) <= input(23);
output(5, 55) <= input(24);
output(5, 56) <= input(25);
output(5, 57) <= input(26);
output(5, 58) <= input(27);
output(5, 59) <= input(28);
output(5, 60) <= input(29);
output(5, 61) <= input(30);
output(5, 62) <= input(31);
output(5, 63) <= input(33);
output(5, 64) <= input(17);
output(5, 65) <= input(18);
output(5, 66) <= input(19);
output(5, 67) <= input(20);
output(5, 68) <= input(21);
output(5, 69) <= input(22);
output(5, 70) <= input(23);
output(5, 71) <= input(24);
output(5, 72) <= input(25);
output(5, 73) <= input(26);
output(5, 74) <= input(27);
output(5, 75) <= input(28);
output(5, 76) <= input(29);
output(5, 77) <= input(30);
output(5, 78) <= input(31);
output(5, 79) <= input(33);
output(5, 80) <= input(17);
output(5, 81) <= input(18);
output(5, 82) <= input(19);
output(5, 83) <= input(20);
output(5, 84) <= input(21);
output(5, 85) <= input(22);
output(5, 86) <= input(23);
output(5, 87) <= input(24);
output(5, 88) <= input(25);
output(5, 89) <= input(26);
output(5, 90) <= input(27);
output(5, 91) <= input(28);
output(5, 92) <= input(29);
output(5, 93) <= input(30);
output(5, 94) <= input(31);
output(5, 95) <= input(33);
output(5, 96) <= input(17);
output(5, 97) <= input(18);
output(5, 98) <= input(19);
output(5, 99) <= input(20);
output(5, 100) <= input(21);
output(5, 101) <= input(22);
output(5, 102) <= input(23);
output(5, 103) <= input(24);
output(5, 104) <= input(25);
output(5, 105) <= input(26);
output(5, 106) <= input(27);
output(5, 107) <= input(28);
output(5, 108) <= input(29);
output(5, 109) <= input(30);
output(5, 110) <= input(31);
output(5, 111) <= input(33);
output(5, 112) <= input(1);
output(5, 113) <= input(2);
output(5, 114) <= input(3);
output(5, 115) <= input(4);
output(5, 116) <= input(5);
output(5, 117) <= input(6);
output(5, 118) <= input(7);
output(5, 119) <= input(8);
output(5, 120) <= input(9);
output(5, 121) <= input(10);
output(5, 122) <= input(11);
output(5, 123) <= input(12);
output(5, 124) <= input(13);
output(5, 125) <= input(14);
output(5, 126) <= input(15);
output(5, 127) <= input(34);
output(5, 128) <= input(1);
output(5, 129) <= input(2);
output(5, 130) <= input(3);
output(5, 131) <= input(4);
output(5, 132) <= input(5);
output(5, 133) <= input(6);
output(5, 134) <= input(7);
output(5, 135) <= input(8);
output(5, 136) <= input(9);
output(5, 137) <= input(10);
output(5, 138) <= input(11);
output(5, 139) <= input(12);
output(5, 140) <= input(13);
output(5, 141) <= input(14);
output(5, 142) <= input(15);
output(5, 143) <= input(34);
output(5, 144) <= input(1);
output(5, 145) <= input(2);
output(5, 146) <= input(3);
output(5, 147) <= input(4);
output(5, 148) <= input(5);
output(5, 149) <= input(6);
output(5, 150) <= input(7);
output(5, 151) <= input(8);
output(5, 152) <= input(9);
output(5, 153) <= input(10);
output(5, 154) <= input(11);
output(5, 155) <= input(12);
output(5, 156) <= input(13);
output(5, 157) <= input(14);
output(5, 158) <= input(15);
output(5, 159) <= input(34);
output(5, 160) <= input(1);
output(5, 161) <= input(2);
output(5, 162) <= input(3);
output(5, 163) <= input(4);
output(5, 164) <= input(5);
output(5, 165) <= input(6);
output(5, 166) <= input(7);
output(5, 167) <= input(8);
output(5, 168) <= input(9);
output(5, 169) <= input(10);
output(5, 170) <= input(11);
output(5, 171) <= input(12);
output(5, 172) <= input(13);
output(5, 173) <= input(14);
output(5, 174) <= input(15);
output(5, 175) <= input(34);
output(5, 176) <= input(1);
output(5, 177) <= input(2);
output(5, 178) <= input(3);
output(5, 179) <= input(4);
output(5, 180) <= input(5);
output(5, 181) <= input(6);
output(5, 182) <= input(7);
output(5, 183) <= input(8);
output(5, 184) <= input(9);
output(5, 185) <= input(10);
output(5, 186) <= input(11);
output(5, 187) <= input(12);
output(5, 188) <= input(13);
output(5, 189) <= input(14);
output(5, 190) <= input(15);
output(5, 191) <= input(34);
output(5, 192) <= input(1);
output(5, 193) <= input(2);
output(5, 194) <= input(3);
output(5, 195) <= input(4);
output(5, 196) <= input(5);
output(5, 197) <= input(6);
output(5, 198) <= input(7);
output(5, 199) <= input(8);
output(5, 200) <= input(9);
output(5, 201) <= input(10);
output(5, 202) <= input(11);
output(5, 203) <= input(12);
output(5, 204) <= input(13);
output(5, 205) <= input(14);
output(5, 206) <= input(15);
output(5, 207) <= input(34);
output(5, 208) <= input(1);
output(5, 209) <= input(2);
output(5, 210) <= input(3);
output(5, 211) <= input(4);
output(5, 212) <= input(5);
output(5, 213) <= input(6);
output(5, 214) <= input(7);
output(5, 215) <= input(8);
output(5, 216) <= input(9);
output(5, 217) <= input(10);
output(5, 218) <= input(11);
output(5, 219) <= input(12);
output(5, 220) <= input(13);
output(5, 221) <= input(14);
output(5, 222) <= input(15);
output(5, 223) <= input(34);
output(5, 224) <= input(1);
output(5, 225) <= input(2);
output(5, 226) <= input(3);
output(5, 227) <= input(4);
output(5, 228) <= input(5);
output(5, 229) <= input(6);
output(5, 230) <= input(7);
output(5, 231) <= input(8);
output(5, 232) <= input(9);
output(5, 233) <= input(10);
output(5, 234) <= input(11);
output(5, 235) <= input(12);
output(5, 236) <= input(13);
output(5, 237) <= input(14);
output(5, 238) <= input(15);
output(5, 239) <= input(34);
output(5, 240) <= input(18);
output(5, 241) <= input(19);
output(5, 242) <= input(20);
output(5, 243) <= input(21);
output(5, 244) <= input(22);
output(5, 245) <= input(23);
output(5, 246) <= input(24);
output(5, 247) <= input(25);
output(5, 248) <= input(26);
output(5, 249) <= input(27);
output(5, 250) <= input(28);
output(5, 251) <= input(29);
output(5, 252) <= input(30);
output(5, 253) <= input(31);
output(5, 254) <= input(33);
output(5, 255) <= input(35);
output(6, 0) <= input(17);
output(6, 1) <= input(18);
output(6, 2) <= input(19);
output(6, 3) <= input(20);
output(6, 4) <= input(21);
output(6, 5) <= input(22);
output(6, 6) <= input(23);
output(6, 7) <= input(24);
output(6, 8) <= input(25);
output(6, 9) <= input(26);
output(6, 10) <= input(27);
output(6, 11) <= input(28);
output(6, 12) <= input(29);
output(6, 13) <= input(30);
output(6, 14) <= input(31);
output(6, 15) <= input(33);
output(6, 16) <= input(17);
output(6, 17) <= input(18);
output(6, 18) <= input(19);
output(6, 19) <= input(20);
output(6, 20) <= input(21);
output(6, 21) <= input(22);
output(6, 22) <= input(23);
output(6, 23) <= input(24);
output(6, 24) <= input(25);
output(6, 25) <= input(26);
output(6, 26) <= input(27);
output(6, 27) <= input(28);
output(6, 28) <= input(29);
output(6, 29) <= input(30);
output(6, 30) <= input(31);
output(6, 31) <= input(33);
output(6, 32) <= input(17);
output(6, 33) <= input(18);
output(6, 34) <= input(19);
output(6, 35) <= input(20);
output(6, 36) <= input(21);
output(6, 37) <= input(22);
output(6, 38) <= input(23);
output(6, 39) <= input(24);
output(6, 40) <= input(25);
output(6, 41) <= input(26);
output(6, 42) <= input(27);
output(6, 43) <= input(28);
output(6, 44) <= input(29);
output(6, 45) <= input(30);
output(6, 46) <= input(31);
output(6, 47) <= input(33);
output(6, 48) <= input(17);
output(6, 49) <= input(18);
output(6, 50) <= input(19);
output(6, 51) <= input(20);
output(6, 52) <= input(21);
output(6, 53) <= input(22);
output(6, 54) <= input(23);
output(6, 55) <= input(24);
output(6, 56) <= input(25);
output(6, 57) <= input(26);
output(6, 58) <= input(27);
output(6, 59) <= input(28);
output(6, 60) <= input(29);
output(6, 61) <= input(30);
output(6, 62) <= input(31);
output(6, 63) <= input(33);
output(6, 64) <= input(17);
output(6, 65) <= input(18);
output(6, 66) <= input(19);
output(6, 67) <= input(20);
output(6, 68) <= input(21);
output(6, 69) <= input(22);
output(6, 70) <= input(23);
output(6, 71) <= input(24);
output(6, 72) <= input(25);
output(6, 73) <= input(26);
output(6, 74) <= input(27);
output(6, 75) <= input(28);
output(6, 76) <= input(29);
output(6, 77) <= input(30);
output(6, 78) <= input(31);
output(6, 79) <= input(33);
output(6, 80) <= input(1);
output(6, 81) <= input(2);
output(6, 82) <= input(3);
output(6, 83) <= input(4);
output(6, 84) <= input(5);
output(6, 85) <= input(6);
output(6, 86) <= input(7);
output(6, 87) <= input(8);
output(6, 88) <= input(9);
output(6, 89) <= input(10);
output(6, 90) <= input(11);
output(6, 91) <= input(12);
output(6, 92) <= input(13);
output(6, 93) <= input(14);
output(6, 94) <= input(15);
output(6, 95) <= input(34);
output(6, 96) <= input(1);
output(6, 97) <= input(2);
output(6, 98) <= input(3);
output(6, 99) <= input(4);
output(6, 100) <= input(5);
output(6, 101) <= input(6);
output(6, 102) <= input(7);
output(6, 103) <= input(8);
output(6, 104) <= input(9);
output(6, 105) <= input(10);
output(6, 106) <= input(11);
output(6, 107) <= input(12);
output(6, 108) <= input(13);
output(6, 109) <= input(14);
output(6, 110) <= input(15);
output(6, 111) <= input(34);
output(6, 112) <= input(1);
output(6, 113) <= input(2);
output(6, 114) <= input(3);
output(6, 115) <= input(4);
output(6, 116) <= input(5);
output(6, 117) <= input(6);
output(6, 118) <= input(7);
output(6, 119) <= input(8);
output(6, 120) <= input(9);
output(6, 121) <= input(10);
output(6, 122) <= input(11);
output(6, 123) <= input(12);
output(6, 124) <= input(13);
output(6, 125) <= input(14);
output(6, 126) <= input(15);
output(6, 127) <= input(34);
output(6, 128) <= input(1);
output(6, 129) <= input(2);
output(6, 130) <= input(3);
output(6, 131) <= input(4);
output(6, 132) <= input(5);
output(6, 133) <= input(6);
output(6, 134) <= input(7);
output(6, 135) <= input(8);
output(6, 136) <= input(9);
output(6, 137) <= input(10);
output(6, 138) <= input(11);
output(6, 139) <= input(12);
output(6, 140) <= input(13);
output(6, 141) <= input(14);
output(6, 142) <= input(15);
output(6, 143) <= input(34);
output(6, 144) <= input(1);
output(6, 145) <= input(2);
output(6, 146) <= input(3);
output(6, 147) <= input(4);
output(6, 148) <= input(5);
output(6, 149) <= input(6);
output(6, 150) <= input(7);
output(6, 151) <= input(8);
output(6, 152) <= input(9);
output(6, 153) <= input(10);
output(6, 154) <= input(11);
output(6, 155) <= input(12);
output(6, 156) <= input(13);
output(6, 157) <= input(14);
output(6, 158) <= input(15);
output(6, 159) <= input(34);
output(6, 160) <= input(18);
output(6, 161) <= input(19);
output(6, 162) <= input(20);
output(6, 163) <= input(21);
output(6, 164) <= input(22);
output(6, 165) <= input(23);
output(6, 166) <= input(24);
output(6, 167) <= input(25);
output(6, 168) <= input(26);
output(6, 169) <= input(27);
output(6, 170) <= input(28);
output(6, 171) <= input(29);
output(6, 172) <= input(30);
output(6, 173) <= input(31);
output(6, 174) <= input(33);
output(6, 175) <= input(35);
output(6, 176) <= input(18);
output(6, 177) <= input(19);
output(6, 178) <= input(20);
output(6, 179) <= input(21);
output(6, 180) <= input(22);
output(6, 181) <= input(23);
output(6, 182) <= input(24);
output(6, 183) <= input(25);
output(6, 184) <= input(26);
output(6, 185) <= input(27);
output(6, 186) <= input(28);
output(6, 187) <= input(29);
output(6, 188) <= input(30);
output(6, 189) <= input(31);
output(6, 190) <= input(33);
output(6, 191) <= input(35);
output(6, 192) <= input(18);
output(6, 193) <= input(19);
output(6, 194) <= input(20);
output(6, 195) <= input(21);
output(6, 196) <= input(22);
output(6, 197) <= input(23);
output(6, 198) <= input(24);
output(6, 199) <= input(25);
output(6, 200) <= input(26);
output(6, 201) <= input(27);
output(6, 202) <= input(28);
output(6, 203) <= input(29);
output(6, 204) <= input(30);
output(6, 205) <= input(31);
output(6, 206) <= input(33);
output(6, 207) <= input(35);
output(6, 208) <= input(18);
output(6, 209) <= input(19);
output(6, 210) <= input(20);
output(6, 211) <= input(21);
output(6, 212) <= input(22);
output(6, 213) <= input(23);
output(6, 214) <= input(24);
output(6, 215) <= input(25);
output(6, 216) <= input(26);
output(6, 217) <= input(27);
output(6, 218) <= input(28);
output(6, 219) <= input(29);
output(6, 220) <= input(30);
output(6, 221) <= input(31);
output(6, 222) <= input(33);
output(6, 223) <= input(35);
output(6, 224) <= input(18);
output(6, 225) <= input(19);
output(6, 226) <= input(20);
output(6, 227) <= input(21);
output(6, 228) <= input(22);
output(6, 229) <= input(23);
output(6, 230) <= input(24);
output(6, 231) <= input(25);
output(6, 232) <= input(26);
output(6, 233) <= input(27);
output(6, 234) <= input(28);
output(6, 235) <= input(29);
output(6, 236) <= input(30);
output(6, 237) <= input(31);
output(6, 238) <= input(33);
output(6, 239) <= input(35);
output(6, 240) <= input(2);
output(6, 241) <= input(3);
output(6, 242) <= input(4);
output(6, 243) <= input(5);
output(6, 244) <= input(6);
output(6, 245) <= input(7);
output(6, 246) <= input(8);
output(6, 247) <= input(9);
output(6, 248) <= input(10);
output(6, 249) <= input(11);
output(6, 250) <= input(12);
output(6, 251) <= input(13);
output(6, 252) <= input(14);
output(6, 253) <= input(15);
output(6, 254) <= input(34);
output(6, 255) <= input(36);
output(7, 0) <= input(17);
output(7, 1) <= input(18);
output(7, 2) <= input(19);
output(7, 3) <= input(20);
output(7, 4) <= input(21);
output(7, 5) <= input(22);
output(7, 6) <= input(23);
output(7, 7) <= input(24);
output(7, 8) <= input(25);
output(7, 9) <= input(26);
output(7, 10) <= input(27);
output(7, 11) <= input(28);
output(7, 12) <= input(29);
output(7, 13) <= input(30);
output(7, 14) <= input(31);
output(7, 15) <= input(33);
output(7, 16) <= input(17);
output(7, 17) <= input(18);
output(7, 18) <= input(19);
output(7, 19) <= input(20);
output(7, 20) <= input(21);
output(7, 21) <= input(22);
output(7, 22) <= input(23);
output(7, 23) <= input(24);
output(7, 24) <= input(25);
output(7, 25) <= input(26);
output(7, 26) <= input(27);
output(7, 27) <= input(28);
output(7, 28) <= input(29);
output(7, 29) <= input(30);
output(7, 30) <= input(31);
output(7, 31) <= input(33);
output(7, 32) <= input(17);
output(7, 33) <= input(18);
output(7, 34) <= input(19);
output(7, 35) <= input(20);
output(7, 36) <= input(21);
output(7, 37) <= input(22);
output(7, 38) <= input(23);
output(7, 39) <= input(24);
output(7, 40) <= input(25);
output(7, 41) <= input(26);
output(7, 42) <= input(27);
output(7, 43) <= input(28);
output(7, 44) <= input(29);
output(7, 45) <= input(30);
output(7, 46) <= input(31);
output(7, 47) <= input(33);
output(7, 48) <= input(1);
output(7, 49) <= input(2);
output(7, 50) <= input(3);
output(7, 51) <= input(4);
output(7, 52) <= input(5);
output(7, 53) <= input(6);
output(7, 54) <= input(7);
output(7, 55) <= input(8);
output(7, 56) <= input(9);
output(7, 57) <= input(10);
output(7, 58) <= input(11);
output(7, 59) <= input(12);
output(7, 60) <= input(13);
output(7, 61) <= input(14);
output(7, 62) <= input(15);
output(7, 63) <= input(34);
output(7, 64) <= input(1);
output(7, 65) <= input(2);
output(7, 66) <= input(3);
output(7, 67) <= input(4);
output(7, 68) <= input(5);
output(7, 69) <= input(6);
output(7, 70) <= input(7);
output(7, 71) <= input(8);
output(7, 72) <= input(9);
output(7, 73) <= input(10);
output(7, 74) <= input(11);
output(7, 75) <= input(12);
output(7, 76) <= input(13);
output(7, 77) <= input(14);
output(7, 78) <= input(15);
output(7, 79) <= input(34);
output(7, 80) <= input(1);
output(7, 81) <= input(2);
output(7, 82) <= input(3);
output(7, 83) <= input(4);
output(7, 84) <= input(5);
output(7, 85) <= input(6);
output(7, 86) <= input(7);
output(7, 87) <= input(8);
output(7, 88) <= input(9);
output(7, 89) <= input(10);
output(7, 90) <= input(11);
output(7, 91) <= input(12);
output(7, 92) <= input(13);
output(7, 93) <= input(14);
output(7, 94) <= input(15);
output(7, 95) <= input(34);
output(7, 96) <= input(1);
output(7, 97) <= input(2);
output(7, 98) <= input(3);
output(7, 99) <= input(4);
output(7, 100) <= input(5);
output(7, 101) <= input(6);
output(7, 102) <= input(7);
output(7, 103) <= input(8);
output(7, 104) <= input(9);
output(7, 105) <= input(10);
output(7, 106) <= input(11);
output(7, 107) <= input(12);
output(7, 108) <= input(13);
output(7, 109) <= input(14);
output(7, 110) <= input(15);
output(7, 111) <= input(34);
output(7, 112) <= input(18);
output(7, 113) <= input(19);
output(7, 114) <= input(20);
output(7, 115) <= input(21);
output(7, 116) <= input(22);
output(7, 117) <= input(23);
output(7, 118) <= input(24);
output(7, 119) <= input(25);
output(7, 120) <= input(26);
output(7, 121) <= input(27);
output(7, 122) <= input(28);
output(7, 123) <= input(29);
output(7, 124) <= input(30);
output(7, 125) <= input(31);
output(7, 126) <= input(33);
output(7, 127) <= input(35);
output(7, 128) <= input(18);
output(7, 129) <= input(19);
output(7, 130) <= input(20);
output(7, 131) <= input(21);
output(7, 132) <= input(22);
output(7, 133) <= input(23);
output(7, 134) <= input(24);
output(7, 135) <= input(25);
output(7, 136) <= input(26);
output(7, 137) <= input(27);
output(7, 138) <= input(28);
output(7, 139) <= input(29);
output(7, 140) <= input(30);
output(7, 141) <= input(31);
output(7, 142) <= input(33);
output(7, 143) <= input(35);
output(7, 144) <= input(18);
output(7, 145) <= input(19);
output(7, 146) <= input(20);
output(7, 147) <= input(21);
output(7, 148) <= input(22);
output(7, 149) <= input(23);
output(7, 150) <= input(24);
output(7, 151) <= input(25);
output(7, 152) <= input(26);
output(7, 153) <= input(27);
output(7, 154) <= input(28);
output(7, 155) <= input(29);
output(7, 156) <= input(30);
output(7, 157) <= input(31);
output(7, 158) <= input(33);
output(7, 159) <= input(35);
output(7, 160) <= input(18);
output(7, 161) <= input(19);
output(7, 162) <= input(20);
output(7, 163) <= input(21);
output(7, 164) <= input(22);
output(7, 165) <= input(23);
output(7, 166) <= input(24);
output(7, 167) <= input(25);
output(7, 168) <= input(26);
output(7, 169) <= input(27);
output(7, 170) <= input(28);
output(7, 171) <= input(29);
output(7, 172) <= input(30);
output(7, 173) <= input(31);
output(7, 174) <= input(33);
output(7, 175) <= input(35);
output(7, 176) <= input(2);
output(7, 177) <= input(3);
output(7, 178) <= input(4);
output(7, 179) <= input(5);
output(7, 180) <= input(6);
output(7, 181) <= input(7);
output(7, 182) <= input(8);
output(7, 183) <= input(9);
output(7, 184) <= input(10);
output(7, 185) <= input(11);
output(7, 186) <= input(12);
output(7, 187) <= input(13);
output(7, 188) <= input(14);
output(7, 189) <= input(15);
output(7, 190) <= input(34);
output(7, 191) <= input(36);
output(7, 192) <= input(2);
output(7, 193) <= input(3);
output(7, 194) <= input(4);
output(7, 195) <= input(5);
output(7, 196) <= input(6);
output(7, 197) <= input(7);
output(7, 198) <= input(8);
output(7, 199) <= input(9);
output(7, 200) <= input(10);
output(7, 201) <= input(11);
output(7, 202) <= input(12);
output(7, 203) <= input(13);
output(7, 204) <= input(14);
output(7, 205) <= input(15);
output(7, 206) <= input(34);
output(7, 207) <= input(36);
output(7, 208) <= input(2);
output(7, 209) <= input(3);
output(7, 210) <= input(4);
output(7, 211) <= input(5);
output(7, 212) <= input(6);
output(7, 213) <= input(7);
output(7, 214) <= input(8);
output(7, 215) <= input(9);
output(7, 216) <= input(10);
output(7, 217) <= input(11);
output(7, 218) <= input(12);
output(7, 219) <= input(13);
output(7, 220) <= input(14);
output(7, 221) <= input(15);
output(7, 222) <= input(34);
output(7, 223) <= input(36);
output(7, 224) <= input(2);
output(7, 225) <= input(3);
output(7, 226) <= input(4);
output(7, 227) <= input(5);
output(7, 228) <= input(6);
output(7, 229) <= input(7);
output(7, 230) <= input(8);
output(7, 231) <= input(9);
output(7, 232) <= input(10);
output(7, 233) <= input(11);
output(7, 234) <= input(12);
output(7, 235) <= input(13);
output(7, 236) <= input(14);
output(7, 237) <= input(15);
output(7, 238) <= input(34);
output(7, 239) <= input(36);
output(7, 240) <= input(19);
output(7, 241) <= input(20);
output(7, 242) <= input(21);
output(7, 243) <= input(22);
output(7, 244) <= input(23);
output(7, 245) <= input(24);
output(7, 246) <= input(25);
output(7, 247) <= input(26);
output(7, 248) <= input(27);
output(7, 249) <= input(28);
output(7, 250) <= input(29);
output(7, 251) <= input(30);
output(7, 252) <= input(31);
output(7, 253) <= input(33);
output(7, 254) <= input(35);
output(7, 255) <= input(37);
when "1110" =>
output(0, 0) <= input(0);
output(0, 1) <= input(1);
output(0, 2) <= input(2);
output(0, 3) <= input(3);
output(0, 4) <= input(4);
output(0, 5) <= input(5);
output(0, 6) <= input(6);
output(0, 7) <= input(7);
output(0, 8) <= input(8);
output(0, 9) <= input(9);
output(0, 10) <= input(10);
output(0, 11) <= input(11);
output(0, 12) <= input(12);
output(0, 13) <= input(13);
output(0, 14) <= input(14);
output(0, 15) <= input(15);
output(0, 16) <= input(0);
output(0, 17) <= input(1);
output(0, 18) <= input(2);
output(0, 19) <= input(3);
output(0, 20) <= input(4);
output(0, 21) <= input(5);
output(0, 22) <= input(6);
output(0, 23) <= input(7);
output(0, 24) <= input(8);
output(0, 25) <= input(9);
output(0, 26) <= input(10);
output(0, 27) <= input(11);
output(0, 28) <= input(12);
output(0, 29) <= input(13);
output(0, 30) <= input(14);
output(0, 31) <= input(15);
output(0, 32) <= input(16);
output(0, 33) <= input(17);
output(0, 34) <= input(18);
output(0, 35) <= input(19);
output(0, 36) <= input(20);
output(0, 37) <= input(21);
output(0, 38) <= input(22);
output(0, 39) <= input(23);
output(0, 40) <= input(24);
output(0, 41) <= input(25);
output(0, 42) <= input(26);
output(0, 43) <= input(27);
output(0, 44) <= input(28);
output(0, 45) <= input(29);
output(0, 46) <= input(30);
output(0, 47) <= input(31);
output(0, 48) <= input(16);
output(0, 49) <= input(17);
output(0, 50) <= input(18);
output(0, 51) <= input(19);
output(0, 52) <= input(20);
output(0, 53) <= input(21);
output(0, 54) <= input(22);
output(0, 55) <= input(23);
output(0, 56) <= input(24);
output(0, 57) <= input(25);
output(0, 58) <= input(26);
output(0, 59) <= input(27);
output(0, 60) <= input(28);
output(0, 61) <= input(29);
output(0, 62) <= input(30);
output(0, 63) <= input(31);
output(0, 64) <= input(16);
output(0, 65) <= input(17);
output(0, 66) <= input(18);
output(0, 67) <= input(19);
output(0, 68) <= input(20);
output(0, 69) <= input(21);
output(0, 70) <= input(22);
output(0, 71) <= input(23);
output(0, 72) <= input(24);
output(0, 73) <= input(25);
output(0, 74) <= input(26);
output(0, 75) <= input(27);
output(0, 76) <= input(28);
output(0, 77) <= input(29);
output(0, 78) <= input(30);
output(0, 79) <= input(31);
output(0, 80) <= input(1);
output(0, 81) <= input(2);
output(0, 82) <= input(3);
output(0, 83) <= input(4);
output(0, 84) <= input(5);
output(0, 85) <= input(6);
output(0, 86) <= input(7);
output(0, 87) <= input(8);
output(0, 88) <= input(9);
output(0, 89) <= input(10);
output(0, 90) <= input(11);
output(0, 91) <= input(12);
output(0, 92) <= input(13);
output(0, 93) <= input(14);
output(0, 94) <= input(15);
output(0, 95) <= input(32);
output(0, 96) <= input(1);
output(0, 97) <= input(2);
output(0, 98) <= input(3);
output(0, 99) <= input(4);
output(0, 100) <= input(5);
output(0, 101) <= input(6);
output(0, 102) <= input(7);
output(0, 103) <= input(8);
output(0, 104) <= input(9);
output(0, 105) <= input(10);
output(0, 106) <= input(11);
output(0, 107) <= input(12);
output(0, 108) <= input(13);
output(0, 109) <= input(14);
output(0, 110) <= input(15);
output(0, 111) <= input(32);
output(0, 112) <= input(17);
output(0, 113) <= input(18);
output(0, 114) <= input(19);
output(0, 115) <= input(20);
output(0, 116) <= input(21);
output(0, 117) <= input(22);
output(0, 118) <= input(23);
output(0, 119) <= input(24);
output(0, 120) <= input(25);
output(0, 121) <= input(26);
output(0, 122) <= input(27);
output(0, 123) <= input(28);
output(0, 124) <= input(29);
output(0, 125) <= input(30);
output(0, 126) <= input(31);
output(0, 127) <= input(33);
output(0, 128) <= input(17);
output(0, 129) <= input(18);
output(0, 130) <= input(19);
output(0, 131) <= input(20);
output(0, 132) <= input(21);
output(0, 133) <= input(22);
output(0, 134) <= input(23);
output(0, 135) <= input(24);
output(0, 136) <= input(25);
output(0, 137) <= input(26);
output(0, 138) <= input(27);
output(0, 139) <= input(28);
output(0, 140) <= input(29);
output(0, 141) <= input(30);
output(0, 142) <= input(31);
output(0, 143) <= input(33);
output(0, 144) <= input(17);
output(0, 145) <= input(18);
output(0, 146) <= input(19);
output(0, 147) <= input(20);
output(0, 148) <= input(21);
output(0, 149) <= input(22);
output(0, 150) <= input(23);
output(0, 151) <= input(24);
output(0, 152) <= input(25);
output(0, 153) <= input(26);
output(0, 154) <= input(27);
output(0, 155) <= input(28);
output(0, 156) <= input(29);
output(0, 157) <= input(30);
output(0, 158) <= input(31);
output(0, 159) <= input(33);
output(0, 160) <= input(2);
output(0, 161) <= input(3);
output(0, 162) <= input(4);
output(0, 163) <= input(5);
output(0, 164) <= input(6);
output(0, 165) <= input(7);
output(0, 166) <= input(8);
output(0, 167) <= input(9);
output(0, 168) <= input(10);
output(0, 169) <= input(11);
output(0, 170) <= input(12);
output(0, 171) <= input(13);
output(0, 172) <= input(14);
output(0, 173) <= input(15);
output(0, 174) <= input(32);
output(0, 175) <= input(34);
output(0, 176) <= input(2);
output(0, 177) <= input(3);
output(0, 178) <= input(4);
output(0, 179) <= input(5);
output(0, 180) <= input(6);
output(0, 181) <= input(7);
output(0, 182) <= input(8);
output(0, 183) <= input(9);
output(0, 184) <= input(10);
output(0, 185) <= input(11);
output(0, 186) <= input(12);
output(0, 187) <= input(13);
output(0, 188) <= input(14);
output(0, 189) <= input(15);
output(0, 190) <= input(32);
output(0, 191) <= input(34);
output(0, 192) <= input(2);
output(0, 193) <= input(3);
output(0, 194) <= input(4);
output(0, 195) <= input(5);
output(0, 196) <= input(6);
output(0, 197) <= input(7);
output(0, 198) <= input(8);
output(0, 199) <= input(9);
output(0, 200) <= input(10);
output(0, 201) <= input(11);
output(0, 202) <= input(12);
output(0, 203) <= input(13);
output(0, 204) <= input(14);
output(0, 205) <= input(15);
output(0, 206) <= input(32);
output(0, 207) <= input(34);
output(0, 208) <= input(18);
output(0, 209) <= input(19);
output(0, 210) <= input(20);
output(0, 211) <= input(21);
output(0, 212) <= input(22);
output(0, 213) <= input(23);
output(0, 214) <= input(24);
output(0, 215) <= input(25);
output(0, 216) <= input(26);
output(0, 217) <= input(27);
output(0, 218) <= input(28);
output(0, 219) <= input(29);
output(0, 220) <= input(30);
output(0, 221) <= input(31);
output(0, 222) <= input(33);
output(0, 223) <= input(35);
output(0, 224) <= input(18);
output(0, 225) <= input(19);
output(0, 226) <= input(20);
output(0, 227) <= input(21);
output(0, 228) <= input(22);
output(0, 229) <= input(23);
output(0, 230) <= input(24);
output(0, 231) <= input(25);
output(0, 232) <= input(26);
output(0, 233) <= input(27);
output(0, 234) <= input(28);
output(0, 235) <= input(29);
output(0, 236) <= input(30);
output(0, 237) <= input(31);
output(0, 238) <= input(33);
output(0, 239) <= input(35);
output(0, 240) <= input(3);
output(0, 241) <= input(4);
output(0, 242) <= input(5);
output(0, 243) <= input(6);
output(0, 244) <= input(7);
output(0, 245) <= input(8);
output(0, 246) <= input(9);
output(0, 247) <= input(10);
output(0, 248) <= input(11);
output(0, 249) <= input(12);
output(0, 250) <= input(13);
output(0, 251) <= input(14);
output(0, 252) <= input(15);
output(0, 253) <= input(32);
output(0, 254) <= input(34);
output(0, 255) <= input(36);
output(1, 0) <= input(0);
output(1, 1) <= input(1);
output(1, 2) <= input(2);
output(1, 3) <= input(3);
output(1, 4) <= input(4);
output(1, 5) <= input(5);
output(1, 6) <= input(6);
output(1, 7) <= input(7);
output(1, 8) <= input(8);
output(1, 9) <= input(9);
output(1, 10) <= input(10);
output(1, 11) <= input(11);
output(1, 12) <= input(12);
output(1, 13) <= input(13);
output(1, 14) <= input(14);
output(1, 15) <= input(15);
output(1, 16) <= input(16);
output(1, 17) <= input(17);
output(1, 18) <= input(18);
output(1, 19) <= input(19);
output(1, 20) <= input(20);
output(1, 21) <= input(21);
output(1, 22) <= input(22);
output(1, 23) <= input(23);
output(1, 24) <= input(24);
output(1, 25) <= input(25);
output(1, 26) <= input(26);
output(1, 27) <= input(27);
output(1, 28) <= input(28);
output(1, 29) <= input(29);
output(1, 30) <= input(30);
output(1, 31) <= input(31);
output(1, 32) <= input(16);
output(1, 33) <= input(17);
output(1, 34) <= input(18);
output(1, 35) <= input(19);
output(1, 36) <= input(20);
output(1, 37) <= input(21);
output(1, 38) <= input(22);
output(1, 39) <= input(23);
output(1, 40) <= input(24);
output(1, 41) <= input(25);
output(1, 42) <= input(26);
output(1, 43) <= input(27);
output(1, 44) <= input(28);
output(1, 45) <= input(29);
output(1, 46) <= input(30);
output(1, 47) <= input(31);
output(1, 48) <= input(1);
output(1, 49) <= input(2);
output(1, 50) <= input(3);
output(1, 51) <= input(4);
output(1, 52) <= input(5);
output(1, 53) <= input(6);
output(1, 54) <= input(7);
output(1, 55) <= input(8);
output(1, 56) <= input(9);
output(1, 57) <= input(10);
output(1, 58) <= input(11);
output(1, 59) <= input(12);
output(1, 60) <= input(13);
output(1, 61) <= input(14);
output(1, 62) <= input(15);
output(1, 63) <= input(32);
output(1, 64) <= input(1);
output(1, 65) <= input(2);
output(1, 66) <= input(3);
output(1, 67) <= input(4);
output(1, 68) <= input(5);
output(1, 69) <= input(6);
output(1, 70) <= input(7);
output(1, 71) <= input(8);
output(1, 72) <= input(9);
output(1, 73) <= input(10);
output(1, 74) <= input(11);
output(1, 75) <= input(12);
output(1, 76) <= input(13);
output(1, 77) <= input(14);
output(1, 78) <= input(15);
output(1, 79) <= input(32);
output(1, 80) <= input(17);
output(1, 81) <= input(18);
output(1, 82) <= input(19);
output(1, 83) <= input(20);
output(1, 84) <= input(21);
output(1, 85) <= input(22);
output(1, 86) <= input(23);
output(1, 87) <= input(24);
output(1, 88) <= input(25);
output(1, 89) <= input(26);
output(1, 90) <= input(27);
output(1, 91) <= input(28);
output(1, 92) <= input(29);
output(1, 93) <= input(30);
output(1, 94) <= input(31);
output(1, 95) <= input(33);
output(1, 96) <= input(17);
output(1, 97) <= input(18);
output(1, 98) <= input(19);
output(1, 99) <= input(20);
output(1, 100) <= input(21);
output(1, 101) <= input(22);
output(1, 102) <= input(23);
output(1, 103) <= input(24);
output(1, 104) <= input(25);
output(1, 105) <= input(26);
output(1, 106) <= input(27);
output(1, 107) <= input(28);
output(1, 108) <= input(29);
output(1, 109) <= input(30);
output(1, 110) <= input(31);
output(1, 111) <= input(33);
output(1, 112) <= input(2);
output(1, 113) <= input(3);
output(1, 114) <= input(4);
output(1, 115) <= input(5);
output(1, 116) <= input(6);
output(1, 117) <= input(7);
output(1, 118) <= input(8);
output(1, 119) <= input(9);
output(1, 120) <= input(10);
output(1, 121) <= input(11);
output(1, 122) <= input(12);
output(1, 123) <= input(13);
output(1, 124) <= input(14);
output(1, 125) <= input(15);
output(1, 126) <= input(32);
output(1, 127) <= input(34);
output(1, 128) <= input(2);
output(1, 129) <= input(3);
output(1, 130) <= input(4);
output(1, 131) <= input(5);
output(1, 132) <= input(6);
output(1, 133) <= input(7);
output(1, 134) <= input(8);
output(1, 135) <= input(9);
output(1, 136) <= input(10);
output(1, 137) <= input(11);
output(1, 138) <= input(12);
output(1, 139) <= input(13);
output(1, 140) <= input(14);
output(1, 141) <= input(15);
output(1, 142) <= input(32);
output(1, 143) <= input(34);
output(1, 144) <= input(18);
output(1, 145) <= input(19);
output(1, 146) <= input(20);
output(1, 147) <= input(21);
output(1, 148) <= input(22);
output(1, 149) <= input(23);
output(1, 150) <= input(24);
output(1, 151) <= input(25);
output(1, 152) <= input(26);
output(1, 153) <= input(27);
output(1, 154) <= input(28);
output(1, 155) <= input(29);
output(1, 156) <= input(30);
output(1, 157) <= input(31);
output(1, 158) <= input(33);
output(1, 159) <= input(35);
output(1, 160) <= input(18);
output(1, 161) <= input(19);
output(1, 162) <= input(20);
output(1, 163) <= input(21);
output(1, 164) <= input(22);
output(1, 165) <= input(23);
output(1, 166) <= input(24);
output(1, 167) <= input(25);
output(1, 168) <= input(26);
output(1, 169) <= input(27);
output(1, 170) <= input(28);
output(1, 171) <= input(29);
output(1, 172) <= input(30);
output(1, 173) <= input(31);
output(1, 174) <= input(33);
output(1, 175) <= input(35);
output(1, 176) <= input(3);
output(1, 177) <= input(4);
output(1, 178) <= input(5);
output(1, 179) <= input(6);
output(1, 180) <= input(7);
output(1, 181) <= input(8);
output(1, 182) <= input(9);
output(1, 183) <= input(10);
output(1, 184) <= input(11);
output(1, 185) <= input(12);
output(1, 186) <= input(13);
output(1, 187) <= input(14);
output(1, 188) <= input(15);
output(1, 189) <= input(32);
output(1, 190) <= input(34);
output(1, 191) <= input(36);
output(1, 192) <= input(3);
output(1, 193) <= input(4);
output(1, 194) <= input(5);
output(1, 195) <= input(6);
output(1, 196) <= input(7);
output(1, 197) <= input(8);
output(1, 198) <= input(9);
output(1, 199) <= input(10);
output(1, 200) <= input(11);
output(1, 201) <= input(12);
output(1, 202) <= input(13);
output(1, 203) <= input(14);
output(1, 204) <= input(15);
output(1, 205) <= input(32);
output(1, 206) <= input(34);
output(1, 207) <= input(36);
output(1, 208) <= input(19);
output(1, 209) <= input(20);
output(1, 210) <= input(21);
output(1, 211) <= input(22);
output(1, 212) <= input(23);
output(1, 213) <= input(24);
output(1, 214) <= input(25);
output(1, 215) <= input(26);
output(1, 216) <= input(27);
output(1, 217) <= input(28);
output(1, 218) <= input(29);
output(1, 219) <= input(30);
output(1, 220) <= input(31);
output(1, 221) <= input(33);
output(1, 222) <= input(35);
output(1, 223) <= input(37);
output(1, 224) <= input(19);
output(1, 225) <= input(20);
output(1, 226) <= input(21);
output(1, 227) <= input(22);
output(1, 228) <= input(23);
output(1, 229) <= input(24);
output(1, 230) <= input(25);
output(1, 231) <= input(26);
output(1, 232) <= input(27);
output(1, 233) <= input(28);
output(1, 234) <= input(29);
output(1, 235) <= input(30);
output(1, 236) <= input(31);
output(1, 237) <= input(33);
output(1, 238) <= input(35);
output(1, 239) <= input(37);
output(1, 240) <= input(4);
output(1, 241) <= input(5);
output(1, 242) <= input(6);
output(1, 243) <= input(7);
output(1, 244) <= input(8);
output(1, 245) <= input(9);
output(1, 246) <= input(10);
output(1, 247) <= input(11);
output(1, 248) <= input(12);
output(1, 249) <= input(13);
output(1, 250) <= input(14);
output(1, 251) <= input(15);
output(1, 252) <= input(32);
output(1, 253) <= input(34);
output(1, 254) <= input(36);
output(1, 255) <= input(38);
output(2, 0) <= input(0);
output(2, 1) <= input(1);
output(2, 2) <= input(2);
output(2, 3) <= input(3);
output(2, 4) <= input(4);
output(2, 5) <= input(5);
output(2, 6) <= input(6);
output(2, 7) <= input(7);
output(2, 8) <= input(8);
output(2, 9) <= input(9);
output(2, 10) <= input(10);
output(2, 11) <= input(11);
output(2, 12) <= input(12);
output(2, 13) <= input(13);
output(2, 14) <= input(14);
output(2, 15) <= input(15);
output(2, 16) <= input(16);
output(2, 17) <= input(17);
output(2, 18) <= input(18);
output(2, 19) <= input(19);
output(2, 20) <= input(20);
output(2, 21) <= input(21);
output(2, 22) <= input(22);
output(2, 23) <= input(23);
output(2, 24) <= input(24);
output(2, 25) <= input(25);
output(2, 26) <= input(26);
output(2, 27) <= input(27);
output(2, 28) <= input(28);
output(2, 29) <= input(29);
output(2, 30) <= input(30);
output(2, 31) <= input(31);
output(2, 32) <= input(16);
output(2, 33) <= input(17);
output(2, 34) <= input(18);
output(2, 35) <= input(19);
output(2, 36) <= input(20);
output(2, 37) <= input(21);
output(2, 38) <= input(22);
output(2, 39) <= input(23);
output(2, 40) <= input(24);
output(2, 41) <= input(25);
output(2, 42) <= input(26);
output(2, 43) <= input(27);
output(2, 44) <= input(28);
output(2, 45) <= input(29);
output(2, 46) <= input(30);
output(2, 47) <= input(31);
output(2, 48) <= input(1);
output(2, 49) <= input(2);
output(2, 50) <= input(3);
output(2, 51) <= input(4);
output(2, 52) <= input(5);
output(2, 53) <= input(6);
output(2, 54) <= input(7);
output(2, 55) <= input(8);
output(2, 56) <= input(9);
output(2, 57) <= input(10);
output(2, 58) <= input(11);
output(2, 59) <= input(12);
output(2, 60) <= input(13);
output(2, 61) <= input(14);
output(2, 62) <= input(15);
output(2, 63) <= input(32);
output(2, 64) <= input(17);
output(2, 65) <= input(18);
output(2, 66) <= input(19);
output(2, 67) <= input(20);
output(2, 68) <= input(21);
output(2, 69) <= input(22);
output(2, 70) <= input(23);
output(2, 71) <= input(24);
output(2, 72) <= input(25);
output(2, 73) <= input(26);
output(2, 74) <= input(27);
output(2, 75) <= input(28);
output(2, 76) <= input(29);
output(2, 77) <= input(30);
output(2, 78) <= input(31);
output(2, 79) <= input(33);
output(2, 80) <= input(17);
output(2, 81) <= input(18);
output(2, 82) <= input(19);
output(2, 83) <= input(20);
output(2, 84) <= input(21);
output(2, 85) <= input(22);
output(2, 86) <= input(23);
output(2, 87) <= input(24);
output(2, 88) <= input(25);
output(2, 89) <= input(26);
output(2, 90) <= input(27);
output(2, 91) <= input(28);
output(2, 92) <= input(29);
output(2, 93) <= input(30);
output(2, 94) <= input(31);
output(2, 95) <= input(33);
output(2, 96) <= input(2);
output(2, 97) <= input(3);
output(2, 98) <= input(4);
output(2, 99) <= input(5);
output(2, 100) <= input(6);
output(2, 101) <= input(7);
output(2, 102) <= input(8);
output(2, 103) <= input(9);
output(2, 104) <= input(10);
output(2, 105) <= input(11);
output(2, 106) <= input(12);
output(2, 107) <= input(13);
output(2, 108) <= input(14);
output(2, 109) <= input(15);
output(2, 110) <= input(32);
output(2, 111) <= input(34);
output(2, 112) <= input(18);
output(2, 113) <= input(19);
output(2, 114) <= input(20);
output(2, 115) <= input(21);
output(2, 116) <= input(22);
output(2, 117) <= input(23);
output(2, 118) <= input(24);
output(2, 119) <= input(25);
output(2, 120) <= input(26);
output(2, 121) <= input(27);
output(2, 122) <= input(28);
output(2, 123) <= input(29);
output(2, 124) <= input(30);
output(2, 125) <= input(31);
output(2, 126) <= input(33);
output(2, 127) <= input(35);
output(2, 128) <= input(18);
output(2, 129) <= input(19);
output(2, 130) <= input(20);
output(2, 131) <= input(21);
output(2, 132) <= input(22);
output(2, 133) <= input(23);
output(2, 134) <= input(24);
output(2, 135) <= input(25);
output(2, 136) <= input(26);
output(2, 137) <= input(27);
output(2, 138) <= input(28);
output(2, 139) <= input(29);
output(2, 140) <= input(30);
output(2, 141) <= input(31);
output(2, 142) <= input(33);
output(2, 143) <= input(35);
output(2, 144) <= input(3);
output(2, 145) <= input(4);
output(2, 146) <= input(5);
output(2, 147) <= input(6);
output(2, 148) <= input(7);
output(2, 149) <= input(8);
output(2, 150) <= input(9);
output(2, 151) <= input(10);
output(2, 152) <= input(11);
output(2, 153) <= input(12);
output(2, 154) <= input(13);
output(2, 155) <= input(14);
output(2, 156) <= input(15);
output(2, 157) <= input(32);
output(2, 158) <= input(34);
output(2, 159) <= input(36);
output(2, 160) <= input(3);
output(2, 161) <= input(4);
output(2, 162) <= input(5);
output(2, 163) <= input(6);
output(2, 164) <= input(7);
output(2, 165) <= input(8);
output(2, 166) <= input(9);
output(2, 167) <= input(10);
output(2, 168) <= input(11);
output(2, 169) <= input(12);
output(2, 170) <= input(13);
output(2, 171) <= input(14);
output(2, 172) <= input(15);
output(2, 173) <= input(32);
output(2, 174) <= input(34);
output(2, 175) <= input(36);
output(2, 176) <= input(19);
output(2, 177) <= input(20);
output(2, 178) <= input(21);
output(2, 179) <= input(22);
output(2, 180) <= input(23);
output(2, 181) <= input(24);
output(2, 182) <= input(25);
output(2, 183) <= input(26);
output(2, 184) <= input(27);
output(2, 185) <= input(28);
output(2, 186) <= input(29);
output(2, 187) <= input(30);
output(2, 188) <= input(31);
output(2, 189) <= input(33);
output(2, 190) <= input(35);
output(2, 191) <= input(37);
output(2, 192) <= input(4);
output(2, 193) <= input(5);
output(2, 194) <= input(6);
output(2, 195) <= input(7);
output(2, 196) <= input(8);
output(2, 197) <= input(9);
output(2, 198) <= input(10);
output(2, 199) <= input(11);
output(2, 200) <= input(12);
output(2, 201) <= input(13);
output(2, 202) <= input(14);
output(2, 203) <= input(15);
output(2, 204) <= input(32);
output(2, 205) <= input(34);
output(2, 206) <= input(36);
output(2, 207) <= input(38);
output(2, 208) <= input(4);
output(2, 209) <= input(5);
output(2, 210) <= input(6);
output(2, 211) <= input(7);
output(2, 212) <= input(8);
output(2, 213) <= input(9);
output(2, 214) <= input(10);
output(2, 215) <= input(11);
output(2, 216) <= input(12);
output(2, 217) <= input(13);
output(2, 218) <= input(14);
output(2, 219) <= input(15);
output(2, 220) <= input(32);
output(2, 221) <= input(34);
output(2, 222) <= input(36);
output(2, 223) <= input(38);
output(2, 224) <= input(20);
output(2, 225) <= input(21);
output(2, 226) <= input(22);
output(2, 227) <= input(23);
output(2, 228) <= input(24);
output(2, 229) <= input(25);
output(2, 230) <= input(26);
output(2, 231) <= input(27);
output(2, 232) <= input(28);
output(2, 233) <= input(29);
output(2, 234) <= input(30);
output(2, 235) <= input(31);
output(2, 236) <= input(33);
output(2, 237) <= input(35);
output(2, 238) <= input(37);
output(2, 239) <= input(39);
output(2, 240) <= input(5);
output(2, 241) <= input(6);
output(2, 242) <= input(7);
output(2, 243) <= input(8);
output(2, 244) <= input(9);
output(2, 245) <= input(10);
output(2, 246) <= input(11);
output(2, 247) <= input(12);
output(2, 248) <= input(13);
output(2, 249) <= input(14);
output(2, 250) <= input(15);
output(2, 251) <= input(32);
output(2, 252) <= input(34);
output(2, 253) <= input(36);
output(2, 254) <= input(38);
output(2, 255) <= input(40);
output(3, 0) <= input(0);
output(3, 1) <= input(1);
output(3, 2) <= input(2);
output(3, 3) <= input(3);
output(3, 4) <= input(4);
output(3, 5) <= input(5);
output(3, 6) <= input(6);
output(3, 7) <= input(7);
output(3, 8) <= input(8);
output(3, 9) <= input(9);
output(3, 10) <= input(10);
output(3, 11) <= input(11);
output(3, 12) <= input(12);
output(3, 13) <= input(13);
output(3, 14) <= input(14);
output(3, 15) <= input(15);
output(3, 16) <= input(16);
output(3, 17) <= input(17);
output(3, 18) <= input(18);
output(3, 19) <= input(19);
output(3, 20) <= input(20);
output(3, 21) <= input(21);
output(3, 22) <= input(22);
output(3, 23) <= input(23);
output(3, 24) <= input(24);
output(3, 25) <= input(25);
output(3, 26) <= input(26);
output(3, 27) <= input(27);
output(3, 28) <= input(28);
output(3, 29) <= input(29);
output(3, 30) <= input(30);
output(3, 31) <= input(31);
output(3, 32) <= input(1);
output(3, 33) <= input(2);
output(3, 34) <= input(3);
output(3, 35) <= input(4);
output(3, 36) <= input(5);
output(3, 37) <= input(6);
output(3, 38) <= input(7);
output(3, 39) <= input(8);
output(3, 40) <= input(9);
output(3, 41) <= input(10);
output(3, 42) <= input(11);
output(3, 43) <= input(12);
output(3, 44) <= input(13);
output(3, 45) <= input(14);
output(3, 46) <= input(15);
output(3, 47) <= input(32);
output(3, 48) <= input(17);
output(3, 49) <= input(18);
output(3, 50) <= input(19);
output(3, 51) <= input(20);
output(3, 52) <= input(21);
output(3, 53) <= input(22);
output(3, 54) <= input(23);
output(3, 55) <= input(24);
output(3, 56) <= input(25);
output(3, 57) <= input(26);
output(3, 58) <= input(27);
output(3, 59) <= input(28);
output(3, 60) <= input(29);
output(3, 61) <= input(30);
output(3, 62) <= input(31);
output(3, 63) <= input(33);
output(3, 64) <= input(17);
output(3, 65) <= input(18);
output(3, 66) <= input(19);
output(3, 67) <= input(20);
output(3, 68) <= input(21);
output(3, 69) <= input(22);
output(3, 70) <= input(23);
output(3, 71) <= input(24);
output(3, 72) <= input(25);
output(3, 73) <= input(26);
output(3, 74) <= input(27);
output(3, 75) <= input(28);
output(3, 76) <= input(29);
output(3, 77) <= input(30);
output(3, 78) <= input(31);
output(3, 79) <= input(33);
output(3, 80) <= input(2);
output(3, 81) <= input(3);
output(3, 82) <= input(4);
output(3, 83) <= input(5);
output(3, 84) <= input(6);
output(3, 85) <= input(7);
output(3, 86) <= input(8);
output(3, 87) <= input(9);
output(3, 88) <= input(10);
output(3, 89) <= input(11);
output(3, 90) <= input(12);
output(3, 91) <= input(13);
output(3, 92) <= input(14);
output(3, 93) <= input(15);
output(3, 94) <= input(32);
output(3, 95) <= input(34);
output(3, 96) <= input(18);
output(3, 97) <= input(19);
output(3, 98) <= input(20);
output(3, 99) <= input(21);
output(3, 100) <= input(22);
output(3, 101) <= input(23);
output(3, 102) <= input(24);
output(3, 103) <= input(25);
output(3, 104) <= input(26);
output(3, 105) <= input(27);
output(3, 106) <= input(28);
output(3, 107) <= input(29);
output(3, 108) <= input(30);
output(3, 109) <= input(31);
output(3, 110) <= input(33);
output(3, 111) <= input(35);
output(3, 112) <= input(3);
output(3, 113) <= input(4);
output(3, 114) <= input(5);
output(3, 115) <= input(6);
output(3, 116) <= input(7);
output(3, 117) <= input(8);
output(3, 118) <= input(9);
output(3, 119) <= input(10);
output(3, 120) <= input(11);
output(3, 121) <= input(12);
output(3, 122) <= input(13);
output(3, 123) <= input(14);
output(3, 124) <= input(15);
output(3, 125) <= input(32);
output(3, 126) <= input(34);
output(3, 127) <= input(36);
output(3, 128) <= input(3);
output(3, 129) <= input(4);
output(3, 130) <= input(5);
output(3, 131) <= input(6);
output(3, 132) <= input(7);
output(3, 133) <= input(8);
output(3, 134) <= input(9);
output(3, 135) <= input(10);
output(3, 136) <= input(11);
output(3, 137) <= input(12);
output(3, 138) <= input(13);
output(3, 139) <= input(14);
output(3, 140) <= input(15);
output(3, 141) <= input(32);
output(3, 142) <= input(34);
output(3, 143) <= input(36);
output(3, 144) <= input(19);
output(3, 145) <= input(20);
output(3, 146) <= input(21);
output(3, 147) <= input(22);
output(3, 148) <= input(23);
output(3, 149) <= input(24);
output(3, 150) <= input(25);
output(3, 151) <= input(26);
output(3, 152) <= input(27);
output(3, 153) <= input(28);
output(3, 154) <= input(29);
output(3, 155) <= input(30);
output(3, 156) <= input(31);
output(3, 157) <= input(33);
output(3, 158) <= input(35);
output(3, 159) <= input(37);
output(3, 160) <= input(4);
output(3, 161) <= input(5);
output(3, 162) <= input(6);
output(3, 163) <= input(7);
output(3, 164) <= input(8);
output(3, 165) <= input(9);
output(3, 166) <= input(10);
output(3, 167) <= input(11);
output(3, 168) <= input(12);
output(3, 169) <= input(13);
output(3, 170) <= input(14);
output(3, 171) <= input(15);
output(3, 172) <= input(32);
output(3, 173) <= input(34);
output(3, 174) <= input(36);
output(3, 175) <= input(38);
output(3, 176) <= input(20);
output(3, 177) <= input(21);
output(3, 178) <= input(22);
output(3, 179) <= input(23);
output(3, 180) <= input(24);
output(3, 181) <= input(25);
output(3, 182) <= input(26);
output(3, 183) <= input(27);
output(3, 184) <= input(28);
output(3, 185) <= input(29);
output(3, 186) <= input(30);
output(3, 187) <= input(31);
output(3, 188) <= input(33);
output(3, 189) <= input(35);
output(3, 190) <= input(37);
output(3, 191) <= input(39);
output(3, 192) <= input(20);
output(3, 193) <= input(21);
output(3, 194) <= input(22);
output(3, 195) <= input(23);
output(3, 196) <= input(24);
output(3, 197) <= input(25);
output(3, 198) <= input(26);
output(3, 199) <= input(27);
output(3, 200) <= input(28);
output(3, 201) <= input(29);
output(3, 202) <= input(30);
output(3, 203) <= input(31);
output(3, 204) <= input(33);
output(3, 205) <= input(35);
output(3, 206) <= input(37);
output(3, 207) <= input(39);
output(3, 208) <= input(5);
output(3, 209) <= input(6);
output(3, 210) <= input(7);
output(3, 211) <= input(8);
output(3, 212) <= input(9);
output(3, 213) <= input(10);
output(3, 214) <= input(11);
output(3, 215) <= input(12);
output(3, 216) <= input(13);
output(3, 217) <= input(14);
output(3, 218) <= input(15);
output(3, 219) <= input(32);
output(3, 220) <= input(34);
output(3, 221) <= input(36);
output(3, 222) <= input(38);
output(3, 223) <= input(40);
output(3, 224) <= input(21);
output(3, 225) <= input(22);
output(3, 226) <= input(23);
output(3, 227) <= input(24);
output(3, 228) <= input(25);
output(3, 229) <= input(26);
output(3, 230) <= input(27);
output(3, 231) <= input(28);
output(3, 232) <= input(29);
output(3, 233) <= input(30);
output(3, 234) <= input(31);
output(3, 235) <= input(33);
output(3, 236) <= input(35);
output(3, 237) <= input(37);
output(3, 238) <= input(39);
output(3, 239) <= input(41);
output(3, 240) <= input(6);
output(3, 241) <= input(7);
output(3, 242) <= input(8);
output(3, 243) <= input(9);
output(3, 244) <= input(10);
output(3, 245) <= input(11);
output(3, 246) <= input(12);
output(3, 247) <= input(13);
output(3, 248) <= input(14);
output(3, 249) <= input(15);
output(3, 250) <= input(32);
output(3, 251) <= input(34);
output(3, 252) <= input(36);
output(3, 253) <= input(38);
output(3, 254) <= input(40);
output(3, 255) <= input(42);
output(4, 0) <= input(0);
output(4, 1) <= input(1);
output(4, 2) <= input(2);
output(4, 3) <= input(3);
output(4, 4) <= input(4);
output(4, 5) <= input(5);
output(4, 6) <= input(6);
output(4, 7) <= input(7);
output(4, 8) <= input(8);
output(4, 9) <= input(9);
output(4, 10) <= input(10);
output(4, 11) <= input(11);
output(4, 12) <= input(12);
output(4, 13) <= input(13);
output(4, 14) <= input(14);
output(4, 15) <= input(15);
output(4, 16) <= input(16);
output(4, 17) <= input(17);
output(4, 18) <= input(18);
output(4, 19) <= input(19);
output(4, 20) <= input(20);
output(4, 21) <= input(21);
output(4, 22) <= input(22);
output(4, 23) <= input(23);
output(4, 24) <= input(24);
output(4, 25) <= input(25);
output(4, 26) <= input(26);
output(4, 27) <= input(27);
output(4, 28) <= input(28);
output(4, 29) <= input(29);
output(4, 30) <= input(30);
output(4, 31) <= input(31);
output(4, 32) <= input(1);
output(4, 33) <= input(2);
output(4, 34) <= input(3);
output(4, 35) <= input(4);
output(4, 36) <= input(5);
output(4, 37) <= input(6);
output(4, 38) <= input(7);
output(4, 39) <= input(8);
output(4, 40) <= input(9);
output(4, 41) <= input(10);
output(4, 42) <= input(11);
output(4, 43) <= input(12);
output(4, 44) <= input(13);
output(4, 45) <= input(14);
output(4, 46) <= input(15);
output(4, 47) <= input(32);
output(4, 48) <= input(17);
output(4, 49) <= input(18);
output(4, 50) <= input(19);
output(4, 51) <= input(20);
output(4, 52) <= input(21);
output(4, 53) <= input(22);
output(4, 54) <= input(23);
output(4, 55) <= input(24);
output(4, 56) <= input(25);
output(4, 57) <= input(26);
output(4, 58) <= input(27);
output(4, 59) <= input(28);
output(4, 60) <= input(29);
output(4, 61) <= input(30);
output(4, 62) <= input(31);
output(4, 63) <= input(33);
output(4, 64) <= input(2);
output(4, 65) <= input(3);
output(4, 66) <= input(4);
output(4, 67) <= input(5);
output(4, 68) <= input(6);
output(4, 69) <= input(7);
output(4, 70) <= input(8);
output(4, 71) <= input(9);
output(4, 72) <= input(10);
output(4, 73) <= input(11);
output(4, 74) <= input(12);
output(4, 75) <= input(13);
output(4, 76) <= input(14);
output(4, 77) <= input(15);
output(4, 78) <= input(32);
output(4, 79) <= input(34);
output(4, 80) <= input(18);
output(4, 81) <= input(19);
output(4, 82) <= input(20);
output(4, 83) <= input(21);
output(4, 84) <= input(22);
output(4, 85) <= input(23);
output(4, 86) <= input(24);
output(4, 87) <= input(25);
output(4, 88) <= input(26);
output(4, 89) <= input(27);
output(4, 90) <= input(28);
output(4, 91) <= input(29);
output(4, 92) <= input(30);
output(4, 93) <= input(31);
output(4, 94) <= input(33);
output(4, 95) <= input(35);
output(4, 96) <= input(3);
output(4, 97) <= input(4);
output(4, 98) <= input(5);
output(4, 99) <= input(6);
output(4, 100) <= input(7);
output(4, 101) <= input(8);
output(4, 102) <= input(9);
output(4, 103) <= input(10);
output(4, 104) <= input(11);
output(4, 105) <= input(12);
output(4, 106) <= input(13);
output(4, 107) <= input(14);
output(4, 108) <= input(15);
output(4, 109) <= input(32);
output(4, 110) <= input(34);
output(4, 111) <= input(36);
output(4, 112) <= input(19);
output(4, 113) <= input(20);
output(4, 114) <= input(21);
output(4, 115) <= input(22);
output(4, 116) <= input(23);
output(4, 117) <= input(24);
output(4, 118) <= input(25);
output(4, 119) <= input(26);
output(4, 120) <= input(27);
output(4, 121) <= input(28);
output(4, 122) <= input(29);
output(4, 123) <= input(30);
output(4, 124) <= input(31);
output(4, 125) <= input(33);
output(4, 126) <= input(35);
output(4, 127) <= input(37);
output(4, 128) <= input(19);
output(4, 129) <= input(20);
output(4, 130) <= input(21);
output(4, 131) <= input(22);
output(4, 132) <= input(23);
output(4, 133) <= input(24);
output(4, 134) <= input(25);
output(4, 135) <= input(26);
output(4, 136) <= input(27);
output(4, 137) <= input(28);
output(4, 138) <= input(29);
output(4, 139) <= input(30);
output(4, 140) <= input(31);
output(4, 141) <= input(33);
output(4, 142) <= input(35);
output(4, 143) <= input(37);
output(4, 144) <= input(4);
output(4, 145) <= input(5);
output(4, 146) <= input(6);
output(4, 147) <= input(7);
output(4, 148) <= input(8);
output(4, 149) <= input(9);
output(4, 150) <= input(10);
output(4, 151) <= input(11);
output(4, 152) <= input(12);
output(4, 153) <= input(13);
output(4, 154) <= input(14);
output(4, 155) <= input(15);
output(4, 156) <= input(32);
output(4, 157) <= input(34);
output(4, 158) <= input(36);
output(4, 159) <= input(38);
output(4, 160) <= input(20);
output(4, 161) <= input(21);
output(4, 162) <= input(22);
output(4, 163) <= input(23);
output(4, 164) <= input(24);
output(4, 165) <= input(25);
output(4, 166) <= input(26);
output(4, 167) <= input(27);
output(4, 168) <= input(28);
output(4, 169) <= input(29);
output(4, 170) <= input(30);
output(4, 171) <= input(31);
output(4, 172) <= input(33);
output(4, 173) <= input(35);
output(4, 174) <= input(37);
output(4, 175) <= input(39);
output(4, 176) <= input(5);
output(4, 177) <= input(6);
output(4, 178) <= input(7);
output(4, 179) <= input(8);
output(4, 180) <= input(9);
output(4, 181) <= input(10);
output(4, 182) <= input(11);
output(4, 183) <= input(12);
output(4, 184) <= input(13);
output(4, 185) <= input(14);
output(4, 186) <= input(15);
output(4, 187) <= input(32);
output(4, 188) <= input(34);
output(4, 189) <= input(36);
output(4, 190) <= input(38);
output(4, 191) <= input(40);
output(4, 192) <= input(21);
output(4, 193) <= input(22);
output(4, 194) <= input(23);
output(4, 195) <= input(24);
output(4, 196) <= input(25);
output(4, 197) <= input(26);
output(4, 198) <= input(27);
output(4, 199) <= input(28);
output(4, 200) <= input(29);
output(4, 201) <= input(30);
output(4, 202) <= input(31);
output(4, 203) <= input(33);
output(4, 204) <= input(35);
output(4, 205) <= input(37);
output(4, 206) <= input(39);
output(4, 207) <= input(41);
output(4, 208) <= input(6);
output(4, 209) <= input(7);
output(4, 210) <= input(8);
output(4, 211) <= input(9);
output(4, 212) <= input(10);
output(4, 213) <= input(11);
output(4, 214) <= input(12);
output(4, 215) <= input(13);
output(4, 216) <= input(14);
output(4, 217) <= input(15);
output(4, 218) <= input(32);
output(4, 219) <= input(34);
output(4, 220) <= input(36);
output(4, 221) <= input(38);
output(4, 222) <= input(40);
output(4, 223) <= input(42);
output(4, 224) <= input(22);
output(4, 225) <= input(23);
output(4, 226) <= input(24);
output(4, 227) <= input(25);
output(4, 228) <= input(26);
output(4, 229) <= input(27);
output(4, 230) <= input(28);
output(4, 231) <= input(29);
output(4, 232) <= input(30);
output(4, 233) <= input(31);
output(4, 234) <= input(33);
output(4, 235) <= input(35);
output(4, 236) <= input(37);
output(4, 237) <= input(39);
output(4, 238) <= input(41);
output(4, 239) <= input(43);
output(4, 240) <= input(7);
output(4, 241) <= input(8);
output(4, 242) <= input(9);
output(4, 243) <= input(10);
output(4, 244) <= input(11);
output(4, 245) <= input(12);
output(4, 246) <= input(13);
output(4, 247) <= input(14);
output(4, 248) <= input(15);
output(4, 249) <= input(32);
output(4, 250) <= input(34);
output(4, 251) <= input(36);
output(4, 252) <= input(38);
output(4, 253) <= input(40);
output(4, 254) <= input(42);
output(4, 255) <= input(44);
output(5, 0) <= input(16);
output(5, 1) <= input(17);
output(5, 2) <= input(18);
output(5, 3) <= input(19);
output(5, 4) <= input(20);
output(5, 5) <= input(21);
output(5, 6) <= input(22);
output(5, 7) <= input(23);
output(5, 8) <= input(24);
output(5, 9) <= input(25);
output(5, 10) <= input(26);
output(5, 11) <= input(27);
output(5, 12) <= input(28);
output(5, 13) <= input(29);
output(5, 14) <= input(30);
output(5, 15) <= input(31);
output(5, 16) <= input(1);
output(5, 17) <= input(2);
output(5, 18) <= input(3);
output(5, 19) <= input(4);
output(5, 20) <= input(5);
output(5, 21) <= input(6);
output(5, 22) <= input(7);
output(5, 23) <= input(8);
output(5, 24) <= input(9);
output(5, 25) <= input(10);
output(5, 26) <= input(11);
output(5, 27) <= input(12);
output(5, 28) <= input(13);
output(5, 29) <= input(14);
output(5, 30) <= input(15);
output(5, 31) <= input(32);
output(5, 32) <= input(17);
output(5, 33) <= input(18);
output(5, 34) <= input(19);
output(5, 35) <= input(20);
output(5, 36) <= input(21);
output(5, 37) <= input(22);
output(5, 38) <= input(23);
output(5, 39) <= input(24);
output(5, 40) <= input(25);
output(5, 41) <= input(26);
output(5, 42) <= input(27);
output(5, 43) <= input(28);
output(5, 44) <= input(29);
output(5, 45) <= input(30);
output(5, 46) <= input(31);
output(5, 47) <= input(33);
output(5, 48) <= input(2);
output(5, 49) <= input(3);
output(5, 50) <= input(4);
output(5, 51) <= input(5);
output(5, 52) <= input(6);
output(5, 53) <= input(7);
output(5, 54) <= input(8);
output(5, 55) <= input(9);
output(5, 56) <= input(10);
output(5, 57) <= input(11);
output(5, 58) <= input(12);
output(5, 59) <= input(13);
output(5, 60) <= input(14);
output(5, 61) <= input(15);
output(5, 62) <= input(32);
output(5, 63) <= input(34);
output(5, 64) <= input(18);
output(5, 65) <= input(19);
output(5, 66) <= input(20);
output(5, 67) <= input(21);
output(5, 68) <= input(22);
output(5, 69) <= input(23);
output(5, 70) <= input(24);
output(5, 71) <= input(25);
output(5, 72) <= input(26);
output(5, 73) <= input(27);
output(5, 74) <= input(28);
output(5, 75) <= input(29);
output(5, 76) <= input(30);
output(5, 77) <= input(31);
output(5, 78) <= input(33);
output(5, 79) <= input(35);
output(5, 80) <= input(3);
output(5, 81) <= input(4);
output(5, 82) <= input(5);
output(5, 83) <= input(6);
output(5, 84) <= input(7);
output(5, 85) <= input(8);
output(5, 86) <= input(9);
output(5, 87) <= input(10);
output(5, 88) <= input(11);
output(5, 89) <= input(12);
output(5, 90) <= input(13);
output(5, 91) <= input(14);
output(5, 92) <= input(15);
output(5, 93) <= input(32);
output(5, 94) <= input(34);
output(5, 95) <= input(36);
output(5, 96) <= input(19);
output(5, 97) <= input(20);
output(5, 98) <= input(21);
output(5, 99) <= input(22);
output(5, 100) <= input(23);
output(5, 101) <= input(24);
output(5, 102) <= input(25);
output(5, 103) <= input(26);
output(5, 104) <= input(27);
output(5, 105) <= input(28);
output(5, 106) <= input(29);
output(5, 107) <= input(30);
output(5, 108) <= input(31);
output(5, 109) <= input(33);
output(5, 110) <= input(35);
output(5, 111) <= input(37);
output(5, 112) <= input(4);
output(5, 113) <= input(5);
output(5, 114) <= input(6);
output(5, 115) <= input(7);
output(5, 116) <= input(8);
output(5, 117) <= input(9);
output(5, 118) <= input(10);
output(5, 119) <= input(11);
output(5, 120) <= input(12);
output(5, 121) <= input(13);
output(5, 122) <= input(14);
output(5, 123) <= input(15);
output(5, 124) <= input(32);
output(5, 125) <= input(34);
output(5, 126) <= input(36);
output(5, 127) <= input(38);
output(5, 128) <= input(20);
output(5, 129) <= input(21);
output(5, 130) <= input(22);
output(5, 131) <= input(23);
output(5, 132) <= input(24);
output(5, 133) <= input(25);
output(5, 134) <= input(26);
output(5, 135) <= input(27);
output(5, 136) <= input(28);
output(5, 137) <= input(29);
output(5, 138) <= input(30);
output(5, 139) <= input(31);
output(5, 140) <= input(33);
output(5, 141) <= input(35);
output(5, 142) <= input(37);
output(5, 143) <= input(39);
output(5, 144) <= input(5);
output(5, 145) <= input(6);
output(5, 146) <= input(7);
output(5, 147) <= input(8);
output(5, 148) <= input(9);
output(5, 149) <= input(10);
output(5, 150) <= input(11);
output(5, 151) <= input(12);
output(5, 152) <= input(13);
output(5, 153) <= input(14);
output(5, 154) <= input(15);
output(5, 155) <= input(32);
output(5, 156) <= input(34);
output(5, 157) <= input(36);
output(5, 158) <= input(38);
output(5, 159) <= input(40);
output(5, 160) <= input(21);
output(5, 161) <= input(22);
output(5, 162) <= input(23);
output(5, 163) <= input(24);
output(5, 164) <= input(25);
output(5, 165) <= input(26);
output(5, 166) <= input(27);
output(5, 167) <= input(28);
output(5, 168) <= input(29);
output(5, 169) <= input(30);
output(5, 170) <= input(31);
output(5, 171) <= input(33);
output(5, 172) <= input(35);
output(5, 173) <= input(37);
output(5, 174) <= input(39);
output(5, 175) <= input(41);
output(5, 176) <= input(6);
output(5, 177) <= input(7);
output(5, 178) <= input(8);
output(5, 179) <= input(9);
output(5, 180) <= input(10);
output(5, 181) <= input(11);
output(5, 182) <= input(12);
output(5, 183) <= input(13);
output(5, 184) <= input(14);
output(5, 185) <= input(15);
output(5, 186) <= input(32);
output(5, 187) <= input(34);
output(5, 188) <= input(36);
output(5, 189) <= input(38);
output(5, 190) <= input(40);
output(5, 191) <= input(42);
output(5, 192) <= input(22);
output(5, 193) <= input(23);
output(5, 194) <= input(24);
output(5, 195) <= input(25);
output(5, 196) <= input(26);
output(5, 197) <= input(27);
output(5, 198) <= input(28);
output(5, 199) <= input(29);
output(5, 200) <= input(30);
output(5, 201) <= input(31);
output(5, 202) <= input(33);
output(5, 203) <= input(35);
output(5, 204) <= input(37);
output(5, 205) <= input(39);
output(5, 206) <= input(41);
output(5, 207) <= input(43);
output(5, 208) <= input(7);
output(5, 209) <= input(8);
output(5, 210) <= input(9);
output(5, 211) <= input(10);
output(5, 212) <= input(11);
output(5, 213) <= input(12);
output(5, 214) <= input(13);
output(5, 215) <= input(14);
output(5, 216) <= input(15);
output(5, 217) <= input(32);
output(5, 218) <= input(34);
output(5, 219) <= input(36);
output(5, 220) <= input(38);
output(5, 221) <= input(40);
output(5, 222) <= input(42);
output(5, 223) <= input(44);
output(5, 224) <= input(23);
output(5, 225) <= input(24);
output(5, 226) <= input(25);
output(5, 227) <= input(26);
output(5, 228) <= input(27);
output(5, 229) <= input(28);
output(5, 230) <= input(29);
output(5, 231) <= input(30);
output(5, 232) <= input(31);
output(5, 233) <= input(33);
output(5, 234) <= input(35);
output(5, 235) <= input(37);
output(5, 236) <= input(39);
output(5, 237) <= input(41);
output(5, 238) <= input(43);
output(5, 239) <= input(45);
output(5, 240) <= input(8);
output(5, 241) <= input(9);
output(5, 242) <= input(10);
output(5, 243) <= input(11);
output(5, 244) <= input(12);
output(5, 245) <= input(13);
output(5, 246) <= input(14);
output(5, 247) <= input(15);
output(5, 248) <= input(32);
output(5, 249) <= input(34);
output(5, 250) <= input(36);
output(5, 251) <= input(38);
output(5, 252) <= input(40);
output(5, 253) <= input(42);
output(5, 254) <= input(44);
output(5, 255) <= input(46);
when "1111" =>
output(0, 0) <= input(0);
output(0, 1) <= input(1);
output(0, 2) <= input(2);
output(0, 3) <= input(3);
output(0, 4) <= input(4);
output(0, 5) <= input(5);
output(0, 6) <= input(6);
output(0, 7) <= input(7);
output(0, 8) <= input(8);
output(0, 9) <= input(9);
output(0, 10) <= input(10);
output(0, 11) <= input(11);
output(0, 12) <= input(12);
output(0, 13) <= input(13);
output(0, 14) <= input(14);
output(0, 15) <= input(15);
output(0, 16) <= input(16);
output(0, 17) <= input(17);
output(0, 18) <= input(18);
output(0, 19) <= input(19);
output(0, 20) <= input(20);
output(0, 21) <= input(21);
output(0, 22) <= input(22);
output(0, 23) <= input(23);
output(0, 24) <= input(24);
output(0, 25) <= input(25);
output(0, 26) <= input(26);
output(0, 27) <= input(27);
output(0, 28) <= input(28);
output(0, 29) <= input(29);
output(0, 30) <= input(30);
output(0, 31) <= input(31);
output(0, 32) <= input(1);
output(0, 33) <= input(2);
output(0, 34) <= input(3);
output(0, 35) <= input(4);
output(0, 36) <= input(5);
output(0, 37) <= input(6);
output(0, 38) <= input(7);
output(0, 39) <= input(8);
output(0, 40) <= input(9);
output(0, 41) <= input(10);
output(0, 42) <= input(11);
output(0, 43) <= input(12);
output(0, 44) <= input(13);
output(0, 45) <= input(14);
output(0, 46) <= input(15);
output(0, 47) <= input(32);
output(0, 48) <= input(17);
output(0, 49) <= input(18);
output(0, 50) <= input(19);
output(0, 51) <= input(20);
output(0, 52) <= input(21);
output(0, 53) <= input(22);
output(0, 54) <= input(23);
output(0, 55) <= input(24);
output(0, 56) <= input(25);
output(0, 57) <= input(26);
output(0, 58) <= input(27);
output(0, 59) <= input(28);
output(0, 60) <= input(29);
output(0, 61) <= input(30);
output(0, 62) <= input(31);
output(0, 63) <= input(33);
output(0, 64) <= input(2);
output(0, 65) <= input(3);
output(0, 66) <= input(4);
output(0, 67) <= input(5);
output(0, 68) <= input(6);
output(0, 69) <= input(7);
output(0, 70) <= input(8);
output(0, 71) <= input(9);
output(0, 72) <= input(10);
output(0, 73) <= input(11);
output(0, 74) <= input(12);
output(0, 75) <= input(13);
output(0, 76) <= input(14);
output(0, 77) <= input(15);
output(0, 78) <= input(32);
output(0, 79) <= input(34);
output(0, 80) <= input(18);
output(0, 81) <= input(19);
output(0, 82) <= input(20);
output(0, 83) <= input(21);
output(0, 84) <= input(22);
output(0, 85) <= input(23);
output(0, 86) <= input(24);
output(0, 87) <= input(25);
output(0, 88) <= input(26);
output(0, 89) <= input(27);
output(0, 90) <= input(28);
output(0, 91) <= input(29);
output(0, 92) <= input(30);
output(0, 93) <= input(31);
output(0, 94) <= input(33);
output(0, 95) <= input(35);
output(0, 96) <= input(3);
output(0, 97) <= input(4);
output(0, 98) <= input(5);
output(0, 99) <= input(6);
output(0, 100) <= input(7);
output(0, 101) <= input(8);
output(0, 102) <= input(9);
output(0, 103) <= input(10);
output(0, 104) <= input(11);
output(0, 105) <= input(12);
output(0, 106) <= input(13);
output(0, 107) <= input(14);
output(0, 108) <= input(15);
output(0, 109) <= input(32);
output(0, 110) <= input(34);
output(0, 111) <= input(36);
output(0, 112) <= input(4);
output(0, 113) <= input(5);
output(0, 114) <= input(6);
output(0, 115) <= input(7);
output(0, 116) <= input(8);
output(0, 117) <= input(9);
output(0, 118) <= input(10);
output(0, 119) <= input(11);
output(0, 120) <= input(12);
output(0, 121) <= input(13);
output(0, 122) <= input(14);
output(0, 123) <= input(15);
output(0, 124) <= input(32);
output(0, 125) <= input(34);
output(0, 126) <= input(36);
output(0, 127) <= input(37);
output(0, 128) <= input(20);
output(0, 129) <= input(21);
output(0, 130) <= input(22);
output(0, 131) <= input(23);
output(0, 132) <= input(24);
output(0, 133) <= input(25);
output(0, 134) <= input(26);
output(0, 135) <= input(27);
output(0, 136) <= input(28);
output(0, 137) <= input(29);
output(0, 138) <= input(30);
output(0, 139) <= input(31);
output(0, 140) <= input(33);
output(0, 141) <= input(35);
output(0, 142) <= input(38);
output(0, 143) <= input(39);
output(0, 144) <= input(5);
output(0, 145) <= input(6);
output(0, 146) <= input(7);
output(0, 147) <= input(8);
output(0, 148) <= input(9);
output(0, 149) <= input(10);
output(0, 150) <= input(11);
output(0, 151) <= input(12);
output(0, 152) <= input(13);
output(0, 153) <= input(14);
output(0, 154) <= input(15);
output(0, 155) <= input(32);
output(0, 156) <= input(34);
output(0, 157) <= input(36);
output(0, 158) <= input(37);
output(0, 159) <= input(40);
output(0, 160) <= input(21);
output(0, 161) <= input(22);
output(0, 162) <= input(23);
output(0, 163) <= input(24);
output(0, 164) <= input(25);
output(0, 165) <= input(26);
output(0, 166) <= input(27);
output(0, 167) <= input(28);
output(0, 168) <= input(29);
output(0, 169) <= input(30);
output(0, 170) <= input(31);
output(0, 171) <= input(33);
output(0, 172) <= input(35);
output(0, 173) <= input(38);
output(0, 174) <= input(39);
output(0, 175) <= input(41);
output(0, 176) <= input(6);
output(0, 177) <= input(7);
output(0, 178) <= input(8);
output(0, 179) <= input(9);
output(0, 180) <= input(10);
output(0, 181) <= input(11);
output(0, 182) <= input(12);
output(0, 183) <= input(13);
output(0, 184) <= input(14);
output(0, 185) <= input(15);
output(0, 186) <= input(32);
output(0, 187) <= input(34);
output(0, 188) <= input(36);
output(0, 189) <= input(37);
output(0, 190) <= input(40);
output(0, 191) <= input(42);
output(0, 192) <= input(22);
output(0, 193) <= input(23);
output(0, 194) <= input(24);
output(0, 195) <= input(25);
output(0, 196) <= input(26);
output(0, 197) <= input(27);
output(0, 198) <= input(28);
output(0, 199) <= input(29);
output(0, 200) <= input(30);
output(0, 201) <= input(31);
output(0, 202) <= input(33);
output(0, 203) <= input(35);
output(0, 204) <= input(38);
output(0, 205) <= input(39);
output(0, 206) <= input(41);
output(0, 207) <= input(43);
output(0, 208) <= input(7);
output(0, 209) <= input(8);
output(0, 210) <= input(9);
output(0, 211) <= input(10);
output(0, 212) <= input(11);
output(0, 213) <= input(12);
output(0, 214) <= input(13);
output(0, 215) <= input(14);
output(0, 216) <= input(15);
output(0, 217) <= input(32);
output(0, 218) <= input(34);
output(0, 219) <= input(36);
output(0, 220) <= input(37);
output(0, 221) <= input(40);
output(0, 222) <= input(42);
output(0, 223) <= input(44);
output(0, 224) <= input(23);
output(0, 225) <= input(24);
output(0, 226) <= input(25);
output(0, 227) <= input(26);
output(0, 228) <= input(27);
output(0, 229) <= input(28);
output(0, 230) <= input(29);
output(0, 231) <= input(30);
output(0, 232) <= input(31);
output(0, 233) <= input(33);
output(0, 234) <= input(35);
output(0, 235) <= input(38);
output(0, 236) <= input(39);
output(0, 237) <= input(41);
output(0, 238) <= input(43);
output(0, 239) <= input(45);
output(0, 240) <= input(24);
output(0, 241) <= input(25);
output(0, 242) <= input(26);
output(0, 243) <= input(27);
output(0, 244) <= input(28);
output(0, 245) <= input(29);
output(0, 246) <= input(30);
output(0, 247) <= input(31);
output(0, 248) <= input(33);
output(0, 249) <= input(35);
output(0, 250) <= input(38);
output(0, 251) <= input(39);
output(0, 252) <= input(41);
output(0, 253) <= input(43);
output(0, 254) <= input(45);
output(0, 255) <= input(46);
output(1, 0) <= input(0);
output(1, 1) <= input(1);
output(1, 2) <= input(2);
output(1, 3) <= input(3);
output(1, 4) <= input(4);
output(1, 5) <= input(5);
output(1, 6) <= input(6);
output(1, 7) <= input(7);
output(1, 8) <= input(8);
output(1, 9) <= input(9);
output(1, 10) <= input(10);
output(1, 11) <= input(11);
output(1, 12) <= input(12);
output(1, 13) <= input(13);
output(1, 14) <= input(14);
output(1, 15) <= input(15);
output(1, 16) <= input(16);
output(1, 17) <= input(17);
output(1, 18) <= input(18);
output(1, 19) <= input(19);
output(1, 20) <= input(20);
output(1, 21) <= input(21);
output(1, 22) <= input(22);
output(1, 23) <= input(23);
output(1, 24) <= input(24);
output(1, 25) <= input(25);
output(1, 26) <= input(26);
output(1, 27) <= input(27);
output(1, 28) <= input(28);
output(1, 29) <= input(29);
output(1, 30) <= input(30);
output(1, 31) <= input(31);
output(1, 32) <= input(1);
output(1, 33) <= input(2);
output(1, 34) <= input(3);
output(1, 35) <= input(4);
output(1, 36) <= input(5);
output(1, 37) <= input(6);
output(1, 38) <= input(7);
output(1, 39) <= input(8);
output(1, 40) <= input(9);
output(1, 41) <= input(10);
output(1, 42) <= input(11);
output(1, 43) <= input(12);
output(1, 44) <= input(13);
output(1, 45) <= input(14);
output(1, 46) <= input(15);
output(1, 47) <= input(32);
output(1, 48) <= input(2);
output(1, 49) <= input(3);
output(1, 50) <= input(4);
output(1, 51) <= input(5);
output(1, 52) <= input(6);
output(1, 53) <= input(7);
output(1, 54) <= input(8);
output(1, 55) <= input(9);
output(1, 56) <= input(10);
output(1, 57) <= input(11);
output(1, 58) <= input(12);
output(1, 59) <= input(13);
output(1, 60) <= input(14);
output(1, 61) <= input(15);
output(1, 62) <= input(32);
output(1, 63) <= input(34);
output(1, 64) <= input(18);
output(1, 65) <= input(19);
output(1, 66) <= input(20);
output(1, 67) <= input(21);
output(1, 68) <= input(22);
output(1, 69) <= input(23);
output(1, 70) <= input(24);
output(1, 71) <= input(25);
output(1, 72) <= input(26);
output(1, 73) <= input(27);
output(1, 74) <= input(28);
output(1, 75) <= input(29);
output(1, 76) <= input(30);
output(1, 77) <= input(31);
output(1, 78) <= input(33);
output(1, 79) <= input(35);
output(1, 80) <= input(3);
output(1, 81) <= input(4);
output(1, 82) <= input(5);
output(1, 83) <= input(6);
output(1, 84) <= input(7);
output(1, 85) <= input(8);
output(1, 86) <= input(9);
output(1, 87) <= input(10);
output(1, 88) <= input(11);
output(1, 89) <= input(12);
output(1, 90) <= input(13);
output(1, 91) <= input(14);
output(1, 92) <= input(15);
output(1, 93) <= input(32);
output(1, 94) <= input(34);
output(1, 95) <= input(36);
output(1, 96) <= input(19);
output(1, 97) <= input(20);
output(1, 98) <= input(21);
output(1, 99) <= input(22);
output(1, 100) <= input(23);
output(1, 101) <= input(24);
output(1, 102) <= input(25);
output(1, 103) <= input(26);
output(1, 104) <= input(27);
output(1, 105) <= input(28);
output(1, 106) <= input(29);
output(1, 107) <= input(30);
output(1, 108) <= input(31);
output(1, 109) <= input(33);
output(1, 110) <= input(35);
output(1, 111) <= input(38);
output(1, 112) <= input(20);
output(1, 113) <= input(21);
output(1, 114) <= input(22);
output(1, 115) <= input(23);
output(1, 116) <= input(24);
output(1, 117) <= input(25);
output(1, 118) <= input(26);
output(1, 119) <= input(27);
output(1, 120) <= input(28);
output(1, 121) <= input(29);
output(1, 122) <= input(30);
output(1, 123) <= input(31);
output(1, 124) <= input(33);
output(1, 125) <= input(35);
output(1, 126) <= input(38);
output(1, 127) <= input(39);
output(1, 128) <= input(5);
output(1, 129) <= input(6);
output(1, 130) <= input(7);
output(1, 131) <= input(8);
output(1, 132) <= input(9);
output(1, 133) <= input(10);
output(1, 134) <= input(11);
output(1, 135) <= input(12);
output(1, 136) <= input(13);
output(1, 137) <= input(14);
output(1, 138) <= input(15);
output(1, 139) <= input(32);
output(1, 140) <= input(34);
output(1, 141) <= input(36);
output(1, 142) <= input(37);
output(1, 143) <= input(40);
output(1, 144) <= input(21);
output(1, 145) <= input(22);
output(1, 146) <= input(23);
output(1, 147) <= input(24);
output(1, 148) <= input(25);
output(1, 149) <= input(26);
output(1, 150) <= input(27);
output(1, 151) <= input(28);
output(1, 152) <= input(29);
output(1, 153) <= input(30);
output(1, 154) <= input(31);
output(1, 155) <= input(33);
output(1, 156) <= input(35);
output(1, 157) <= input(38);
output(1, 158) <= input(39);
output(1, 159) <= input(41);
output(1, 160) <= input(6);
output(1, 161) <= input(7);
output(1, 162) <= input(8);
output(1, 163) <= input(9);
output(1, 164) <= input(10);
output(1, 165) <= input(11);
output(1, 166) <= input(12);
output(1, 167) <= input(13);
output(1, 168) <= input(14);
output(1, 169) <= input(15);
output(1, 170) <= input(32);
output(1, 171) <= input(34);
output(1, 172) <= input(36);
output(1, 173) <= input(37);
output(1, 174) <= input(40);
output(1, 175) <= input(42);
output(1, 176) <= input(7);
output(1, 177) <= input(8);
output(1, 178) <= input(9);
output(1, 179) <= input(10);
output(1, 180) <= input(11);
output(1, 181) <= input(12);
output(1, 182) <= input(13);
output(1, 183) <= input(14);
output(1, 184) <= input(15);
output(1, 185) <= input(32);
output(1, 186) <= input(34);
output(1, 187) <= input(36);
output(1, 188) <= input(37);
output(1, 189) <= input(40);
output(1, 190) <= input(42);
output(1, 191) <= input(44);
output(1, 192) <= input(23);
output(1, 193) <= input(24);
output(1, 194) <= input(25);
output(1, 195) <= input(26);
output(1, 196) <= input(27);
output(1, 197) <= input(28);
output(1, 198) <= input(29);
output(1, 199) <= input(30);
output(1, 200) <= input(31);
output(1, 201) <= input(33);
output(1, 202) <= input(35);
output(1, 203) <= input(38);
output(1, 204) <= input(39);
output(1, 205) <= input(41);
output(1, 206) <= input(43);
output(1, 207) <= input(45);
output(1, 208) <= input(8);
output(1, 209) <= input(9);
output(1, 210) <= input(10);
output(1, 211) <= input(11);
output(1, 212) <= input(12);
output(1, 213) <= input(13);
output(1, 214) <= input(14);
output(1, 215) <= input(15);
output(1, 216) <= input(32);
output(1, 217) <= input(34);
output(1, 218) <= input(36);
output(1, 219) <= input(37);
output(1, 220) <= input(40);
output(1, 221) <= input(42);
output(1, 222) <= input(44);
output(1, 223) <= input(47);
output(1, 224) <= input(24);
output(1, 225) <= input(25);
output(1, 226) <= input(26);
output(1, 227) <= input(27);
output(1, 228) <= input(28);
output(1, 229) <= input(29);
output(1, 230) <= input(30);
output(1, 231) <= input(31);
output(1, 232) <= input(33);
output(1, 233) <= input(35);
output(1, 234) <= input(38);
output(1, 235) <= input(39);
output(1, 236) <= input(41);
output(1, 237) <= input(43);
output(1, 238) <= input(45);
output(1, 239) <= input(46);
output(1, 240) <= input(25);
output(1, 241) <= input(26);
output(1, 242) <= input(27);
output(1, 243) <= input(28);
output(1, 244) <= input(29);
output(1, 245) <= input(30);
output(1, 246) <= input(31);
output(1, 247) <= input(33);
output(1, 248) <= input(35);
output(1, 249) <= input(38);
output(1, 250) <= input(39);
output(1, 251) <= input(41);
output(1, 252) <= input(43);
output(1, 253) <= input(45);
output(1, 254) <= input(46);
output(1, 255) <= input(48);
output(2, 0) <= input(0);
output(2, 1) <= input(1);
output(2, 2) <= input(2);
output(2, 3) <= input(3);
output(2, 4) <= input(4);
output(2, 5) <= input(5);
output(2, 6) <= input(6);
output(2, 7) <= input(7);
output(2, 8) <= input(8);
output(2, 9) <= input(9);
output(2, 10) <= input(10);
output(2, 11) <= input(11);
output(2, 12) <= input(12);
output(2, 13) <= input(13);
output(2, 14) <= input(14);
output(2, 15) <= input(15);
output(2, 16) <= input(16);
output(2, 17) <= input(17);
output(2, 18) <= input(18);
output(2, 19) <= input(19);
output(2, 20) <= input(20);
output(2, 21) <= input(21);
output(2, 22) <= input(22);
output(2, 23) <= input(23);
output(2, 24) <= input(24);
output(2, 25) <= input(25);
output(2, 26) <= input(26);
output(2, 27) <= input(27);
output(2, 28) <= input(28);
output(2, 29) <= input(29);
output(2, 30) <= input(30);
output(2, 31) <= input(31);
output(2, 32) <= input(17);
output(2, 33) <= input(18);
output(2, 34) <= input(19);
output(2, 35) <= input(20);
output(2, 36) <= input(21);
output(2, 37) <= input(22);
output(2, 38) <= input(23);
output(2, 39) <= input(24);
output(2, 40) <= input(25);
output(2, 41) <= input(26);
output(2, 42) <= input(27);
output(2, 43) <= input(28);
output(2, 44) <= input(29);
output(2, 45) <= input(30);
output(2, 46) <= input(31);
output(2, 47) <= input(33);
output(2, 48) <= input(2);
output(2, 49) <= input(3);
output(2, 50) <= input(4);
output(2, 51) <= input(5);
output(2, 52) <= input(6);
output(2, 53) <= input(7);
output(2, 54) <= input(8);
output(2, 55) <= input(9);
output(2, 56) <= input(10);
output(2, 57) <= input(11);
output(2, 58) <= input(12);
output(2, 59) <= input(13);
output(2, 60) <= input(14);
output(2, 61) <= input(15);
output(2, 62) <= input(32);
output(2, 63) <= input(34);
output(2, 64) <= input(3);
output(2, 65) <= input(4);
output(2, 66) <= input(5);
output(2, 67) <= input(6);
output(2, 68) <= input(7);
output(2, 69) <= input(8);
output(2, 70) <= input(9);
output(2, 71) <= input(10);
output(2, 72) <= input(11);
output(2, 73) <= input(12);
output(2, 74) <= input(13);
output(2, 75) <= input(14);
output(2, 76) <= input(15);
output(2, 77) <= input(32);
output(2, 78) <= input(34);
output(2, 79) <= input(36);
output(2, 80) <= input(19);
output(2, 81) <= input(20);
output(2, 82) <= input(21);
output(2, 83) <= input(22);
output(2, 84) <= input(23);
output(2, 85) <= input(24);
output(2, 86) <= input(25);
output(2, 87) <= input(26);
output(2, 88) <= input(27);
output(2, 89) <= input(28);
output(2, 90) <= input(29);
output(2, 91) <= input(30);
output(2, 92) <= input(31);
output(2, 93) <= input(33);
output(2, 94) <= input(35);
output(2, 95) <= input(38);
output(2, 96) <= input(20);
output(2, 97) <= input(21);
output(2, 98) <= input(22);
output(2, 99) <= input(23);
output(2, 100) <= input(24);
output(2, 101) <= input(25);
output(2, 102) <= input(26);
output(2, 103) <= input(27);
output(2, 104) <= input(28);
output(2, 105) <= input(29);
output(2, 106) <= input(30);
output(2, 107) <= input(31);
output(2, 108) <= input(33);
output(2, 109) <= input(35);
output(2, 110) <= input(38);
output(2, 111) <= input(39);
output(2, 112) <= input(5);
output(2, 113) <= input(6);
output(2, 114) <= input(7);
output(2, 115) <= input(8);
output(2, 116) <= input(9);
output(2, 117) <= input(10);
output(2, 118) <= input(11);
output(2, 119) <= input(12);
output(2, 120) <= input(13);
output(2, 121) <= input(14);
output(2, 122) <= input(15);
output(2, 123) <= input(32);
output(2, 124) <= input(34);
output(2, 125) <= input(36);
output(2, 126) <= input(37);
output(2, 127) <= input(40);
output(2, 128) <= input(21);
output(2, 129) <= input(22);
output(2, 130) <= input(23);
output(2, 131) <= input(24);
output(2, 132) <= input(25);
output(2, 133) <= input(26);
output(2, 134) <= input(27);
output(2, 135) <= input(28);
output(2, 136) <= input(29);
output(2, 137) <= input(30);
output(2, 138) <= input(31);
output(2, 139) <= input(33);
output(2, 140) <= input(35);
output(2, 141) <= input(38);
output(2, 142) <= input(39);
output(2, 143) <= input(41);
output(2, 144) <= input(22);
output(2, 145) <= input(23);
output(2, 146) <= input(24);
output(2, 147) <= input(25);
output(2, 148) <= input(26);
output(2, 149) <= input(27);
output(2, 150) <= input(28);
output(2, 151) <= input(29);
output(2, 152) <= input(30);
output(2, 153) <= input(31);
output(2, 154) <= input(33);
output(2, 155) <= input(35);
output(2, 156) <= input(38);
output(2, 157) <= input(39);
output(2, 158) <= input(41);
output(2, 159) <= input(43);
output(2, 160) <= input(7);
output(2, 161) <= input(8);
output(2, 162) <= input(9);
output(2, 163) <= input(10);
output(2, 164) <= input(11);
output(2, 165) <= input(12);
output(2, 166) <= input(13);
output(2, 167) <= input(14);
output(2, 168) <= input(15);
output(2, 169) <= input(32);
output(2, 170) <= input(34);
output(2, 171) <= input(36);
output(2, 172) <= input(37);
output(2, 173) <= input(40);
output(2, 174) <= input(42);
output(2, 175) <= input(44);
output(2, 176) <= input(8);
output(2, 177) <= input(9);
output(2, 178) <= input(10);
output(2, 179) <= input(11);
output(2, 180) <= input(12);
output(2, 181) <= input(13);
output(2, 182) <= input(14);
output(2, 183) <= input(15);
output(2, 184) <= input(32);
output(2, 185) <= input(34);
output(2, 186) <= input(36);
output(2, 187) <= input(37);
output(2, 188) <= input(40);
output(2, 189) <= input(42);
output(2, 190) <= input(44);
output(2, 191) <= input(47);
output(2, 192) <= input(24);
output(2, 193) <= input(25);
output(2, 194) <= input(26);
output(2, 195) <= input(27);
output(2, 196) <= input(28);
output(2, 197) <= input(29);
output(2, 198) <= input(30);
output(2, 199) <= input(31);
output(2, 200) <= input(33);
output(2, 201) <= input(35);
output(2, 202) <= input(38);
output(2, 203) <= input(39);
output(2, 204) <= input(41);
output(2, 205) <= input(43);
output(2, 206) <= input(45);
output(2, 207) <= input(46);
output(2, 208) <= input(25);
output(2, 209) <= input(26);
output(2, 210) <= input(27);
output(2, 211) <= input(28);
output(2, 212) <= input(29);
output(2, 213) <= input(30);
output(2, 214) <= input(31);
output(2, 215) <= input(33);
output(2, 216) <= input(35);
output(2, 217) <= input(38);
output(2, 218) <= input(39);
output(2, 219) <= input(41);
output(2, 220) <= input(43);
output(2, 221) <= input(45);
output(2, 222) <= input(46);
output(2, 223) <= input(48);
output(2, 224) <= input(10);
output(2, 225) <= input(11);
output(2, 226) <= input(12);
output(2, 227) <= input(13);
output(2, 228) <= input(14);
output(2, 229) <= input(15);
output(2, 230) <= input(32);
output(2, 231) <= input(34);
output(2, 232) <= input(36);
output(2, 233) <= input(37);
output(2, 234) <= input(40);
output(2, 235) <= input(42);
output(2, 236) <= input(44);
output(2, 237) <= input(47);
output(2, 238) <= input(49);
output(2, 239) <= input(50);
output(2, 240) <= input(11);
output(2, 241) <= input(12);
output(2, 242) <= input(13);
output(2, 243) <= input(14);
output(2, 244) <= input(15);
output(2, 245) <= input(32);
output(2, 246) <= input(34);
output(2, 247) <= input(36);
output(2, 248) <= input(37);
output(2, 249) <= input(40);
output(2, 250) <= input(42);
output(2, 251) <= input(44);
output(2, 252) <= input(47);
output(2, 253) <= input(49);
output(2, 254) <= input(50);
output(2, 255) <= input(51);
output(3, 0) <= input(0);
output(3, 1) <= input(1);
output(3, 2) <= input(2);
output(3, 3) <= input(3);
output(3, 4) <= input(4);
output(3, 5) <= input(5);
output(3, 6) <= input(6);
output(3, 7) <= input(7);
output(3, 8) <= input(8);
output(3, 9) <= input(9);
output(3, 10) <= input(10);
output(3, 11) <= input(11);
output(3, 12) <= input(12);
output(3, 13) <= input(13);
output(3, 14) <= input(14);
output(3, 15) <= input(15);
output(3, 16) <= input(1);
output(3, 17) <= input(2);
output(3, 18) <= input(3);
output(3, 19) <= input(4);
output(3, 20) <= input(5);
output(3, 21) <= input(6);
output(3, 22) <= input(7);
output(3, 23) <= input(8);
output(3, 24) <= input(9);
output(3, 25) <= input(10);
output(3, 26) <= input(11);
output(3, 27) <= input(12);
output(3, 28) <= input(13);
output(3, 29) <= input(14);
output(3, 30) <= input(15);
output(3, 31) <= input(32);
output(3, 32) <= input(17);
output(3, 33) <= input(18);
output(3, 34) <= input(19);
output(3, 35) <= input(20);
output(3, 36) <= input(21);
output(3, 37) <= input(22);
output(3, 38) <= input(23);
output(3, 39) <= input(24);
output(3, 40) <= input(25);
output(3, 41) <= input(26);
output(3, 42) <= input(27);
output(3, 43) <= input(28);
output(3, 44) <= input(29);
output(3, 45) <= input(30);
output(3, 46) <= input(31);
output(3, 47) <= input(33);
output(3, 48) <= input(18);
output(3, 49) <= input(19);
output(3, 50) <= input(20);
output(3, 51) <= input(21);
output(3, 52) <= input(22);
output(3, 53) <= input(23);
output(3, 54) <= input(24);
output(3, 55) <= input(25);
output(3, 56) <= input(26);
output(3, 57) <= input(27);
output(3, 58) <= input(28);
output(3, 59) <= input(29);
output(3, 60) <= input(30);
output(3, 61) <= input(31);
output(3, 62) <= input(33);
output(3, 63) <= input(35);
output(3, 64) <= input(19);
output(3, 65) <= input(20);
output(3, 66) <= input(21);
output(3, 67) <= input(22);
output(3, 68) <= input(23);
output(3, 69) <= input(24);
output(3, 70) <= input(25);
output(3, 71) <= input(26);
output(3, 72) <= input(27);
output(3, 73) <= input(28);
output(3, 74) <= input(29);
output(3, 75) <= input(30);
output(3, 76) <= input(31);
output(3, 77) <= input(33);
output(3, 78) <= input(35);
output(3, 79) <= input(38);
output(3, 80) <= input(4);
output(3, 81) <= input(5);
output(3, 82) <= input(6);
output(3, 83) <= input(7);
output(3, 84) <= input(8);
output(3, 85) <= input(9);
output(3, 86) <= input(10);
output(3, 87) <= input(11);
output(3, 88) <= input(12);
output(3, 89) <= input(13);
output(3, 90) <= input(14);
output(3, 91) <= input(15);
output(3, 92) <= input(32);
output(3, 93) <= input(34);
output(3, 94) <= input(36);
output(3, 95) <= input(37);
output(3, 96) <= input(5);
output(3, 97) <= input(6);
output(3, 98) <= input(7);
output(3, 99) <= input(8);
output(3, 100) <= input(9);
output(3, 101) <= input(10);
output(3, 102) <= input(11);
output(3, 103) <= input(12);
output(3, 104) <= input(13);
output(3, 105) <= input(14);
output(3, 106) <= input(15);
output(3, 107) <= input(32);
output(3, 108) <= input(34);
output(3, 109) <= input(36);
output(3, 110) <= input(37);
output(3, 111) <= input(40);
output(3, 112) <= input(6);
output(3, 113) <= input(7);
output(3, 114) <= input(8);
output(3, 115) <= input(9);
output(3, 116) <= input(10);
output(3, 117) <= input(11);
output(3, 118) <= input(12);
output(3, 119) <= input(13);
output(3, 120) <= input(14);
output(3, 121) <= input(15);
output(3, 122) <= input(32);
output(3, 123) <= input(34);
output(3, 124) <= input(36);
output(3, 125) <= input(37);
output(3, 126) <= input(40);
output(3, 127) <= input(42);
output(3, 128) <= input(22);
output(3, 129) <= input(23);
output(3, 130) <= input(24);
output(3, 131) <= input(25);
output(3, 132) <= input(26);
output(3, 133) <= input(27);
output(3, 134) <= input(28);
output(3, 135) <= input(29);
output(3, 136) <= input(30);
output(3, 137) <= input(31);
output(3, 138) <= input(33);
output(3, 139) <= input(35);
output(3, 140) <= input(38);
output(3, 141) <= input(39);
output(3, 142) <= input(41);
output(3, 143) <= input(43);
output(3, 144) <= input(23);
output(3, 145) <= input(24);
output(3, 146) <= input(25);
output(3, 147) <= input(26);
output(3, 148) <= input(27);
output(3, 149) <= input(28);
output(3, 150) <= input(29);
output(3, 151) <= input(30);
output(3, 152) <= input(31);
output(3, 153) <= input(33);
output(3, 154) <= input(35);
output(3, 155) <= input(38);
output(3, 156) <= input(39);
output(3, 157) <= input(41);
output(3, 158) <= input(43);
output(3, 159) <= input(45);
output(3, 160) <= input(8);
output(3, 161) <= input(9);
output(3, 162) <= input(10);
output(3, 163) <= input(11);
output(3, 164) <= input(12);
output(3, 165) <= input(13);
output(3, 166) <= input(14);
output(3, 167) <= input(15);
output(3, 168) <= input(32);
output(3, 169) <= input(34);
output(3, 170) <= input(36);
output(3, 171) <= input(37);
output(3, 172) <= input(40);
output(3, 173) <= input(42);
output(3, 174) <= input(44);
output(3, 175) <= input(47);
output(3, 176) <= input(9);
output(3, 177) <= input(10);
output(3, 178) <= input(11);
output(3, 179) <= input(12);
output(3, 180) <= input(13);
output(3, 181) <= input(14);
output(3, 182) <= input(15);
output(3, 183) <= input(32);
output(3, 184) <= input(34);
output(3, 185) <= input(36);
output(3, 186) <= input(37);
output(3, 187) <= input(40);
output(3, 188) <= input(42);
output(3, 189) <= input(44);
output(3, 190) <= input(47);
output(3, 191) <= input(49);
output(3, 192) <= input(10);
output(3, 193) <= input(11);
output(3, 194) <= input(12);
output(3, 195) <= input(13);
output(3, 196) <= input(14);
output(3, 197) <= input(15);
output(3, 198) <= input(32);
output(3, 199) <= input(34);
output(3, 200) <= input(36);
output(3, 201) <= input(37);
output(3, 202) <= input(40);
output(3, 203) <= input(42);
output(3, 204) <= input(44);
output(3, 205) <= input(47);
output(3, 206) <= input(49);
output(3, 207) <= input(50);
output(3, 208) <= input(26);
output(3, 209) <= input(27);
output(3, 210) <= input(28);
output(3, 211) <= input(29);
output(3, 212) <= input(30);
output(3, 213) <= input(31);
output(3, 214) <= input(33);
output(3, 215) <= input(35);
output(3, 216) <= input(38);
output(3, 217) <= input(39);
output(3, 218) <= input(41);
output(3, 219) <= input(43);
output(3, 220) <= input(45);
output(3, 221) <= input(46);
output(3, 222) <= input(48);
output(3, 223) <= input(52);
output(3, 224) <= input(27);
output(3, 225) <= input(28);
output(3, 226) <= input(29);
output(3, 227) <= input(30);
output(3, 228) <= input(31);
output(3, 229) <= input(33);
output(3, 230) <= input(35);
output(3, 231) <= input(38);
output(3, 232) <= input(39);
output(3, 233) <= input(41);
output(3, 234) <= input(43);
output(3, 235) <= input(45);
output(3, 236) <= input(46);
output(3, 237) <= input(48);
output(3, 238) <= input(52);
output(3, 239) <= input(53);
output(3, 240) <= input(28);
output(3, 241) <= input(29);
output(3, 242) <= input(30);
output(3, 243) <= input(31);
output(3, 244) <= input(33);
output(3, 245) <= input(35);
output(3, 246) <= input(38);
output(3, 247) <= input(39);
output(3, 248) <= input(41);
output(3, 249) <= input(43);
output(3, 250) <= input(45);
output(3, 251) <= input(46);
output(3, 252) <= input(48);
output(3, 253) <= input(52);
output(3, 254) <= input(53);
output(3, 255) <= input(54);
output(4, 0) <= input(0);
output(4, 1) <= input(1);
output(4, 2) <= input(2);
output(4, 3) <= input(3);
output(4, 4) <= input(4);
output(4, 5) <= input(5);
output(4, 6) <= input(6);
output(4, 7) <= input(7);
output(4, 8) <= input(8);
output(4, 9) <= input(9);
output(4, 10) <= input(10);
output(4, 11) <= input(11);
output(4, 12) <= input(12);
output(4, 13) <= input(13);
output(4, 14) <= input(14);
output(4, 15) <= input(15);
output(4, 16) <= input(1);
output(4, 17) <= input(2);
output(4, 18) <= input(3);
output(4, 19) <= input(4);
output(4, 20) <= input(5);
output(4, 21) <= input(6);
output(4, 22) <= input(7);
output(4, 23) <= input(8);
output(4, 24) <= input(9);
output(4, 25) <= input(10);
output(4, 26) <= input(11);
output(4, 27) <= input(12);
output(4, 28) <= input(13);
output(4, 29) <= input(14);
output(4, 30) <= input(15);
output(4, 31) <= input(32);
output(4, 32) <= input(2);
output(4, 33) <= input(3);
output(4, 34) <= input(4);
output(4, 35) <= input(5);
output(4, 36) <= input(6);
output(4, 37) <= input(7);
output(4, 38) <= input(8);
output(4, 39) <= input(9);
output(4, 40) <= input(10);
output(4, 41) <= input(11);
output(4, 42) <= input(12);
output(4, 43) <= input(13);
output(4, 44) <= input(14);
output(4, 45) <= input(15);
output(4, 46) <= input(32);
output(4, 47) <= input(34);
output(4, 48) <= input(3);
output(4, 49) <= input(4);
output(4, 50) <= input(5);
output(4, 51) <= input(6);
output(4, 52) <= input(7);
output(4, 53) <= input(8);
output(4, 54) <= input(9);
output(4, 55) <= input(10);
output(4, 56) <= input(11);
output(4, 57) <= input(12);
output(4, 58) <= input(13);
output(4, 59) <= input(14);
output(4, 60) <= input(15);
output(4, 61) <= input(32);
output(4, 62) <= input(34);
output(4, 63) <= input(36);
output(4, 64) <= input(4);
output(4, 65) <= input(5);
output(4, 66) <= input(6);
output(4, 67) <= input(7);
output(4, 68) <= input(8);
output(4, 69) <= input(9);
output(4, 70) <= input(10);
output(4, 71) <= input(11);
output(4, 72) <= input(12);
output(4, 73) <= input(13);
output(4, 74) <= input(14);
output(4, 75) <= input(15);
output(4, 76) <= input(32);
output(4, 77) <= input(34);
output(4, 78) <= input(36);
output(4, 79) <= input(37);
output(4, 80) <= input(20);
output(4, 81) <= input(21);
output(4, 82) <= input(22);
output(4, 83) <= input(23);
output(4, 84) <= input(24);
output(4, 85) <= input(25);
output(4, 86) <= input(26);
output(4, 87) <= input(27);
output(4, 88) <= input(28);
output(4, 89) <= input(29);
output(4, 90) <= input(30);
output(4, 91) <= input(31);
output(4, 92) <= input(33);
output(4, 93) <= input(35);
output(4, 94) <= input(38);
output(4, 95) <= input(39);
output(4, 96) <= input(21);
output(4, 97) <= input(22);
output(4, 98) <= input(23);
output(4, 99) <= input(24);
output(4, 100) <= input(25);
output(4, 101) <= input(26);
output(4, 102) <= input(27);
output(4, 103) <= input(28);
output(4, 104) <= input(29);
output(4, 105) <= input(30);
output(4, 106) <= input(31);
output(4, 107) <= input(33);
output(4, 108) <= input(35);
output(4, 109) <= input(38);
output(4, 110) <= input(39);
output(4, 111) <= input(41);
output(4, 112) <= input(22);
output(4, 113) <= input(23);
output(4, 114) <= input(24);
output(4, 115) <= input(25);
output(4, 116) <= input(26);
output(4, 117) <= input(27);
output(4, 118) <= input(28);
output(4, 119) <= input(29);
output(4, 120) <= input(30);
output(4, 121) <= input(31);
output(4, 122) <= input(33);
output(4, 123) <= input(35);
output(4, 124) <= input(38);
output(4, 125) <= input(39);
output(4, 126) <= input(41);
output(4, 127) <= input(43);
output(4, 128) <= input(23);
output(4, 129) <= input(24);
output(4, 130) <= input(25);
output(4, 131) <= input(26);
output(4, 132) <= input(27);
output(4, 133) <= input(28);
output(4, 134) <= input(29);
output(4, 135) <= input(30);
output(4, 136) <= input(31);
output(4, 137) <= input(33);
output(4, 138) <= input(35);
output(4, 139) <= input(38);
output(4, 140) <= input(39);
output(4, 141) <= input(41);
output(4, 142) <= input(43);
output(4, 143) <= input(45);
output(4, 144) <= input(24);
output(4, 145) <= input(25);
output(4, 146) <= input(26);
output(4, 147) <= input(27);
output(4, 148) <= input(28);
output(4, 149) <= input(29);
output(4, 150) <= input(30);
output(4, 151) <= input(31);
output(4, 152) <= input(33);
output(4, 153) <= input(35);
output(4, 154) <= input(38);
output(4, 155) <= input(39);
output(4, 156) <= input(41);
output(4, 157) <= input(43);
output(4, 158) <= input(45);
output(4, 159) <= input(46);
output(4, 160) <= input(9);
output(4, 161) <= input(10);
output(4, 162) <= input(11);
output(4, 163) <= input(12);
output(4, 164) <= input(13);
output(4, 165) <= input(14);
output(4, 166) <= input(15);
output(4, 167) <= input(32);
output(4, 168) <= input(34);
output(4, 169) <= input(36);
output(4, 170) <= input(37);
output(4, 171) <= input(40);
output(4, 172) <= input(42);
output(4, 173) <= input(44);
output(4, 174) <= input(47);
output(4, 175) <= input(49);
output(4, 176) <= input(10);
output(4, 177) <= input(11);
output(4, 178) <= input(12);
output(4, 179) <= input(13);
output(4, 180) <= input(14);
output(4, 181) <= input(15);
output(4, 182) <= input(32);
output(4, 183) <= input(34);
output(4, 184) <= input(36);
output(4, 185) <= input(37);
output(4, 186) <= input(40);
output(4, 187) <= input(42);
output(4, 188) <= input(44);
output(4, 189) <= input(47);
output(4, 190) <= input(49);
output(4, 191) <= input(50);
output(4, 192) <= input(11);
output(4, 193) <= input(12);
output(4, 194) <= input(13);
output(4, 195) <= input(14);
output(4, 196) <= input(15);
output(4, 197) <= input(32);
output(4, 198) <= input(34);
output(4, 199) <= input(36);
output(4, 200) <= input(37);
output(4, 201) <= input(40);
output(4, 202) <= input(42);
output(4, 203) <= input(44);
output(4, 204) <= input(47);
output(4, 205) <= input(49);
output(4, 206) <= input(50);
output(4, 207) <= input(51);
output(4, 208) <= input(12);
output(4, 209) <= input(13);
output(4, 210) <= input(14);
output(4, 211) <= input(15);
output(4, 212) <= input(32);
output(4, 213) <= input(34);
output(4, 214) <= input(36);
output(4, 215) <= input(37);
output(4, 216) <= input(40);
output(4, 217) <= input(42);
output(4, 218) <= input(44);
output(4, 219) <= input(47);
output(4, 220) <= input(49);
output(4, 221) <= input(50);
output(4, 222) <= input(51);
output(4, 223) <= input(55);
output(4, 224) <= input(13);
output(4, 225) <= input(14);
output(4, 226) <= input(15);
output(4, 227) <= input(32);
output(4, 228) <= input(34);
output(4, 229) <= input(36);
output(4, 230) <= input(37);
output(4, 231) <= input(40);
output(4, 232) <= input(42);
output(4, 233) <= input(44);
output(4, 234) <= input(47);
output(4, 235) <= input(49);
output(4, 236) <= input(50);
output(4, 237) <= input(51);
output(4, 238) <= input(55);
output(4, 239) <= input(56);
output(4, 240) <= input(14);
output(4, 241) <= input(15);
output(4, 242) <= input(32);
output(4, 243) <= input(34);
output(4, 244) <= input(36);
output(4, 245) <= input(37);
output(4, 246) <= input(40);
output(4, 247) <= input(42);
output(4, 248) <= input(44);
output(4, 249) <= input(47);
output(4, 250) <= input(49);
output(4, 251) <= input(50);
output(4, 252) <= input(51);
output(4, 253) <= input(55);
output(4, 254) <= input(56);
output(4, 255) <= input(57);
output(5, 0) <= input(16);
output(5, 1) <= input(17);
output(5, 2) <= input(18);
output(5, 3) <= input(19);
output(5, 4) <= input(20);
output(5, 5) <= input(21);
output(5, 6) <= input(22);
output(5, 7) <= input(23);
output(5, 8) <= input(24);
output(5, 9) <= input(25);
output(5, 10) <= input(26);
output(5, 11) <= input(27);
output(5, 12) <= input(28);
output(5, 13) <= input(29);
output(5, 14) <= input(30);
output(5, 15) <= input(31);
output(5, 16) <= input(17);
output(5, 17) <= input(18);
output(5, 18) <= input(19);
output(5, 19) <= input(20);
output(5, 20) <= input(21);
output(5, 21) <= input(22);
output(5, 22) <= input(23);
output(5, 23) <= input(24);
output(5, 24) <= input(25);
output(5, 25) <= input(26);
output(5, 26) <= input(27);
output(5, 27) <= input(28);
output(5, 28) <= input(29);
output(5, 29) <= input(30);
output(5, 30) <= input(31);
output(5, 31) <= input(33);
output(5, 32) <= input(18);
output(5, 33) <= input(19);
output(5, 34) <= input(20);
output(5, 35) <= input(21);
output(5, 36) <= input(22);
output(5, 37) <= input(23);
output(5, 38) <= input(24);
output(5, 39) <= input(25);
output(5, 40) <= input(26);
output(5, 41) <= input(27);
output(5, 42) <= input(28);
output(5, 43) <= input(29);
output(5, 44) <= input(30);
output(5, 45) <= input(31);
output(5, 46) <= input(33);
output(5, 47) <= input(35);
output(5, 48) <= input(19);
output(5, 49) <= input(20);
output(5, 50) <= input(21);
output(5, 51) <= input(22);
output(5, 52) <= input(23);
output(5, 53) <= input(24);
output(5, 54) <= input(25);
output(5, 55) <= input(26);
output(5, 56) <= input(27);
output(5, 57) <= input(28);
output(5, 58) <= input(29);
output(5, 59) <= input(30);
output(5, 60) <= input(31);
output(5, 61) <= input(33);
output(5, 62) <= input(35);
output(5, 63) <= input(38);
output(5, 64) <= input(20);
output(5, 65) <= input(21);
output(5, 66) <= input(22);
output(5, 67) <= input(23);
output(5, 68) <= input(24);
output(5, 69) <= input(25);
output(5, 70) <= input(26);
output(5, 71) <= input(27);
output(5, 72) <= input(28);
output(5, 73) <= input(29);
output(5, 74) <= input(30);
output(5, 75) <= input(31);
output(5, 76) <= input(33);
output(5, 77) <= input(35);
output(5, 78) <= input(38);
output(5, 79) <= input(39);
output(5, 80) <= input(21);
output(5, 81) <= input(22);
output(5, 82) <= input(23);
output(5, 83) <= input(24);
output(5, 84) <= input(25);
output(5, 85) <= input(26);
output(5, 86) <= input(27);
output(5, 87) <= input(28);
output(5, 88) <= input(29);
output(5, 89) <= input(30);
output(5, 90) <= input(31);
output(5, 91) <= input(33);
output(5, 92) <= input(35);
output(5, 93) <= input(38);
output(5, 94) <= input(39);
output(5, 95) <= input(41);
output(5, 96) <= input(22);
output(5, 97) <= input(23);
output(5, 98) <= input(24);
output(5, 99) <= input(25);
output(5, 100) <= input(26);
output(5, 101) <= input(27);
output(5, 102) <= input(28);
output(5, 103) <= input(29);
output(5, 104) <= input(30);
output(5, 105) <= input(31);
output(5, 106) <= input(33);
output(5, 107) <= input(35);
output(5, 108) <= input(38);
output(5, 109) <= input(39);
output(5, 110) <= input(41);
output(5, 111) <= input(43);
output(5, 112) <= input(23);
output(5, 113) <= input(24);
output(5, 114) <= input(25);
output(5, 115) <= input(26);
output(5, 116) <= input(27);
output(5, 117) <= input(28);
output(5, 118) <= input(29);
output(5, 119) <= input(30);
output(5, 120) <= input(31);
output(5, 121) <= input(33);
output(5, 122) <= input(35);
output(5, 123) <= input(38);
output(5, 124) <= input(39);
output(5, 125) <= input(41);
output(5, 126) <= input(43);
output(5, 127) <= input(45);
output(5, 128) <= input(24);
output(5, 129) <= input(25);
output(5, 130) <= input(26);
output(5, 131) <= input(27);
output(5, 132) <= input(28);
output(5, 133) <= input(29);
output(5, 134) <= input(30);
output(5, 135) <= input(31);
output(5, 136) <= input(33);
output(5, 137) <= input(35);
output(5, 138) <= input(38);
output(5, 139) <= input(39);
output(5, 140) <= input(41);
output(5, 141) <= input(43);
output(5, 142) <= input(45);
output(5, 143) <= input(46);
output(5, 144) <= input(25);
output(5, 145) <= input(26);
output(5, 146) <= input(27);
output(5, 147) <= input(28);
output(5, 148) <= input(29);
output(5, 149) <= input(30);
output(5, 150) <= input(31);
output(5, 151) <= input(33);
output(5, 152) <= input(35);
output(5, 153) <= input(38);
output(5, 154) <= input(39);
output(5, 155) <= input(41);
output(5, 156) <= input(43);
output(5, 157) <= input(45);
output(5, 158) <= input(46);
output(5, 159) <= input(48);
output(5, 160) <= input(26);
output(5, 161) <= input(27);
output(5, 162) <= input(28);
output(5, 163) <= input(29);
output(5, 164) <= input(30);
output(5, 165) <= input(31);
output(5, 166) <= input(33);
output(5, 167) <= input(35);
output(5, 168) <= input(38);
output(5, 169) <= input(39);
output(5, 170) <= input(41);
output(5, 171) <= input(43);
output(5, 172) <= input(45);
output(5, 173) <= input(46);
output(5, 174) <= input(48);
output(5, 175) <= input(52);
output(5, 176) <= input(27);
output(5, 177) <= input(28);
output(5, 178) <= input(29);
output(5, 179) <= input(30);
output(5, 180) <= input(31);
output(5, 181) <= input(33);
output(5, 182) <= input(35);
output(5, 183) <= input(38);
output(5, 184) <= input(39);
output(5, 185) <= input(41);
output(5, 186) <= input(43);
output(5, 187) <= input(45);
output(5, 188) <= input(46);
output(5, 189) <= input(48);
output(5, 190) <= input(52);
output(5, 191) <= input(53);
output(5, 192) <= input(28);
output(5, 193) <= input(29);
output(5, 194) <= input(30);
output(5, 195) <= input(31);
output(5, 196) <= input(33);
output(5, 197) <= input(35);
output(5, 198) <= input(38);
output(5, 199) <= input(39);
output(5, 200) <= input(41);
output(5, 201) <= input(43);
output(5, 202) <= input(45);
output(5, 203) <= input(46);
output(5, 204) <= input(48);
output(5, 205) <= input(52);
output(5, 206) <= input(53);
output(5, 207) <= input(54);
output(5, 208) <= input(29);
output(5, 209) <= input(30);
output(5, 210) <= input(31);
output(5, 211) <= input(33);
output(5, 212) <= input(35);
output(5, 213) <= input(38);
output(5, 214) <= input(39);
output(5, 215) <= input(41);
output(5, 216) <= input(43);
output(5, 217) <= input(45);
output(5, 218) <= input(46);
output(5, 219) <= input(48);
output(5, 220) <= input(52);
output(5, 221) <= input(53);
output(5, 222) <= input(54);
output(5, 223) <= input(58);
output(5, 224) <= input(30);
output(5, 225) <= input(31);
output(5, 226) <= input(33);
output(5, 227) <= input(35);
output(5, 228) <= input(38);
output(5, 229) <= input(39);
output(5, 230) <= input(41);
output(5, 231) <= input(43);
output(5, 232) <= input(45);
output(5, 233) <= input(46);
output(5, 234) <= input(48);
output(5, 235) <= input(52);
output(5, 236) <= input(53);
output(5, 237) <= input(54);
output(5, 238) <= input(58);
output(5, 239) <= input(59);
output(5, 240) <= input(31);
output(5, 241) <= input(33);
output(5, 242) <= input(35);
output(5, 243) <= input(38);
output(5, 244) <= input(39);
output(5, 245) <= input(41);
output(5, 246) <= input(43);
output(5, 247) <= input(45);
output(5, 248) <= input(46);
output(5, 249) <= input(48);
output(5, 250) <= input(52);
output(5, 251) <= input(53);
output(5, 252) <= input(54);
output(5, 253) <= input(58);
output(5, 254) <= input(59);
output(5, 255) <= input(60);
when others => for i in 0 to 7 loop for j in 0 to 255 loop output(i,j) <= "00000000"; end loop; end loop;
end case;
elsif control = "010" then 
case iteration_control is
when "0000" =>
output(0, 0) <= input(0);
output(0, 1) <= input(1);
output(0, 2) <= input(2);
output(0, 3) <= input(3);
output(0, 4) <= input(4);
output(0, 5) <= input(5);
output(0, 6) <= input(6);
output(0, 7) <= input(7);
output(0, 8) <= input(8);
output(0, 9) <= input(9);
output(0, 10) <= input(10);
output(0, 11) <= input(11);
output(0, 12) <= input(12);
output(0, 13) <= input(13);
output(0, 14) <= input(14);
output(0, 15) <= input(15);
output(0, 16) <= input(1);
output(0, 17) <= input(2);
output(0, 18) <= input(3);
output(0, 19) <= input(4);
output(0, 20) <= input(5);
output(0, 21) <= input(6);
output(0, 22) <= input(7);
output(0, 23) <= input(8);
output(0, 24) <= input(9);
output(0, 25) <= input(10);
output(0, 26) <= input(11);
output(0, 27) <= input(12);
output(0, 28) <= input(13);
output(0, 29) <= input(14);
output(0, 30) <= input(15);
output(0, 31) <= input(16);
output(0, 32) <= input(2);
output(0, 33) <= input(3);
output(0, 34) <= input(4);
output(0, 35) <= input(5);
output(0, 36) <= input(6);
output(0, 37) <= input(7);
output(0, 38) <= input(8);
output(0, 39) <= input(9);
output(0, 40) <= input(10);
output(0, 41) <= input(11);
output(0, 42) <= input(12);
output(0, 43) <= input(13);
output(0, 44) <= input(14);
output(0, 45) <= input(15);
output(0, 46) <= input(16);
output(0, 47) <= input(17);
output(0, 48) <= input(3);
output(0, 49) <= input(4);
output(0, 50) <= input(5);
output(0, 51) <= input(6);
output(0, 52) <= input(7);
output(0, 53) <= input(8);
output(0, 54) <= input(9);
output(0, 55) <= input(10);
output(0, 56) <= input(11);
output(0, 57) <= input(12);
output(0, 58) <= input(13);
output(0, 59) <= input(14);
output(0, 60) <= input(15);
output(0, 61) <= input(16);
output(0, 62) <= input(17);
output(0, 63) <= input(18);
output(0, 64) <= input(4);
output(0, 65) <= input(5);
output(0, 66) <= input(6);
output(0, 67) <= input(7);
output(0, 68) <= input(8);
output(0, 69) <= input(9);
output(0, 70) <= input(10);
output(0, 71) <= input(11);
output(0, 72) <= input(12);
output(0, 73) <= input(13);
output(0, 74) <= input(14);
output(0, 75) <= input(15);
output(0, 76) <= input(16);
output(0, 77) <= input(17);
output(0, 78) <= input(18);
output(0, 79) <= input(19);
output(0, 80) <= input(5);
output(0, 81) <= input(6);
output(0, 82) <= input(7);
output(0, 83) <= input(8);
output(0, 84) <= input(9);
output(0, 85) <= input(10);
output(0, 86) <= input(11);
output(0, 87) <= input(12);
output(0, 88) <= input(13);
output(0, 89) <= input(14);
output(0, 90) <= input(15);
output(0, 91) <= input(16);
output(0, 92) <= input(17);
output(0, 93) <= input(18);
output(0, 94) <= input(19);
output(0, 95) <= input(20);
output(0, 96) <= input(6);
output(0, 97) <= input(7);
output(0, 98) <= input(8);
output(0, 99) <= input(9);
output(0, 100) <= input(10);
output(0, 101) <= input(11);
output(0, 102) <= input(12);
output(0, 103) <= input(13);
output(0, 104) <= input(14);
output(0, 105) <= input(15);
output(0, 106) <= input(16);
output(0, 107) <= input(17);
output(0, 108) <= input(18);
output(0, 109) <= input(19);
output(0, 110) <= input(20);
output(0, 111) <= input(21);
output(0, 112) <= input(7);
output(0, 113) <= input(8);
output(0, 114) <= input(9);
output(0, 115) <= input(10);
output(0, 116) <= input(11);
output(0, 117) <= input(12);
output(0, 118) <= input(13);
output(0, 119) <= input(14);
output(0, 120) <= input(15);
output(0, 121) <= input(16);
output(0, 122) <= input(17);
output(0, 123) <= input(18);
output(0, 124) <= input(19);
output(0, 125) <= input(20);
output(0, 126) <= input(21);
output(0, 127) <= input(22);
output(0, 128) <= input(8);
output(0, 129) <= input(9);
output(0, 130) <= input(10);
output(0, 131) <= input(11);
output(0, 132) <= input(12);
output(0, 133) <= input(13);
output(0, 134) <= input(14);
output(0, 135) <= input(15);
output(0, 136) <= input(16);
output(0, 137) <= input(17);
output(0, 138) <= input(18);
output(0, 139) <= input(19);
output(0, 140) <= input(20);
output(0, 141) <= input(21);
output(0, 142) <= input(22);
output(0, 143) <= input(23);
output(0, 144) <= input(9);
output(0, 145) <= input(10);
output(0, 146) <= input(11);
output(0, 147) <= input(12);
output(0, 148) <= input(13);
output(0, 149) <= input(14);
output(0, 150) <= input(15);
output(0, 151) <= input(16);
output(0, 152) <= input(17);
output(0, 153) <= input(18);
output(0, 154) <= input(19);
output(0, 155) <= input(20);
output(0, 156) <= input(21);
output(0, 157) <= input(22);
output(0, 158) <= input(23);
output(0, 159) <= input(24);
output(0, 160) <= input(10);
output(0, 161) <= input(11);
output(0, 162) <= input(12);
output(0, 163) <= input(13);
output(0, 164) <= input(14);
output(0, 165) <= input(15);
output(0, 166) <= input(16);
output(0, 167) <= input(17);
output(0, 168) <= input(18);
output(0, 169) <= input(19);
output(0, 170) <= input(20);
output(0, 171) <= input(21);
output(0, 172) <= input(22);
output(0, 173) <= input(23);
output(0, 174) <= input(24);
output(0, 175) <= input(25);
output(0, 176) <= input(11);
output(0, 177) <= input(12);
output(0, 178) <= input(13);
output(0, 179) <= input(14);
output(0, 180) <= input(15);
output(0, 181) <= input(16);
output(0, 182) <= input(17);
output(0, 183) <= input(18);
output(0, 184) <= input(19);
output(0, 185) <= input(20);
output(0, 186) <= input(21);
output(0, 187) <= input(22);
output(0, 188) <= input(23);
output(0, 189) <= input(24);
output(0, 190) <= input(25);
output(0, 191) <= input(26);
output(0, 192) <= input(12);
output(0, 193) <= input(13);
output(0, 194) <= input(14);
output(0, 195) <= input(15);
output(0, 196) <= input(16);
output(0, 197) <= input(17);
output(0, 198) <= input(18);
output(0, 199) <= input(19);
output(0, 200) <= input(20);
output(0, 201) <= input(21);
output(0, 202) <= input(22);
output(0, 203) <= input(23);
output(0, 204) <= input(24);
output(0, 205) <= input(25);
output(0, 206) <= input(26);
output(0, 207) <= input(27);
output(0, 208) <= input(13);
output(0, 209) <= input(14);
output(0, 210) <= input(15);
output(0, 211) <= input(16);
output(0, 212) <= input(17);
output(0, 213) <= input(18);
output(0, 214) <= input(19);
output(0, 215) <= input(20);
output(0, 216) <= input(21);
output(0, 217) <= input(22);
output(0, 218) <= input(23);
output(0, 219) <= input(24);
output(0, 220) <= input(25);
output(0, 221) <= input(26);
output(0, 222) <= input(27);
output(0, 223) <= input(28);
output(0, 224) <= input(14);
output(0, 225) <= input(15);
output(0, 226) <= input(16);
output(0, 227) <= input(17);
output(0, 228) <= input(18);
output(0, 229) <= input(19);
output(0, 230) <= input(20);
output(0, 231) <= input(21);
output(0, 232) <= input(22);
output(0, 233) <= input(23);
output(0, 234) <= input(24);
output(0, 235) <= input(25);
output(0, 236) <= input(26);
output(0, 237) <= input(27);
output(0, 238) <= input(28);
output(0, 239) <= input(29);
output(0, 240) <= input(15);
output(0, 241) <= input(16);
output(0, 242) <= input(17);
output(0, 243) <= input(18);
output(0, 244) <= input(19);
output(0, 245) <= input(20);
output(0, 246) <= input(21);
output(0, 247) <= input(22);
output(0, 248) <= input(23);
output(0, 249) <= input(24);
output(0, 250) <= input(25);
output(0, 251) <= input(26);
output(0, 252) <= input(27);
output(0, 253) <= input(28);
output(0, 254) <= input(29);
output(0, 255) <= input(30);
output(1, 0) <= input(31);
output(1, 1) <= input(32);
output(1, 2) <= input(33);
output(1, 3) <= input(34);
output(1, 4) <= input(35);
output(1, 5) <= input(36);
output(1, 6) <= input(37);
output(1, 7) <= input(38);
output(1, 8) <= input(39);
output(1, 9) <= input(40);
output(1, 10) <= input(41);
output(1, 11) <= input(42);
output(1, 12) <= input(43);
output(1, 13) <= input(44);
output(1, 14) <= input(45);
output(1, 15) <= input(46);
output(1, 16) <= input(32);
output(1, 17) <= input(33);
output(1, 18) <= input(34);
output(1, 19) <= input(35);
output(1, 20) <= input(36);
output(1, 21) <= input(37);
output(1, 22) <= input(38);
output(1, 23) <= input(39);
output(1, 24) <= input(40);
output(1, 25) <= input(41);
output(1, 26) <= input(42);
output(1, 27) <= input(43);
output(1, 28) <= input(44);
output(1, 29) <= input(45);
output(1, 30) <= input(46);
output(1, 31) <= input(47);
output(1, 32) <= input(33);
output(1, 33) <= input(34);
output(1, 34) <= input(35);
output(1, 35) <= input(36);
output(1, 36) <= input(37);
output(1, 37) <= input(38);
output(1, 38) <= input(39);
output(1, 39) <= input(40);
output(1, 40) <= input(41);
output(1, 41) <= input(42);
output(1, 42) <= input(43);
output(1, 43) <= input(44);
output(1, 44) <= input(45);
output(1, 45) <= input(46);
output(1, 46) <= input(47);
output(1, 47) <= input(48);
output(1, 48) <= input(34);
output(1, 49) <= input(35);
output(1, 50) <= input(36);
output(1, 51) <= input(37);
output(1, 52) <= input(38);
output(1, 53) <= input(39);
output(1, 54) <= input(40);
output(1, 55) <= input(41);
output(1, 56) <= input(42);
output(1, 57) <= input(43);
output(1, 58) <= input(44);
output(1, 59) <= input(45);
output(1, 60) <= input(46);
output(1, 61) <= input(47);
output(1, 62) <= input(48);
output(1, 63) <= input(49);
output(1, 64) <= input(35);
output(1, 65) <= input(36);
output(1, 66) <= input(37);
output(1, 67) <= input(38);
output(1, 68) <= input(39);
output(1, 69) <= input(40);
output(1, 70) <= input(41);
output(1, 71) <= input(42);
output(1, 72) <= input(43);
output(1, 73) <= input(44);
output(1, 74) <= input(45);
output(1, 75) <= input(46);
output(1, 76) <= input(47);
output(1, 77) <= input(48);
output(1, 78) <= input(49);
output(1, 79) <= input(50);
output(1, 80) <= input(4);
output(1, 81) <= input(5);
output(1, 82) <= input(6);
output(1, 83) <= input(7);
output(1, 84) <= input(8);
output(1, 85) <= input(9);
output(1, 86) <= input(10);
output(1, 87) <= input(11);
output(1, 88) <= input(12);
output(1, 89) <= input(13);
output(1, 90) <= input(14);
output(1, 91) <= input(15);
output(1, 92) <= input(16);
output(1, 93) <= input(17);
output(1, 94) <= input(18);
output(1, 95) <= input(19);
output(1, 96) <= input(5);
output(1, 97) <= input(6);
output(1, 98) <= input(7);
output(1, 99) <= input(8);
output(1, 100) <= input(9);
output(1, 101) <= input(10);
output(1, 102) <= input(11);
output(1, 103) <= input(12);
output(1, 104) <= input(13);
output(1, 105) <= input(14);
output(1, 106) <= input(15);
output(1, 107) <= input(16);
output(1, 108) <= input(17);
output(1, 109) <= input(18);
output(1, 110) <= input(19);
output(1, 111) <= input(20);
output(1, 112) <= input(6);
output(1, 113) <= input(7);
output(1, 114) <= input(8);
output(1, 115) <= input(9);
output(1, 116) <= input(10);
output(1, 117) <= input(11);
output(1, 118) <= input(12);
output(1, 119) <= input(13);
output(1, 120) <= input(14);
output(1, 121) <= input(15);
output(1, 122) <= input(16);
output(1, 123) <= input(17);
output(1, 124) <= input(18);
output(1, 125) <= input(19);
output(1, 126) <= input(20);
output(1, 127) <= input(21);
output(1, 128) <= input(7);
output(1, 129) <= input(8);
output(1, 130) <= input(9);
output(1, 131) <= input(10);
output(1, 132) <= input(11);
output(1, 133) <= input(12);
output(1, 134) <= input(13);
output(1, 135) <= input(14);
output(1, 136) <= input(15);
output(1, 137) <= input(16);
output(1, 138) <= input(17);
output(1, 139) <= input(18);
output(1, 140) <= input(19);
output(1, 141) <= input(20);
output(1, 142) <= input(21);
output(1, 143) <= input(22);
output(1, 144) <= input(8);
output(1, 145) <= input(9);
output(1, 146) <= input(10);
output(1, 147) <= input(11);
output(1, 148) <= input(12);
output(1, 149) <= input(13);
output(1, 150) <= input(14);
output(1, 151) <= input(15);
output(1, 152) <= input(16);
output(1, 153) <= input(17);
output(1, 154) <= input(18);
output(1, 155) <= input(19);
output(1, 156) <= input(20);
output(1, 157) <= input(21);
output(1, 158) <= input(22);
output(1, 159) <= input(23);
output(1, 160) <= input(40);
output(1, 161) <= input(41);
output(1, 162) <= input(42);
output(1, 163) <= input(43);
output(1, 164) <= input(44);
output(1, 165) <= input(45);
output(1, 166) <= input(46);
output(1, 167) <= input(47);
output(1, 168) <= input(48);
output(1, 169) <= input(49);
output(1, 170) <= input(50);
output(1, 171) <= input(51);
output(1, 172) <= input(52);
output(1, 173) <= input(53);
output(1, 174) <= input(54);
output(1, 175) <= input(55);
output(1, 176) <= input(41);
output(1, 177) <= input(42);
output(1, 178) <= input(43);
output(1, 179) <= input(44);
output(1, 180) <= input(45);
output(1, 181) <= input(46);
output(1, 182) <= input(47);
output(1, 183) <= input(48);
output(1, 184) <= input(49);
output(1, 185) <= input(50);
output(1, 186) <= input(51);
output(1, 187) <= input(52);
output(1, 188) <= input(53);
output(1, 189) <= input(54);
output(1, 190) <= input(55);
output(1, 191) <= input(56);
output(1, 192) <= input(42);
output(1, 193) <= input(43);
output(1, 194) <= input(44);
output(1, 195) <= input(45);
output(1, 196) <= input(46);
output(1, 197) <= input(47);
output(1, 198) <= input(48);
output(1, 199) <= input(49);
output(1, 200) <= input(50);
output(1, 201) <= input(51);
output(1, 202) <= input(52);
output(1, 203) <= input(53);
output(1, 204) <= input(54);
output(1, 205) <= input(55);
output(1, 206) <= input(56);
output(1, 207) <= input(57);
output(1, 208) <= input(43);
output(1, 209) <= input(44);
output(1, 210) <= input(45);
output(1, 211) <= input(46);
output(1, 212) <= input(47);
output(1, 213) <= input(48);
output(1, 214) <= input(49);
output(1, 215) <= input(50);
output(1, 216) <= input(51);
output(1, 217) <= input(52);
output(1, 218) <= input(53);
output(1, 219) <= input(54);
output(1, 220) <= input(55);
output(1, 221) <= input(56);
output(1, 222) <= input(57);
output(1, 223) <= input(58);
output(1, 224) <= input(44);
output(1, 225) <= input(45);
output(1, 226) <= input(46);
output(1, 227) <= input(47);
output(1, 228) <= input(48);
output(1, 229) <= input(49);
output(1, 230) <= input(50);
output(1, 231) <= input(51);
output(1, 232) <= input(52);
output(1, 233) <= input(53);
output(1, 234) <= input(54);
output(1, 235) <= input(55);
output(1, 236) <= input(56);
output(1, 237) <= input(57);
output(1, 238) <= input(58);
output(1, 239) <= input(59);
output(1, 240) <= input(45);
output(1, 241) <= input(46);
output(1, 242) <= input(47);
output(1, 243) <= input(48);
output(1, 244) <= input(49);
output(1, 245) <= input(50);
output(1, 246) <= input(51);
output(1, 247) <= input(52);
output(1, 248) <= input(53);
output(1, 249) <= input(54);
output(1, 250) <= input(55);
output(1, 251) <= input(56);
output(1, 252) <= input(57);
output(1, 253) <= input(58);
output(1, 254) <= input(59);
output(1, 255) <= input(60);
output(2, 0) <= input(31);
output(2, 1) <= input(32);
output(2, 2) <= input(33);
output(2, 3) <= input(34);
output(2, 4) <= input(35);
output(2, 5) <= input(36);
output(2, 6) <= input(37);
output(2, 7) <= input(38);
output(2, 8) <= input(39);
output(2, 9) <= input(40);
output(2, 10) <= input(41);
output(2, 11) <= input(42);
output(2, 12) <= input(43);
output(2, 13) <= input(44);
output(2, 14) <= input(45);
output(2, 15) <= input(46);
output(2, 16) <= input(32);
output(2, 17) <= input(33);
output(2, 18) <= input(34);
output(2, 19) <= input(35);
output(2, 20) <= input(36);
output(2, 21) <= input(37);
output(2, 22) <= input(38);
output(2, 23) <= input(39);
output(2, 24) <= input(40);
output(2, 25) <= input(41);
output(2, 26) <= input(42);
output(2, 27) <= input(43);
output(2, 28) <= input(44);
output(2, 29) <= input(45);
output(2, 30) <= input(46);
output(2, 31) <= input(47);
output(2, 32) <= input(1);
output(2, 33) <= input(2);
output(2, 34) <= input(3);
output(2, 35) <= input(4);
output(2, 36) <= input(5);
output(2, 37) <= input(6);
output(2, 38) <= input(7);
output(2, 39) <= input(8);
output(2, 40) <= input(9);
output(2, 41) <= input(10);
output(2, 42) <= input(11);
output(2, 43) <= input(12);
output(2, 44) <= input(13);
output(2, 45) <= input(14);
output(2, 46) <= input(15);
output(2, 47) <= input(16);
output(2, 48) <= input(2);
output(2, 49) <= input(3);
output(2, 50) <= input(4);
output(2, 51) <= input(5);
output(2, 52) <= input(6);
output(2, 53) <= input(7);
output(2, 54) <= input(8);
output(2, 55) <= input(9);
output(2, 56) <= input(10);
output(2, 57) <= input(11);
output(2, 58) <= input(12);
output(2, 59) <= input(13);
output(2, 60) <= input(14);
output(2, 61) <= input(15);
output(2, 62) <= input(16);
output(2, 63) <= input(17);
output(2, 64) <= input(3);
output(2, 65) <= input(4);
output(2, 66) <= input(5);
output(2, 67) <= input(6);
output(2, 68) <= input(7);
output(2, 69) <= input(8);
output(2, 70) <= input(9);
output(2, 71) <= input(10);
output(2, 72) <= input(11);
output(2, 73) <= input(12);
output(2, 74) <= input(13);
output(2, 75) <= input(14);
output(2, 76) <= input(15);
output(2, 77) <= input(16);
output(2, 78) <= input(17);
output(2, 79) <= input(18);
output(2, 80) <= input(35);
output(2, 81) <= input(36);
output(2, 82) <= input(37);
output(2, 83) <= input(38);
output(2, 84) <= input(39);
output(2, 85) <= input(40);
output(2, 86) <= input(41);
output(2, 87) <= input(42);
output(2, 88) <= input(43);
output(2, 89) <= input(44);
output(2, 90) <= input(45);
output(2, 91) <= input(46);
output(2, 92) <= input(47);
output(2, 93) <= input(48);
output(2, 94) <= input(49);
output(2, 95) <= input(50);
output(2, 96) <= input(36);
output(2, 97) <= input(37);
output(2, 98) <= input(38);
output(2, 99) <= input(39);
output(2, 100) <= input(40);
output(2, 101) <= input(41);
output(2, 102) <= input(42);
output(2, 103) <= input(43);
output(2, 104) <= input(44);
output(2, 105) <= input(45);
output(2, 106) <= input(46);
output(2, 107) <= input(47);
output(2, 108) <= input(48);
output(2, 109) <= input(49);
output(2, 110) <= input(50);
output(2, 111) <= input(51);
output(2, 112) <= input(37);
output(2, 113) <= input(38);
output(2, 114) <= input(39);
output(2, 115) <= input(40);
output(2, 116) <= input(41);
output(2, 117) <= input(42);
output(2, 118) <= input(43);
output(2, 119) <= input(44);
output(2, 120) <= input(45);
output(2, 121) <= input(46);
output(2, 122) <= input(47);
output(2, 123) <= input(48);
output(2, 124) <= input(49);
output(2, 125) <= input(50);
output(2, 126) <= input(51);
output(2, 127) <= input(52);
output(2, 128) <= input(6);
output(2, 129) <= input(7);
output(2, 130) <= input(8);
output(2, 131) <= input(9);
output(2, 132) <= input(10);
output(2, 133) <= input(11);
output(2, 134) <= input(12);
output(2, 135) <= input(13);
output(2, 136) <= input(14);
output(2, 137) <= input(15);
output(2, 138) <= input(16);
output(2, 139) <= input(17);
output(2, 140) <= input(18);
output(2, 141) <= input(19);
output(2, 142) <= input(20);
output(2, 143) <= input(21);
output(2, 144) <= input(7);
output(2, 145) <= input(8);
output(2, 146) <= input(9);
output(2, 147) <= input(10);
output(2, 148) <= input(11);
output(2, 149) <= input(12);
output(2, 150) <= input(13);
output(2, 151) <= input(14);
output(2, 152) <= input(15);
output(2, 153) <= input(16);
output(2, 154) <= input(17);
output(2, 155) <= input(18);
output(2, 156) <= input(19);
output(2, 157) <= input(20);
output(2, 158) <= input(21);
output(2, 159) <= input(22);
output(2, 160) <= input(39);
output(2, 161) <= input(40);
output(2, 162) <= input(41);
output(2, 163) <= input(42);
output(2, 164) <= input(43);
output(2, 165) <= input(44);
output(2, 166) <= input(45);
output(2, 167) <= input(46);
output(2, 168) <= input(47);
output(2, 169) <= input(48);
output(2, 170) <= input(49);
output(2, 171) <= input(50);
output(2, 172) <= input(51);
output(2, 173) <= input(52);
output(2, 174) <= input(53);
output(2, 175) <= input(54);
output(2, 176) <= input(40);
output(2, 177) <= input(41);
output(2, 178) <= input(42);
output(2, 179) <= input(43);
output(2, 180) <= input(44);
output(2, 181) <= input(45);
output(2, 182) <= input(46);
output(2, 183) <= input(47);
output(2, 184) <= input(48);
output(2, 185) <= input(49);
output(2, 186) <= input(50);
output(2, 187) <= input(51);
output(2, 188) <= input(52);
output(2, 189) <= input(53);
output(2, 190) <= input(54);
output(2, 191) <= input(55);
output(2, 192) <= input(41);
output(2, 193) <= input(42);
output(2, 194) <= input(43);
output(2, 195) <= input(44);
output(2, 196) <= input(45);
output(2, 197) <= input(46);
output(2, 198) <= input(47);
output(2, 199) <= input(48);
output(2, 200) <= input(49);
output(2, 201) <= input(50);
output(2, 202) <= input(51);
output(2, 203) <= input(52);
output(2, 204) <= input(53);
output(2, 205) <= input(54);
output(2, 206) <= input(55);
output(2, 207) <= input(56);
output(2, 208) <= input(10);
output(2, 209) <= input(11);
output(2, 210) <= input(12);
output(2, 211) <= input(13);
output(2, 212) <= input(14);
output(2, 213) <= input(15);
output(2, 214) <= input(16);
output(2, 215) <= input(17);
output(2, 216) <= input(18);
output(2, 217) <= input(19);
output(2, 218) <= input(20);
output(2, 219) <= input(21);
output(2, 220) <= input(22);
output(2, 221) <= input(23);
output(2, 222) <= input(24);
output(2, 223) <= input(25);
output(2, 224) <= input(11);
output(2, 225) <= input(12);
output(2, 226) <= input(13);
output(2, 227) <= input(14);
output(2, 228) <= input(15);
output(2, 229) <= input(16);
output(2, 230) <= input(17);
output(2, 231) <= input(18);
output(2, 232) <= input(19);
output(2, 233) <= input(20);
output(2, 234) <= input(21);
output(2, 235) <= input(22);
output(2, 236) <= input(23);
output(2, 237) <= input(24);
output(2, 238) <= input(25);
output(2, 239) <= input(26);
output(2, 240) <= input(12);
output(2, 241) <= input(13);
output(2, 242) <= input(14);
output(2, 243) <= input(15);
output(2, 244) <= input(16);
output(2, 245) <= input(17);
output(2, 246) <= input(18);
output(2, 247) <= input(19);
output(2, 248) <= input(20);
output(2, 249) <= input(21);
output(2, 250) <= input(22);
output(2, 251) <= input(23);
output(2, 252) <= input(24);
output(2, 253) <= input(25);
output(2, 254) <= input(26);
output(2, 255) <= input(27);
output(3, 0) <= input(31);
output(3, 1) <= input(32);
output(3, 2) <= input(33);
output(3, 3) <= input(34);
output(3, 4) <= input(35);
output(3, 5) <= input(36);
output(3, 6) <= input(37);
output(3, 7) <= input(38);
output(3, 8) <= input(39);
output(3, 9) <= input(40);
output(3, 10) <= input(41);
output(3, 11) <= input(42);
output(3, 12) <= input(43);
output(3, 13) <= input(44);
output(3, 14) <= input(45);
output(3, 15) <= input(46);
output(3, 16) <= input(0);
output(3, 17) <= input(1);
output(3, 18) <= input(2);
output(3, 19) <= input(3);
output(3, 20) <= input(4);
output(3, 21) <= input(5);
output(3, 22) <= input(6);
output(3, 23) <= input(7);
output(3, 24) <= input(8);
output(3, 25) <= input(9);
output(3, 26) <= input(10);
output(3, 27) <= input(11);
output(3, 28) <= input(12);
output(3, 29) <= input(13);
output(3, 30) <= input(14);
output(3, 31) <= input(15);
output(3, 32) <= input(1);
output(3, 33) <= input(2);
output(3, 34) <= input(3);
output(3, 35) <= input(4);
output(3, 36) <= input(5);
output(3, 37) <= input(6);
output(3, 38) <= input(7);
output(3, 39) <= input(8);
output(3, 40) <= input(9);
output(3, 41) <= input(10);
output(3, 42) <= input(11);
output(3, 43) <= input(12);
output(3, 44) <= input(13);
output(3, 45) <= input(14);
output(3, 46) <= input(15);
output(3, 47) <= input(16);
output(3, 48) <= input(33);
output(3, 49) <= input(34);
output(3, 50) <= input(35);
output(3, 51) <= input(36);
output(3, 52) <= input(37);
output(3, 53) <= input(38);
output(3, 54) <= input(39);
output(3, 55) <= input(40);
output(3, 56) <= input(41);
output(3, 57) <= input(42);
output(3, 58) <= input(43);
output(3, 59) <= input(44);
output(3, 60) <= input(45);
output(3, 61) <= input(46);
output(3, 62) <= input(47);
output(3, 63) <= input(48);
output(3, 64) <= input(34);
output(3, 65) <= input(35);
output(3, 66) <= input(36);
output(3, 67) <= input(37);
output(3, 68) <= input(38);
output(3, 69) <= input(39);
output(3, 70) <= input(40);
output(3, 71) <= input(41);
output(3, 72) <= input(42);
output(3, 73) <= input(43);
output(3, 74) <= input(44);
output(3, 75) <= input(45);
output(3, 76) <= input(46);
output(3, 77) <= input(47);
output(3, 78) <= input(48);
output(3, 79) <= input(49);
output(3, 80) <= input(3);
output(3, 81) <= input(4);
output(3, 82) <= input(5);
output(3, 83) <= input(6);
output(3, 84) <= input(7);
output(3, 85) <= input(8);
output(3, 86) <= input(9);
output(3, 87) <= input(10);
output(3, 88) <= input(11);
output(3, 89) <= input(12);
output(3, 90) <= input(13);
output(3, 91) <= input(14);
output(3, 92) <= input(15);
output(3, 93) <= input(16);
output(3, 94) <= input(17);
output(3, 95) <= input(18);
output(3, 96) <= input(4);
output(3, 97) <= input(5);
output(3, 98) <= input(6);
output(3, 99) <= input(7);
output(3, 100) <= input(8);
output(3, 101) <= input(9);
output(3, 102) <= input(10);
output(3, 103) <= input(11);
output(3, 104) <= input(12);
output(3, 105) <= input(13);
output(3, 106) <= input(14);
output(3, 107) <= input(15);
output(3, 108) <= input(16);
output(3, 109) <= input(17);
output(3, 110) <= input(18);
output(3, 111) <= input(19);
output(3, 112) <= input(36);
output(3, 113) <= input(37);
output(3, 114) <= input(38);
output(3, 115) <= input(39);
output(3, 116) <= input(40);
output(3, 117) <= input(41);
output(3, 118) <= input(42);
output(3, 119) <= input(43);
output(3, 120) <= input(44);
output(3, 121) <= input(45);
output(3, 122) <= input(46);
output(3, 123) <= input(47);
output(3, 124) <= input(48);
output(3, 125) <= input(49);
output(3, 126) <= input(50);
output(3, 127) <= input(51);
output(3, 128) <= input(5);
output(3, 129) <= input(6);
output(3, 130) <= input(7);
output(3, 131) <= input(8);
output(3, 132) <= input(9);
output(3, 133) <= input(10);
output(3, 134) <= input(11);
output(3, 135) <= input(12);
output(3, 136) <= input(13);
output(3, 137) <= input(14);
output(3, 138) <= input(15);
output(3, 139) <= input(16);
output(3, 140) <= input(17);
output(3, 141) <= input(18);
output(3, 142) <= input(19);
output(3, 143) <= input(20);
output(3, 144) <= input(6);
output(3, 145) <= input(7);
output(3, 146) <= input(8);
output(3, 147) <= input(9);
output(3, 148) <= input(10);
output(3, 149) <= input(11);
output(3, 150) <= input(12);
output(3, 151) <= input(13);
output(3, 152) <= input(14);
output(3, 153) <= input(15);
output(3, 154) <= input(16);
output(3, 155) <= input(17);
output(3, 156) <= input(18);
output(3, 157) <= input(19);
output(3, 158) <= input(20);
output(3, 159) <= input(21);
output(3, 160) <= input(38);
output(3, 161) <= input(39);
output(3, 162) <= input(40);
output(3, 163) <= input(41);
output(3, 164) <= input(42);
output(3, 165) <= input(43);
output(3, 166) <= input(44);
output(3, 167) <= input(45);
output(3, 168) <= input(46);
output(3, 169) <= input(47);
output(3, 170) <= input(48);
output(3, 171) <= input(49);
output(3, 172) <= input(50);
output(3, 173) <= input(51);
output(3, 174) <= input(52);
output(3, 175) <= input(53);
output(3, 176) <= input(39);
output(3, 177) <= input(40);
output(3, 178) <= input(41);
output(3, 179) <= input(42);
output(3, 180) <= input(43);
output(3, 181) <= input(44);
output(3, 182) <= input(45);
output(3, 183) <= input(46);
output(3, 184) <= input(47);
output(3, 185) <= input(48);
output(3, 186) <= input(49);
output(3, 187) <= input(50);
output(3, 188) <= input(51);
output(3, 189) <= input(52);
output(3, 190) <= input(53);
output(3, 191) <= input(54);
output(3, 192) <= input(8);
output(3, 193) <= input(9);
output(3, 194) <= input(10);
output(3, 195) <= input(11);
output(3, 196) <= input(12);
output(3, 197) <= input(13);
output(3, 198) <= input(14);
output(3, 199) <= input(15);
output(3, 200) <= input(16);
output(3, 201) <= input(17);
output(3, 202) <= input(18);
output(3, 203) <= input(19);
output(3, 204) <= input(20);
output(3, 205) <= input(21);
output(3, 206) <= input(22);
output(3, 207) <= input(23);
output(3, 208) <= input(9);
output(3, 209) <= input(10);
output(3, 210) <= input(11);
output(3, 211) <= input(12);
output(3, 212) <= input(13);
output(3, 213) <= input(14);
output(3, 214) <= input(15);
output(3, 215) <= input(16);
output(3, 216) <= input(17);
output(3, 217) <= input(18);
output(3, 218) <= input(19);
output(3, 219) <= input(20);
output(3, 220) <= input(21);
output(3, 221) <= input(22);
output(3, 222) <= input(23);
output(3, 223) <= input(24);
output(3, 224) <= input(41);
output(3, 225) <= input(42);
output(3, 226) <= input(43);
output(3, 227) <= input(44);
output(3, 228) <= input(45);
output(3, 229) <= input(46);
output(3, 230) <= input(47);
output(3, 231) <= input(48);
output(3, 232) <= input(49);
output(3, 233) <= input(50);
output(3, 234) <= input(51);
output(3, 235) <= input(52);
output(3, 236) <= input(53);
output(3, 237) <= input(54);
output(3, 238) <= input(55);
output(3, 239) <= input(56);
output(3, 240) <= input(42);
output(3, 241) <= input(43);
output(3, 242) <= input(44);
output(3, 243) <= input(45);
output(3, 244) <= input(46);
output(3, 245) <= input(47);
output(3, 246) <= input(48);
output(3, 247) <= input(49);
output(3, 248) <= input(50);
output(3, 249) <= input(51);
output(3, 250) <= input(52);
output(3, 251) <= input(53);
output(3, 252) <= input(54);
output(3, 253) <= input(55);
output(3, 254) <= input(56);
output(3, 255) <= input(57);
output(4, 0) <= input(31);
output(4, 1) <= input(32);
output(4, 2) <= input(33);
output(4, 3) <= input(34);
output(4, 4) <= input(35);
output(4, 5) <= input(36);
output(4, 6) <= input(37);
output(4, 7) <= input(38);
output(4, 8) <= input(39);
output(4, 9) <= input(40);
output(4, 10) <= input(41);
output(4, 11) <= input(42);
output(4, 12) <= input(43);
output(4, 13) <= input(44);
output(4, 14) <= input(45);
output(4, 15) <= input(46);
output(4, 16) <= input(0);
output(4, 17) <= input(1);
output(4, 18) <= input(2);
output(4, 19) <= input(3);
output(4, 20) <= input(4);
output(4, 21) <= input(5);
output(4, 22) <= input(6);
output(4, 23) <= input(7);
output(4, 24) <= input(8);
output(4, 25) <= input(9);
output(4, 26) <= input(10);
output(4, 27) <= input(11);
output(4, 28) <= input(12);
output(4, 29) <= input(13);
output(4, 30) <= input(14);
output(4, 31) <= input(15);
output(4, 32) <= input(32);
output(4, 33) <= input(33);
output(4, 34) <= input(34);
output(4, 35) <= input(35);
output(4, 36) <= input(36);
output(4, 37) <= input(37);
output(4, 38) <= input(38);
output(4, 39) <= input(39);
output(4, 40) <= input(40);
output(4, 41) <= input(41);
output(4, 42) <= input(42);
output(4, 43) <= input(43);
output(4, 44) <= input(44);
output(4, 45) <= input(45);
output(4, 46) <= input(46);
output(4, 47) <= input(47);
output(4, 48) <= input(33);
output(4, 49) <= input(34);
output(4, 50) <= input(35);
output(4, 51) <= input(36);
output(4, 52) <= input(37);
output(4, 53) <= input(38);
output(4, 54) <= input(39);
output(4, 55) <= input(40);
output(4, 56) <= input(41);
output(4, 57) <= input(42);
output(4, 58) <= input(43);
output(4, 59) <= input(44);
output(4, 60) <= input(45);
output(4, 61) <= input(46);
output(4, 62) <= input(47);
output(4, 63) <= input(48);
output(4, 64) <= input(2);
output(4, 65) <= input(3);
output(4, 66) <= input(4);
output(4, 67) <= input(5);
output(4, 68) <= input(6);
output(4, 69) <= input(7);
output(4, 70) <= input(8);
output(4, 71) <= input(9);
output(4, 72) <= input(10);
output(4, 73) <= input(11);
output(4, 74) <= input(12);
output(4, 75) <= input(13);
output(4, 76) <= input(14);
output(4, 77) <= input(15);
output(4, 78) <= input(16);
output(4, 79) <= input(17);
output(4, 80) <= input(34);
output(4, 81) <= input(35);
output(4, 82) <= input(36);
output(4, 83) <= input(37);
output(4, 84) <= input(38);
output(4, 85) <= input(39);
output(4, 86) <= input(40);
output(4, 87) <= input(41);
output(4, 88) <= input(42);
output(4, 89) <= input(43);
output(4, 90) <= input(44);
output(4, 91) <= input(45);
output(4, 92) <= input(46);
output(4, 93) <= input(47);
output(4, 94) <= input(48);
output(4, 95) <= input(49);
output(4, 96) <= input(3);
output(4, 97) <= input(4);
output(4, 98) <= input(5);
output(4, 99) <= input(6);
output(4, 100) <= input(7);
output(4, 101) <= input(8);
output(4, 102) <= input(9);
output(4, 103) <= input(10);
output(4, 104) <= input(11);
output(4, 105) <= input(12);
output(4, 106) <= input(13);
output(4, 107) <= input(14);
output(4, 108) <= input(15);
output(4, 109) <= input(16);
output(4, 110) <= input(17);
output(4, 111) <= input(18);
output(4, 112) <= input(4);
output(4, 113) <= input(5);
output(4, 114) <= input(6);
output(4, 115) <= input(7);
output(4, 116) <= input(8);
output(4, 117) <= input(9);
output(4, 118) <= input(10);
output(4, 119) <= input(11);
output(4, 120) <= input(12);
output(4, 121) <= input(13);
output(4, 122) <= input(14);
output(4, 123) <= input(15);
output(4, 124) <= input(16);
output(4, 125) <= input(17);
output(4, 126) <= input(18);
output(4, 127) <= input(19);
output(4, 128) <= input(36);
output(4, 129) <= input(37);
output(4, 130) <= input(38);
output(4, 131) <= input(39);
output(4, 132) <= input(40);
output(4, 133) <= input(41);
output(4, 134) <= input(42);
output(4, 135) <= input(43);
output(4, 136) <= input(44);
output(4, 137) <= input(45);
output(4, 138) <= input(46);
output(4, 139) <= input(47);
output(4, 140) <= input(48);
output(4, 141) <= input(49);
output(4, 142) <= input(50);
output(4, 143) <= input(51);
output(4, 144) <= input(5);
output(4, 145) <= input(6);
output(4, 146) <= input(7);
output(4, 147) <= input(8);
output(4, 148) <= input(9);
output(4, 149) <= input(10);
output(4, 150) <= input(11);
output(4, 151) <= input(12);
output(4, 152) <= input(13);
output(4, 153) <= input(14);
output(4, 154) <= input(15);
output(4, 155) <= input(16);
output(4, 156) <= input(17);
output(4, 157) <= input(18);
output(4, 158) <= input(19);
output(4, 159) <= input(20);
output(4, 160) <= input(37);
output(4, 161) <= input(38);
output(4, 162) <= input(39);
output(4, 163) <= input(40);
output(4, 164) <= input(41);
output(4, 165) <= input(42);
output(4, 166) <= input(43);
output(4, 167) <= input(44);
output(4, 168) <= input(45);
output(4, 169) <= input(46);
output(4, 170) <= input(47);
output(4, 171) <= input(48);
output(4, 172) <= input(49);
output(4, 173) <= input(50);
output(4, 174) <= input(51);
output(4, 175) <= input(52);
output(4, 176) <= input(38);
output(4, 177) <= input(39);
output(4, 178) <= input(40);
output(4, 179) <= input(41);
output(4, 180) <= input(42);
output(4, 181) <= input(43);
output(4, 182) <= input(44);
output(4, 183) <= input(45);
output(4, 184) <= input(46);
output(4, 185) <= input(47);
output(4, 186) <= input(48);
output(4, 187) <= input(49);
output(4, 188) <= input(50);
output(4, 189) <= input(51);
output(4, 190) <= input(52);
output(4, 191) <= input(53);
output(4, 192) <= input(7);
output(4, 193) <= input(8);
output(4, 194) <= input(9);
output(4, 195) <= input(10);
output(4, 196) <= input(11);
output(4, 197) <= input(12);
output(4, 198) <= input(13);
output(4, 199) <= input(14);
output(4, 200) <= input(15);
output(4, 201) <= input(16);
output(4, 202) <= input(17);
output(4, 203) <= input(18);
output(4, 204) <= input(19);
output(4, 205) <= input(20);
output(4, 206) <= input(21);
output(4, 207) <= input(22);
output(4, 208) <= input(39);
output(4, 209) <= input(40);
output(4, 210) <= input(41);
output(4, 211) <= input(42);
output(4, 212) <= input(43);
output(4, 213) <= input(44);
output(4, 214) <= input(45);
output(4, 215) <= input(46);
output(4, 216) <= input(47);
output(4, 217) <= input(48);
output(4, 218) <= input(49);
output(4, 219) <= input(50);
output(4, 220) <= input(51);
output(4, 221) <= input(52);
output(4, 222) <= input(53);
output(4, 223) <= input(54);
output(4, 224) <= input(8);
output(4, 225) <= input(9);
output(4, 226) <= input(10);
output(4, 227) <= input(11);
output(4, 228) <= input(12);
output(4, 229) <= input(13);
output(4, 230) <= input(14);
output(4, 231) <= input(15);
output(4, 232) <= input(16);
output(4, 233) <= input(17);
output(4, 234) <= input(18);
output(4, 235) <= input(19);
output(4, 236) <= input(20);
output(4, 237) <= input(21);
output(4, 238) <= input(22);
output(4, 239) <= input(23);
output(4, 240) <= input(9);
output(4, 241) <= input(10);
output(4, 242) <= input(11);
output(4, 243) <= input(12);
output(4, 244) <= input(13);
output(4, 245) <= input(14);
output(4, 246) <= input(15);
output(4, 247) <= input(16);
output(4, 248) <= input(17);
output(4, 249) <= input(18);
output(4, 250) <= input(19);
output(4, 251) <= input(20);
output(4, 252) <= input(21);
output(4, 253) <= input(22);
output(4, 254) <= input(23);
output(4, 255) <= input(24);
output(5, 0) <= input(31);
output(5, 1) <= input(32);
output(5, 2) <= input(33);
output(5, 3) <= input(34);
output(5, 4) <= input(35);
output(5, 5) <= input(36);
output(5, 6) <= input(37);
output(5, 7) <= input(38);
output(5, 8) <= input(39);
output(5, 9) <= input(40);
output(5, 10) <= input(41);
output(5, 11) <= input(42);
output(5, 12) <= input(43);
output(5, 13) <= input(44);
output(5, 14) <= input(45);
output(5, 15) <= input(46);
output(5, 16) <= input(0);
output(5, 17) <= input(1);
output(5, 18) <= input(2);
output(5, 19) <= input(3);
output(5, 20) <= input(4);
output(5, 21) <= input(5);
output(5, 22) <= input(6);
output(5, 23) <= input(7);
output(5, 24) <= input(8);
output(5, 25) <= input(9);
output(5, 26) <= input(10);
output(5, 27) <= input(11);
output(5, 28) <= input(12);
output(5, 29) <= input(13);
output(5, 30) <= input(14);
output(5, 31) <= input(15);
output(5, 32) <= input(32);
output(5, 33) <= input(33);
output(5, 34) <= input(34);
output(5, 35) <= input(35);
output(5, 36) <= input(36);
output(5, 37) <= input(37);
output(5, 38) <= input(38);
output(5, 39) <= input(39);
output(5, 40) <= input(40);
output(5, 41) <= input(41);
output(5, 42) <= input(42);
output(5, 43) <= input(43);
output(5, 44) <= input(44);
output(5, 45) <= input(45);
output(5, 46) <= input(46);
output(5, 47) <= input(47);
output(5, 48) <= input(1);
output(5, 49) <= input(2);
output(5, 50) <= input(3);
output(5, 51) <= input(4);
output(5, 52) <= input(5);
output(5, 53) <= input(6);
output(5, 54) <= input(7);
output(5, 55) <= input(8);
output(5, 56) <= input(9);
output(5, 57) <= input(10);
output(5, 58) <= input(11);
output(5, 59) <= input(12);
output(5, 60) <= input(13);
output(5, 61) <= input(14);
output(5, 62) <= input(15);
output(5, 63) <= input(16);
output(5, 64) <= input(33);
output(5, 65) <= input(34);
output(5, 66) <= input(35);
output(5, 67) <= input(36);
output(5, 68) <= input(37);
output(5, 69) <= input(38);
output(5, 70) <= input(39);
output(5, 71) <= input(40);
output(5, 72) <= input(41);
output(5, 73) <= input(42);
output(5, 74) <= input(43);
output(5, 75) <= input(44);
output(5, 76) <= input(45);
output(5, 77) <= input(46);
output(5, 78) <= input(47);
output(5, 79) <= input(48);
output(5, 80) <= input(2);
output(5, 81) <= input(3);
output(5, 82) <= input(4);
output(5, 83) <= input(5);
output(5, 84) <= input(6);
output(5, 85) <= input(7);
output(5, 86) <= input(8);
output(5, 87) <= input(9);
output(5, 88) <= input(10);
output(5, 89) <= input(11);
output(5, 90) <= input(12);
output(5, 91) <= input(13);
output(5, 92) <= input(14);
output(5, 93) <= input(15);
output(5, 94) <= input(16);
output(5, 95) <= input(17);
output(5, 96) <= input(34);
output(5, 97) <= input(35);
output(5, 98) <= input(36);
output(5, 99) <= input(37);
output(5, 100) <= input(38);
output(5, 101) <= input(39);
output(5, 102) <= input(40);
output(5, 103) <= input(41);
output(5, 104) <= input(42);
output(5, 105) <= input(43);
output(5, 106) <= input(44);
output(5, 107) <= input(45);
output(5, 108) <= input(46);
output(5, 109) <= input(47);
output(5, 110) <= input(48);
output(5, 111) <= input(49);
output(5, 112) <= input(35);
output(5, 113) <= input(36);
output(5, 114) <= input(37);
output(5, 115) <= input(38);
output(5, 116) <= input(39);
output(5, 117) <= input(40);
output(5, 118) <= input(41);
output(5, 119) <= input(42);
output(5, 120) <= input(43);
output(5, 121) <= input(44);
output(5, 122) <= input(45);
output(5, 123) <= input(46);
output(5, 124) <= input(47);
output(5, 125) <= input(48);
output(5, 126) <= input(49);
output(5, 127) <= input(50);
output(5, 128) <= input(4);
output(5, 129) <= input(5);
output(5, 130) <= input(6);
output(5, 131) <= input(7);
output(5, 132) <= input(8);
output(5, 133) <= input(9);
output(5, 134) <= input(10);
output(5, 135) <= input(11);
output(5, 136) <= input(12);
output(5, 137) <= input(13);
output(5, 138) <= input(14);
output(5, 139) <= input(15);
output(5, 140) <= input(16);
output(5, 141) <= input(17);
output(5, 142) <= input(18);
output(5, 143) <= input(19);
output(5, 144) <= input(36);
output(5, 145) <= input(37);
output(5, 146) <= input(38);
output(5, 147) <= input(39);
output(5, 148) <= input(40);
output(5, 149) <= input(41);
output(5, 150) <= input(42);
output(5, 151) <= input(43);
output(5, 152) <= input(44);
output(5, 153) <= input(45);
output(5, 154) <= input(46);
output(5, 155) <= input(47);
output(5, 156) <= input(48);
output(5, 157) <= input(49);
output(5, 158) <= input(50);
output(5, 159) <= input(51);
output(5, 160) <= input(5);
output(5, 161) <= input(6);
output(5, 162) <= input(7);
output(5, 163) <= input(8);
output(5, 164) <= input(9);
output(5, 165) <= input(10);
output(5, 166) <= input(11);
output(5, 167) <= input(12);
output(5, 168) <= input(13);
output(5, 169) <= input(14);
output(5, 170) <= input(15);
output(5, 171) <= input(16);
output(5, 172) <= input(17);
output(5, 173) <= input(18);
output(5, 174) <= input(19);
output(5, 175) <= input(20);
output(5, 176) <= input(37);
output(5, 177) <= input(38);
output(5, 178) <= input(39);
output(5, 179) <= input(40);
output(5, 180) <= input(41);
output(5, 181) <= input(42);
output(5, 182) <= input(43);
output(5, 183) <= input(44);
output(5, 184) <= input(45);
output(5, 185) <= input(46);
output(5, 186) <= input(47);
output(5, 187) <= input(48);
output(5, 188) <= input(49);
output(5, 189) <= input(50);
output(5, 190) <= input(51);
output(5, 191) <= input(52);
output(5, 192) <= input(6);
output(5, 193) <= input(7);
output(5, 194) <= input(8);
output(5, 195) <= input(9);
output(5, 196) <= input(10);
output(5, 197) <= input(11);
output(5, 198) <= input(12);
output(5, 199) <= input(13);
output(5, 200) <= input(14);
output(5, 201) <= input(15);
output(5, 202) <= input(16);
output(5, 203) <= input(17);
output(5, 204) <= input(18);
output(5, 205) <= input(19);
output(5, 206) <= input(20);
output(5, 207) <= input(21);
output(5, 208) <= input(38);
output(5, 209) <= input(39);
output(5, 210) <= input(40);
output(5, 211) <= input(41);
output(5, 212) <= input(42);
output(5, 213) <= input(43);
output(5, 214) <= input(44);
output(5, 215) <= input(45);
output(5, 216) <= input(46);
output(5, 217) <= input(47);
output(5, 218) <= input(48);
output(5, 219) <= input(49);
output(5, 220) <= input(50);
output(5, 221) <= input(51);
output(5, 222) <= input(52);
output(5, 223) <= input(53);
output(5, 224) <= input(7);
output(5, 225) <= input(8);
output(5, 226) <= input(9);
output(5, 227) <= input(10);
output(5, 228) <= input(11);
output(5, 229) <= input(12);
output(5, 230) <= input(13);
output(5, 231) <= input(14);
output(5, 232) <= input(15);
output(5, 233) <= input(16);
output(5, 234) <= input(17);
output(5, 235) <= input(18);
output(5, 236) <= input(19);
output(5, 237) <= input(20);
output(5, 238) <= input(21);
output(5, 239) <= input(22);
output(5, 240) <= input(8);
output(5, 241) <= input(9);
output(5, 242) <= input(10);
output(5, 243) <= input(11);
output(5, 244) <= input(12);
output(5, 245) <= input(13);
output(5, 246) <= input(14);
output(5, 247) <= input(15);
output(5, 248) <= input(16);
output(5, 249) <= input(17);
output(5, 250) <= input(18);
output(5, 251) <= input(19);
output(5, 252) <= input(20);
output(5, 253) <= input(21);
output(5, 254) <= input(22);
output(5, 255) <= input(23);
when "0001" =>
output(0, 0) <= input(0);
output(0, 1) <= input(1);
output(0, 2) <= input(2);
output(0, 3) <= input(3);
output(0, 4) <= input(4);
output(0, 5) <= input(5);
output(0, 6) <= input(6);
output(0, 7) <= input(7);
output(0, 8) <= input(8);
output(0, 9) <= input(9);
output(0, 10) <= input(10);
output(0, 11) <= input(11);
output(0, 12) <= input(12);
output(0, 13) <= input(13);
output(0, 14) <= input(14);
output(0, 15) <= input(15);
output(0, 16) <= input(16);
output(0, 17) <= input(17);
output(0, 18) <= input(18);
output(0, 19) <= input(19);
output(0, 20) <= input(20);
output(0, 21) <= input(21);
output(0, 22) <= input(22);
output(0, 23) <= input(23);
output(0, 24) <= input(24);
output(0, 25) <= input(25);
output(0, 26) <= input(26);
output(0, 27) <= input(27);
output(0, 28) <= input(28);
output(0, 29) <= input(29);
output(0, 30) <= input(30);
output(0, 31) <= input(31);
output(0, 32) <= input(1);
output(0, 33) <= input(2);
output(0, 34) <= input(3);
output(0, 35) <= input(4);
output(0, 36) <= input(5);
output(0, 37) <= input(6);
output(0, 38) <= input(7);
output(0, 39) <= input(8);
output(0, 40) <= input(9);
output(0, 41) <= input(10);
output(0, 42) <= input(11);
output(0, 43) <= input(12);
output(0, 44) <= input(13);
output(0, 45) <= input(14);
output(0, 46) <= input(15);
output(0, 47) <= input(32);
output(0, 48) <= input(17);
output(0, 49) <= input(18);
output(0, 50) <= input(19);
output(0, 51) <= input(20);
output(0, 52) <= input(21);
output(0, 53) <= input(22);
output(0, 54) <= input(23);
output(0, 55) <= input(24);
output(0, 56) <= input(25);
output(0, 57) <= input(26);
output(0, 58) <= input(27);
output(0, 59) <= input(28);
output(0, 60) <= input(29);
output(0, 61) <= input(30);
output(0, 62) <= input(31);
output(0, 63) <= input(33);
output(0, 64) <= input(2);
output(0, 65) <= input(3);
output(0, 66) <= input(4);
output(0, 67) <= input(5);
output(0, 68) <= input(6);
output(0, 69) <= input(7);
output(0, 70) <= input(8);
output(0, 71) <= input(9);
output(0, 72) <= input(10);
output(0, 73) <= input(11);
output(0, 74) <= input(12);
output(0, 75) <= input(13);
output(0, 76) <= input(14);
output(0, 77) <= input(15);
output(0, 78) <= input(32);
output(0, 79) <= input(34);
output(0, 80) <= input(18);
output(0, 81) <= input(19);
output(0, 82) <= input(20);
output(0, 83) <= input(21);
output(0, 84) <= input(22);
output(0, 85) <= input(23);
output(0, 86) <= input(24);
output(0, 87) <= input(25);
output(0, 88) <= input(26);
output(0, 89) <= input(27);
output(0, 90) <= input(28);
output(0, 91) <= input(29);
output(0, 92) <= input(30);
output(0, 93) <= input(31);
output(0, 94) <= input(33);
output(0, 95) <= input(35);
output(0, 96) <= input(3);
output(0, 97) <= input(4);
output(0, 98) <= input(5);
output(0, 99) <= input(6);
output(0, 100) <= input(7);
output(0, 101) <= input(8);
output(0, 102) <= input(9);
output(0, 103) <= input(10);
output(0, 104) <= input(11);
output(0, 105) <= input(12);
output(0, 106) <= input(13);
output(0, 107) <= input(14);
output(0, 108) <= input(15);
output(0, 109) <= input(32);
output(0, 110) <= input(34);
output(0, 111) <= input(36);
output(0, 112) <= input(19);
output(0, 113) <= input(20);
output(0, 114) <= input(21);
output(0, 115) <= input(22);
output(0, 116) <= input(23);
output(0, 117) <= input(24);
output(0, 118) <= input(25);
output(0, 119) <= input(26);
output(0, 120) <= input(27);
output(0, 121) <= input(28);
output(0, 122) <= input(29);
output(0, 123) <= input(30);
output(0, 124) <= input(31);
output(0, 125) <= input(33);
output(0, 126) <= input(35);
output(0, 127) <= input(37);
output(0, 128) <= input(4);
output(0, 129) <= input(5);
output(0, 130) <= input(6);
output(0, 131) <= input(7);
output(0, 132) <= input(8);
output(0, 133) <= input(9);
output(0, 134) <= input(10);
output(0, 135) <= input(11);
output(0, 136) <= input(12);
output(0, 137) <= input(13);
output(0, 138) <= input(14);
output(0, 139) <= input(15);
output(0, 140) <= input(32);
output(0, 141) <= input(34);
output(0, 142) <= input(36);
output(0, 143) <= input(38);
output(0, 144) <= input(20);
output(0, 145) <= input(21);
output(0, 146) <= input(22);
output(0, 147) <= input(23);
output(0, 148) <= input(24);
output(0, 149) <= input(25);
output(0, 150) <= input(26);
output(0, 151) <= input(27);
output(0, 152) <= input(28);
output(0, 153) <= input(29);
output(0, 154) <= input(30);
output(0, 155) <= input(31);
output(0, 156) <= input(33);
output(0, 157) <= input(35);
output(0, 158) <= input(37);
output(0, 159) <= input(39);
output(0, 160) <= input(5);
output(0, 161) <= input(6);
output(0, 162) <= input(7);
output(0, 163) <= input(8);
output(0, 164) <= input(9);
output(0, 165) <= input(10);
output(0, 166) <= input(11);
output(0, 167) <= input(12);
output(0, 168) <= input(13);
output(0, 169) <= input(14);
output(0, 170) <= input(15);
output(0, 171) <= input(32);
output(0, 172) <= input(34);
output(0, 173) <= input(36);
output(0, 174) <= input(38);
output(0, 175) <= input(40);
output(0, 176) <= input(21);
output(0, 177) <= input(22);
output(0, 178) <= input(23);
output(0, 179) <= input(24);
output(0, 180) <= input(25);
output(0, 181) <= input(26);
output(0, 182) <= input(27);
output(0, 183) <= input(28);
output(0, 184) <= input(29);
output(0, 185) <= input(30);
output(0, 186) <= input(31);
output(0, 187) <= input(33);
output(0, 188) <= input(35);
output(0, 189) <= input(37);
output(0, 190) <= input(39);
output(0, 191) <= input(41);
output(0, 192) <= input(6);
output(0, 193) <= input(7);
output(0, 194) <= input(8);
output(0, 195) <= input(9);
output(0, 196) <= input(10);
output(0, 197) <= input(11);
output(0, 198) <= input(12);
output(0, 199) <= input(13);
output(0, 200) <= input(14);
output(0, 201) <= input(15);
output(0, 202) <= input(32);
output(0, 203) <= input(34);
output(0, 204) <= input(36);
output(0, 205) <= input(38);
output(0, 206) <= input(40);
output(0, 207) <= input(42);
output(0, 208) <= input(22);
output(0, 209) <= input(23);
output(0, 210) <= input(24);
output(0, 211) <= input(25);
output(0, 212) <= input(26);
output(0, 213) <= input(27);
output(0, 214) <= input(28);
output(0, 215) <= input(29);
output(0, 216) <= input(30);
output(0, 217) <= input(31);
output(0, 218) <= input(33);
output(0, 219) <= input(35);
output(0, 220) <= input(37);
output(0, 221) <= input(39);
output(0, 222) <= input(41);
output(0, 223) <= input(43);
output(0, 224) <= input(7);
output(0, 225) <= input(8);
output(0, 226) <= input(9);
output(0, 227) <= input(10);
output(0, 228) <= input(11);
output(0, 229) <= input(12);
output(0, 230) <= input(13);
output(0, 231) <= input(14);
output(0, 232) <= input(15);
output(0, 233) <= input(32);
output(0, 234) <= input(34);
output(0, 235) <= input(36);
output(0, 236) <= input(38);
output(0, 237) <= input(40);
output(0, 238) <= input(42);
output(0, 239) <= input(44);
output(0, 240) <= input(23);
output(0, 241) <= input(24);
output(0, 242) <= input(25);
output(0, 243) <= input(26);
output(0, 244) <= input(27);
output(0, 245) <= input(28);
output(0, 246) <= input(29);
output(0, 247) <= input(30);
output(0, 248) <= input(31);
output(0, 249) <= input(33);
output(0, 250) <= input(35);
output(0, 251) <= input(37);
output(0, 252) <= input(39);
output(0, 253) <= input(41);
output(0, 254) <= input(43);
output(0, 255) <= input(45);
output(1, 0) <= input(46);
output(1, 1) <= input(16);
output(1, 2) <= input(17);
output(1, 3) <= input(18);
output(1, 4) <= input(19);
output(1, 5) <= input(20);
output(1, 6) <= input(21);
output(1, 7) <= input(22);
output(1, 8) <= input(23);
output(1, 9) <= input(24);
output(1, 10) <= input(25);
output(1, 11) <= input(26);
output(1, 12) <= input(27);
output(1, 13) <= input(28);
output(1, 14) <= input(29);
output(1, 15) <= input(30);
output(1, 16) <= input(0);
output(1, 17) <= input(1);
output(1, 18) <= input(2);
output(1, 19) <= input(3);
output(1, 20) <= input(4);
output(1, 21) <= input(5);
output(1, 22) <= input(6);
output(1, 23) <= input(7);
output(1, 24) <= input(8);
output(1, 25) <= input(9);
output(1, 26) <= input(10);
output(1, 27) <= input(11);
output(1, 28) <= input(12);
output(1, 29) <= input(13);
output(1, 30) <= input(14);
output(1, 31) <= input(15);
output(1, 32) <= input(16);
output(1, 33) <= input(17);
output(1, 34) <= input(18);
output(1, 35) <= input(19);
output(1, 36) <= input(20);
output(1, 37) <= input(21);
output(1, 38) <= input(22);
output(1, 39) <= input(23);
output(1, 40) <= input(24);
output(1, 41) <= input(25);
output(1, 42) <= input(26);
output(1, 43) <= input(27);
output(1, 44) <= input(28);
output(1, 45) <= input(29);
output(1, 46) <= input(30);
output(1, 47) <= input(31);
output(1, 48) <= input(1);
output(1, 49) <= input(2);
output(1, 50) <= input(3);
output(1, 51) <= input(4);
output(1, 52) <= input(5);
output(1, 53) <= input(6);
output(1, 54) <= input(7);
output(1, 55) <= input(8);
output(1, 56) <= input(9);
output(1, 57) <= input(10);
output(1, 58) <= input(11);
output(1, 59) <= input(12);
output(1, 60) <= input(13);
output(1, 61) <= input(14);
output(1, 62) <= input(15);
output(1, 63) <= input(32);
output(1, 64) <= input(17);
output(1, 65) <= input(18);
output(1, 66) <= input(19);
output(1, 67) <= input(20);
output(1, 68) <= input(21);
output(1, 69) <= input(22);
output(1, 70) <= input(23);
output(1, 71) <= input(24);
output(1, 72) <= input(25);
output(1, 73) <= input(26);
output(1, 74) <= input(27);
output(1, 75) <= input(28);
output(1, 76) <= input(29);
output(1, 77) <= input(30);
output(1, 78) <= input(31);
output(1, 79) <= input(33);
output(1, 80) <= input(2);
output(1, 81) <= input(3);
output(1, 82) <= input(4);
output(1, 83) <= input(5);
output(1, 84) <= input(6);
output(1, 85) <= input(7);
output(1, 86) <= input(8);
output(1, 87) <= input(9);
output(1, 88) <= input(10);
output(1, 89) <= input(11);
output(1, 90) <= input(12);
output(1, 91) <= input(13);
output(1, 92) <= input(14);
output(1, 93) <= input(15);
output(1, 94) <= input(32);
output(1, 95) <= input(34);
output(1, 96) <= input(18);
output(1, 97) <= input(19);
output(1, 98) <= input(20);
output(1, 99) <= input(21);
output(1, 100) <= input(22);
output(1, 101) <= input(23);
output(1, 102) <= input(24);
output(1, 103) <= input(25);
output(1, 104) <= input(26);
output(1, 105) <= input(27);
output(1, 106) <= input(28);
output(1, 107) <= input(29);
output(1, 108) <= input(30);
output(1, 109) <= input(31);
output(1, 110) <= input(33);
output(1, 111) <= input(35);
output(1, 112) <= input(3);
output(1, 113) <= input(4);
output(1, 114) <= input(5);
output(1, 115) <= input(6);
output(1, 116) <= input(7);
output(1, 117) <= input(8);
output(1, 118) <= input(9);
output(1, 119) <= input(10);
output(1, 120) <= input(11);
output(1, 121) <= input(12);
output(1, 122) <= input(13);
output(1, 123) <= input(14);
output(1, 124) <= input(15);
output(1, 125) <= input(32);
output(1, 126) <= input(34);
output(1, 127) <= input(36);
output(1, 128) <= input(3);
output(1, 129) <= input(4);
output(1, 130) <= input(5);
output(1, 131) <= input(6);
output(1, 132) <= input(7);
output(1, 133) <= input(8);
output(1, 134) <= input(9);
output(1, 135) <= input(10);
output(1, 136) <= input(11);
output(1, 137) <= input(12);
output(1, 138) <= input(13);
output(1, 139) <= input(14);
output(1, 140) <= input(15);
output(1, 141) <= input(32);
output(1, 142) <= input(34);
output(1, 143) <= input(36);
output(1, 144) <= input(19);
output(1, 145) <= input(20);
output(1, 146) <= input(21);
output(1, 147) <= input(22);
output(1, 148) <= input(23);
output(1, 149) <= input(24);
output(1, 150) <= input(25);
output(1, 151) <= input(26);
output(1, 152) <= input(27);
output(1, 153) <= input(28);
output(1, 154) <= input(29);
output(1, 155) <= input(30);
output(1, 156) <= input(31);
output(1, 157) <= input(33);
output(1, 158) <= input(35);
output(1, 159) <= input(37);
output(1, 160) <= input(4);
output(1, 161) <= input(5);
output(1, 162) <= input(6);
output(1, 163) <= input(7);
output(1, 164) <= input(8);
output(1, 165) <= input(9);
output(1, 166) <= input(10);
output(1, 167) <= input(11);
output(1, 168) <= input(12);
output(1, 169) <= input(13);
output(1, 170) <= input(14);
output(1, 171) <= input(15);
output(1, 172) <= input(32);
output(1, 173) <= input(34);
output(1, 174) <= input(36);
output(1, 175) <= input(38);
output(1, 176) <= input(20);
output(1, 177) <= input(21);
output(1, 178) <= input(22);
output(1, 179) <= input(23);
output(1, 180) <= input(24);
output(1, 181) <= input(25);
output(1, 182) <= input(26);
output(1, 183) <= input(27);
output(1, 184) <= input(28);
output(1, 185) <= input(29);
output(1, 186) <= input(30);
output(1, 187) <= input(31);
output(1, 188) <= input(33);
output(1, 189) <= input(35);
output(1, 190) <= input(37);
output(1, 191) <= input(39);
output(1, 192) <= input(5);
output(1, 193) <= input(6);
output(1, 194) <= input(7);
output(1, 195) <= input(8);
output(1, 196) <= input(9);
output(1, 197) <= input(10);
output(1, 198) <= input(11);
output(1, 199) <= input(12);
output(1, 200) <= input(13);
output(1, 201) <= input(14);
output(1, 202) <= input(15);
output(1, 203) <= input(32);
output(1, 204) <= input(34);
output(1, 205) <= input(36);
output(1, 206) <= input(38);
output(1, 207) <= input(40);
output(1, 208) <= input(21);
output(1, 209) <= input(22);
output(1, 210) <= input(23);
output(1, 211) <= input(24);
output(1, 212) <= input(25);
output(1, 213) <= input(26);
output(1, 214) <= input(27);
output(1, 215) <= input(28);
output(1, 216) <= input(29);
output(1, 217) <= input(30);
output(1, 218) <= input(31);
output(1, 219) <= input(33);
output(1, 220) <= input(35);
output(1, 221) <= input(37);
output(1, 222) <= input(39);
output(1, 223) <= input(41);
output(1, 224) <= input(6);
output(1, 225) <= input(7);
output(1, 226) <= input(8);
output(1, 227) <= input(9);
output(1, 228) <= input(10);
output(1, 229) <= input(11);
output(1, 230) <= input(12);
output(1, 231) <= input(13);
output(1, 232) <= input(14);
output(1, 233) <= input(15);
output(1, 234) <= input(32);
output(1, 235) <= input(34);
output(1, 236) <= input(36);
output(1, 237) <= input(38);
output(1, 238) <= input(40);
output(1, 239) <= input(42);
output(1, 240) <= input(22);
output(1, 241) <= input(23);
output(1, 242) <= input(24);
output(1, 243) <= input(25);
output(1, 244) <= input(26);
output(1, 245) <= input(27);
output(1, 246) <= input(28);
output(1, 247) <= input(29);
output(1, 248) <= input(30);
output(1, 249) <= input(31);
output(1, 250) <= input(33);
output(1, 251) <= input(35);
output(1, 252) <= input(37);
output(1, 253) <= input(39);
output(1, 254) <= input(41);
output(1, 255) <= input(43);
output(2, 0) <= input(46);
output(2, 1) <= input(16);
output(2, 2) <= input(17);
output(2, 3) <= input(18);
output(2, 4) <= input(19);
output(2, 5) <= input(20);
output(2, 6) <= input(21);
output(2, 7) <= input(22);
output(2, 8) <= input(23);
output(2, 9) <= input(24);
output(2, 10) <= input(25);
output(2, 11) <= input(26);
output(2, 12) <= input(27);
output(2, 13) <= input(28);
output(2, 14) <= input(29);
output(2, 15) <= input(30);
output(2, 16) <= input(0);
output(2, 17) <= input(1);
output(2, 18) <= input(2);
output(2, 19) <= input(3);
output(2, 20) <= input(4);
output(2, 21) <= input(5);
output(2, 22) <= input(6);
output(2, 23) <= input(7);
output(2, 24) <= input(8);
output(2, 25) <= input(9);
output(2, 26) <= input(10);
output(2, 27) <= input(11);
output(2, 28) <= input(12);
output(2, 29) <= input(13);
output(2, 30) <= input(14);
output(2, 31) <= input(15);
output(2, 32) <= input(16);
output(2, 33) <= input(17);
output(2, 34) <= input(18);
output(2, 35) <= input(19);
output(2, 36) <= input(20);
output(2, 37) <= input(21);
output(2, 38) <= input(22);
output(2, 39) <= input(23);
output(2, 40) <= input(24);
output(2, 41) <= input(25);
output(2, 42) <= input(26);
output(2, 43) <= input(27);
output(2, 44) <= input(28);
output(2, 45) <= input(29);
output(2, 46) <= input(30);
output(2, 47) <= input(31);
output(2, 48) <= input(1);
output(2, 49) <= input(2);
output(2, 50) <= input(3);
output(2, 51) <= input(4);
output(2, 52) <= input(5);
output(2, 53) <= input(6);
output(2, 54) <= input(7);
output(2, 55) <= input(8);
output(2, 56) <= input(9);
output(2, 57) <= input(10);
output(2, 58) <= input(11);
output(2, 59) <= input(12);
output(2, 60) <= input(13);
output(2, 61) <= input(14);
output(2, 62) <= input(15);
output(2, 63) <= input(32);
output(2, 64) <= input(1);
output(2, 65) <= input(2);
output(2, 66) <= input(3);
output(2, 67) <= input(4);
output(2, 68) <= input(5);
output(2, 69) <= input(6);
output(2, 70) <= input(7);
output(2, 71) <= input(8);
output(2, 72) <= input(9);
output(2, 73) <= input(10);
output(2, 74) <= input(11);
output(2, 75) <= input(12);
output(2, 76) <= input(13);
output(2, 77) <= input(14);
output(2, 78) <= input(15);
output(2, 79) <= input(32);
output(2, 80) <= input(17);
output(2, 81) <= input(18);
output(2, 82) <= input(19);
output(2, 83) <= input(20);
output(2, 84) <= input(21);
output(2, 85) <= input(22);
output(2, 86) <= input(23);
output(2, 87) <= input(24);
output(2, 88) <= input(25);
output(2, 89) <= input(26);
output(2, 90) <= input(27);
output(2, 91) <= input(28);
output(2, 92) <= input(29);
output(2, 93) <= input(30);
output(2, 94) <= input(31);
output(2, 95) <= input(33);
output(2, 96) <= input(2);
output(2, 97) <= input(3);
output(2, 98) <= input(4);
output(2, 99) <= input(5);
output(2, 100) <= input(6);
output(2, 101) <= input(7);
output(2, 102) <= input(8);
output(2, 103) <= input(9);
output(2, 104) <= input(10);
output(2, 105) <= input(11);
output(2, 106) <= input(12);
output(2, 107) <= input(13);
output(2, 108) <= input(14);
output(2, 109) <= input(15);
output(2, 110) <= input(32);
output(2, 111) <= input(34);
output(2, 112) <= input(18);
output(2, 113) <= input(19);
output(2, 114) <= input(20);
output(2, 115) <= input(21);
output(2, 116) <= input(22);
output(2, 117) <= input(23);
output(2, 118) <= input(24);
output(2, 119) <= input(25);
output(2, 120) <= input(26);
output(2, 121) <= input(27);
output(2, 122) <= input(28);
output(2, 123) <= input(29);
output(2, 124) <= input(30);
output(2, 125) <= input(31);
output(2, 126) <= input(33);
output(2, 127) <= input(35);
output(2, 128) <= input(18);
output(2, 129) <= input(19);
output(2, 130) <= input(20);
output(2, 131) <= input(21);
output(2, 132) <= input(22);
output(2, 133) <= input(23);
output(2, 134) <= input(24);
output(2, 135) <= input(25);
output(2, 136) <= input(26);
output(2, 137) <= input(27);
output(2, 138) <= input(28);
output(2, 139) <= input(29);
output(2, 140) <= input(30);
output(2, 141) <= input(31);
output(2, 142) <= input(33);
output(2, 143) <= input(35);
output(2, 144) <= input(3);
output(2, 145) <= input(4);
output(2, 146) <= input(5);
output(2, 147) <= input(6);
output(2, 148) <= input(7);
output(2, 149) <= input(8);
output(2, 150) <= input(9);
output(2, 151) <= input(10);
output(2, 152) <= input(11);
output(2, 153) <= input(12);
output(2, 154) <= input(13);
output(2, 155) <= input(14);
output(2, 156) <= input(15);
output(2, 157) <= input(32);
output(2, 158) <= input(34);
output(2, 159) <= input(36);
output(2, 160) <= input(19);
output(2, 161) <= input(20);
output(2, 162) <= input(21);
output(2, 163) <= input(22);
output(2, 164) <= input(23);
output(2, 165) <= input(24);
output(2, 166) <= input(25);
output(2, 167) <= input(26);
output(2, 168) <= input(27);
output(2, 169) <= input(28);
output(2, 170) <= input(29);
output(2, 171) <= input(30);
output(2, 172) <= input(31);
output(2, 173) <= input(33);
output(2, 174) <= input(35);
output(2, 175) <= input(37);
output(2, 176) <= input(4);
output(2, 177) <= input(5);
output(2, 178) <= input(6);
output(2, 179) <= input(7);
output(2, 180) <= input(8);
output(2, 181) <= input(9);
output(2, 182) <= input(10);
output(2, 183) <= input(11);
output(2, 184) <= input(12);
output(2, 185) <= input(13);
output(2, 186) <= input(14);
output(2, 187) <= input(15);
output(2, 188) <= input(32);
output(2, 189) <= input(34);
output(2, 190) <= input(36);
output(2, 191) <= input(38);
output(2, 192) <= input(4);
output(2, 193) <= input(5);
output(2, 194) <= input(6);
output(2, 195) <= input(7);
output(2, 196) <= input(8);
output(2, 197) <= input(9);
output(2, 198) <= input(10);
output(2, 199) <= input(11);
output(2, 200) <= input(12);
output(2, 201) <= input(13);
output(2, 202) <= input(14);
output(2, 203) <= input(15);
output(2, 204) <= input(32);
output(2, 205) <= input(34);
output(2, 206) <= input(36);
output(2, 207) <= input(38);
output(2, 208) <= input(20);
output(2, 209) <= input(21);
output(2, 210) <= input(22);
output(2, 211) <= input(23);
output(2, 212) <= input(24);
output(2, 213) <= input(25);
output(2, 214) <= input(26);
output(2, 215) <= input(27);
output(2, 216) <= input(28);
output(2, 217) <= input(29);
output(2, 218) <= input(30);
output(2, 219) <= input(31);
output(2, 220) <= input(33);
output(2, 221) <= input(35);
output(2, 222) <= input(37);
output(2, 223) <= input(39);
output(2, 224) <= input(5);
output(2, 225) <= input(6);
output(2, 226) <= input(7);
output(2, 227) <= input(8);
output(2, 228) <= input(9);
output(2, 229) <= input(10);
output(2, 230) <= input(11);
output(2, 231) <= input(12);
output(2, 232) <= input(13);
output(2, 233) <= input(14);
output(2, 234) <= input(15);
output(2, 235) <= input(32);
output(2, 236) <= input(34);
output(2, 237) <= input(36);
output(2, 238) <= input(38);
output(2, 239) <= input(40);
output(2, 240) <= input(21);
output(2, 241) <= input(22);
output(2, 242) <= input(23);
output(2, 243) <= input(24);
output(2, 244) <= input(25);
output(2, 245) <= input(26);
output(2, 246) <= input(27);
output(2, 247) <= input(28);
output(2, 248) <= input(29);
output(2, 249) <= input(30);
output(2, 250) <= input(31);
output(2, 251) <= input(33);
output(2, 252) <= input(35);
output(2, 253) <= input(37);
output(2, 254) <= input(39);
output(2, 255) <= input(41);
output(3, 0) <= input(46);
output(3, 1) <= input(16);
output(3, 2) <= input(17);
output(3, 3) <= input(18);
output(3, 4) <= input(19);
output(3, 5) <= input(20);
output(3, 6) <= input(21);
output(3, 7) <= input(22);
output(3, 8) <= input(23);
output(3, 9) <= input(24);
output(3, 10) <= input(25);
output(3, 11) <= input(26);
output(3, 12) <= input(27);
output(3, 13) <= input(28);
output(3, 14) <= input(29);
output(3, 15) <= input(30);
output(3, 16) <= input(0);
output(3, 17) <= input(1);
output(3, 18) <= input(2);
output(3, 19) <= input(3);
output(3, 20) <= input(4);
output(3, 21) <= input(5);
output(3, 22) <= input(6);
output(3, 23) <= input(7);
output(3, 24) <= input(8);
output(3, 25) <= input(9);
output(3, 26) <= input(10);
output(3, 27) <= input(11);
output(3, 28) <= input(12);
output(3, 29) <= input(13);
output(3, 30) <= input(14);
output(3, 31) <= input(15);
output(3, 32) <= input(0);
output(3, 33) <= input(1);
output(3, 34) <= input(2);
output(3, 35) <= input(3);
output(3, 36) <= input(4);
output(3, 37) <= input(5);
output(3, 38) <= input(6);
output(3, 39) <= input(7);
output(3, 40) <= input(8);
output(3, 41) <= input(9);
output(3, 42) <= input(10);
output(3, 43) <= input(11);
output(3, 44) <= input(12);
output(3, 45) <= input(13);
output(3, 46) <= input(14);
output(3, 47) <= input(15);
output(3, 48) <= input(16);
output(3, 49) <= input(17);
output(3, 50) <= input(18);
output(3, 51) <= input(19);
output(3, 52) <= input(20);
output(3, 53) <= input(21);
output(3, 54) <= input(22);
output(3, 55) <= input(23);
output(3, 56) <= input(24);
output(3, 57) <= input(25);
output(3, 58) <= input(26);
output(3, 59) <= input(27);
output(3, 60) <= input(28);
output(3, 61) <= input(29);
output(3, 62) <= input(30);
output(3, 63) <= input(31);
output(3, 64) <= input(1);
output(3, 65) <= input(2);
output(3, 66) <= input(3);
output(3, 67) <= input(4);
output(3, 68) <= input(5);
output(3, 69) <= input(6);
output(3, 70) <= input(7);
output(3, 71) <= input(8);
output(3, 72) <= input(9);
output(3, 73) <= input(10);
output(3, 74) <= input(11);
output(3, 75) <= input(12);
output(3, 76) <= input(13);
output(3, 77) <= input(14);
output(3, 78) <= input(15);
output(3, 79) <= input(32);
output(3, 80) <= input(1);
output(3, 81) <= input(2);
output(3, 82) <= input(3);
output(3, 83) <= input(4);
output(3, 84) <= input(5);
output(3, 85) <= input(6);
output(3, 86) <= input(7);
output(3, 87) <= input(8);
output(3, 88) <= input(9);
output(3, 89) <= input(10);
output(3, 90) <= input(11);
output(3, 91) <= input(12);
output(3, 92) <= input(13);
output(3, 93) <= input(14);
output(3, 94) <= input(15);
output(3, 95) <= input(32);
output(3, 96) <= input(17);
output(3, 97) <= input(18);
output(3, 98) <= input(19);
output(3, 99) <= input(20);
output(3, 100) <= input(21);
output(3, 101) <= input(22);
output(3, 102) <= input(23);
output(3, 103) <= input(24);
output(3, 104) <= input(25);
output(3, 105) <= input(26);
output(3, 106) <= input(27);
output(3, 107) <= input(28);
output(3, 108) <= input(29);
output(3, 109) <= input(30);
output(3, 110) <= input(31);
output(3, 111) <= input(33);
output(3, 112) <= input(2);
output(3, 113) <= input(3);
output(3, 114) <= input(4);
output(3, 115) <= input(5);
output(3, 116) <= input(6);
output(3, 117) <= input(7);
output(3, 118) <= input(8);
output(3, 119) <= input(9);
output(3, 120) <= input(10);
output(3, 121) <= input(11);
output(3, 122) <= input(12);
output(3, 123) <= input(13);
output(3, 124) <= input(14);
output(3, 125) <= input(15);
output(3, 126) <= input(32);
output(3, 127) <= input(34);
output(3, 128) <= input(2);
output(3, 129) <= input(3);
output(3, 130) <= input(4);
output(3, 131) <= input(5);
output(3, 132) <= input(6);
output(3, 133) <= input(7);
output(3, 134) <= input(8);
output(3, 135) <= input(9);
output(3, 136) <= input(10);
output(3, 137) <= input(11);
output(3, 138) <= input(12);
output(3, 139) <= input(13);
output(3, 140) <= input(14);
output(3, 141) <= input(15);
output(3, 142) <= input(32);
output(3, 143) <= input(34);
output(3, 144) <= input(18);
output(3, 145) <= input(19);
output(3, 146) <= input(20);
output(3, 147) <= input(21);
output(3, 148) <= input(22);
output(3, 149) <= input(23);
output(3, 150) <= input(24);
output(3, 151) <= input(25);
output(3, 152) <= input(26);
output(3, 153) <= input(27);
output(3, 154) <= input(28);
output(3, 155) <= input(29);
output(3, 156) <= input(30);
output(3, 157) <= input(31);
output(3, 158) <= input(33);
output(3, 159) <= input(35);
output(3, 160) <= input(18);
output(3, 161) <= input(19);
output(3, 162) <= input(20);
output(3, 163) <= input(21);
output(3, 164) <= input(22);
output(3, 165) <= input(23);
output(3, 166) <= input(24);
output(3, 167) <= input(25);
output(3, 168) <= input(26);
output(3, 169) <= input(27);
output(3, 170) <= input(28);
output(3, 171) <= input(29);
output(3, 172) <= input(30);
output(3, 173) <= input(31);
output(3, 174) <= input(33);
output(3, 175) <= input(35);
output(3, 176) <= input(3);
output(3, 177) <= input(4);
output(3, 178) <= input(5);
output(3, 179) <= input(6);
output(3, 180) <= input(7);
output(3, 181) <= input(8);
output(3, 182) <= input(9);
output(3, 183) <= input(10);
output(3, 184) <= input(11);
output(3, 185) <= input(12);
output(3, 186) <= input(13);
output(3, 187) <= input(14);
output(3, 188) <= input(15);
output(3, 189) <= input(32);
output(3, 190) <= input(34);
output(3, 191) <= input(36);
output(3, 192) <= input(19);
output(3, 193) <= input(20);
output(3, 194) <= input(21);
output(3, 195) <= input(22);
output(3, 196) <= input(23);
output(3, 197) <= input(24);
output(3, 198) <= input(25);
output(3, 199) <= input(26);
output(3, 200) <= input(27);
output(3, 201) <= input(28);
output(3, 202) <= input(29);
output(3, 203) <= input(30);
output(3, 204) <= input(31);
output(3, 205) <= input(33);
output(3, 206) <= input(35);
output(3, 207) <= input(37);
output(3, 208) <= input(19);
output(3, 209) <= input(20);
output(3, 210) <= input(21);
output(3, 211) <= input(22);
output(3, 212) <= input(23);
output(3, 213) <= input(24);
output(3, 214) <= input(25);
output(3, 215) <= input(26);
output(3, 216) <= input(27);
output(3, 217) <= input(28);
output(3, 218) <= input(29);
output(3, 219) <= input(30);
output(3, 220) <= input(31);
output(3, 221) <= input(33);
output(3, 222) <= input(35);
output(3, 223) <= input(37);
output(3, 224) <= input(4);
output(3, 225) <= input(5);
output(3, 226) <= input(6);
output(3, 227) <= input(7);
output(3, 228) <= input(8);
output(3, 229) <= input(9);
output(3, 230) <= input(10);
output(3, 231) <= input(11);
output(3, 232) <= input(12);
output(3, 233) <= input(13);
output(3, 234) <= input(14);
output(3, 235) <= input(15);
output(3, 236) <= input(32);
output(3, 237) <= input(34);
output(3, 238) <= input(36);
output(3, 239) <= input(38);
output(3, 240) <= input(20);
output(3, 241) <= input(21);
output(3, 242) <= input(22);
output(3, 243) <= input(23);
output(3, 244) <= input(24);
output(3, 245) <= input(25);
output(3, 246) <= input(26);
output(3, 247) <= input(27);
output(3, 248) <= input(28);
output(3, 249) <= input(29);
output(3, 250) <= input(30);
output(3, 251) <= input(31);
output(3, 252) <= input(33);
output(3, 253) <= input(35);
output(3, 254) <= input(37);
output(3, 255) <= input(39);
output(4, 0) <= input(46);
output(4, 1) <= input(16);
output(4, 2) <= input(17);
output(4, 3) <= input(18);
output(4, 4) <= input(19);
output(4, 5) <= input(20);
output(4, 6) <= input(21);
output(4, 7) <= input(22);
output(4, 8) <= input(23);
output(4, 9) <= input(24);
output(4, 10) <= input(25);
output(4, 11) <= input(26);
output(4, 12) <= input(27);
output(4, 13) <= input(28);
output(4, 14) <= input(29);
output(4, 15) <= input(30);
output(4, 16) <= input(0);
output(4, 17) <= input(1);
output(4, 18) <= input(2);
output(4, 19) <= input(3);
output(4, 20) <= input(4);
output(4, 21) <= input(5);
output(4, 22) <= input(6);
output(4, 23) <= input(7);
output(4, 24) <= input(8);
output(4, 25) <= input(9);
output(4, 26) <= input(10);
output(4, 27) <= input(11);
output(4, 28) <= input(12);
output(4, 29) <= input(13);
output(4, 30) <= input(14);
output(4, 31) <= input(15);
output(4, 32) <= input(0);
output(4, 33) <= input(1);
output(4, 34) <= input(2);
output(4, 35) <= input(3);
output(4, 36) <= input(4);
output(4, 37) <= input(5);
output(4, 38) <= input(6);
output(4, 39) <= input(7);
output(4, 40) <= input(8);
output(4, 41) <= input(9);
output(4, 42) <= input(10);
output(4, 43) <= input(11);
output(4, 44) <= input(12);
output(4, 45) <= input(13);
output(4, 46) <= input(14);
output(4, 47) <= input(15);
output(4, 48) <= input(16);
output(4, 49) <= input(17);
output(4, 50) <= input(18);
output(4, 51) <= input(19);
output(4, 52) <= input(20);
output(4, 53) <= input(21);
output(4, 54) <= input(22);
output(4, 55) <= input(23);
output(4, 56) <= input(24);
output(4, 57) <= input(25);
output(4, 58) <= input(26);
output(4, 59) <= input(27);
output(4, 60) <= input(28);
output(4, 61) <= input(29);
output(4, 62) <= input(30);
output(4, 63) <= input(31);
output(4, 64) <= input(16);
output(4, 65) <= input(17);
output(4, 66) <= input(18);
output(4, 67) <= input(19);
output(4, 68) <= input(20);
output(4, 69) <= input(21);
output(4, 70) <= input(22);
output(4, 71) <= input(23);
output(4, 72) <= input(24);
output(4, 73) <= input(25);
output(4, 74) <= input(26);
output(4, 75) <= input(27);
output(4, 76) <= input(28);
output(4, 77) <= input(29);
output(4, 78) <= input(30);
output(4, 79) <= input(31);
output(4, 80) <= input(1);
output(4, 81) <= input(2);
output(4, 82) <= input(3);
output(4, 83) <= input(4);
output(4, 84) <= input(5);
output(4, 85) <= input(6);
output(4, 86) <= input(7);
output(4, 87) <= input(8);
output(4, 88) <= input(9);
output(4, 89) <= input(10);
output(4, 90) <= input(11);
output(4, 91) <= input(12);
output(4, 92) <= input(13);
output(4, 93) <= input(14);
output(4, 94) <= input(15);
output(4, 95) <= input(32);
output(4, 96) <= input(1);
output(4, 97) <= input(2);
output(4, 98) <= input(3);
output(4, 99) <= input(4);
output(4, 100) <= input(5);
output(4, 101) <= input(6);
output(4, 102) <= input(7);
output(4, 103) <= input(8);
output(4, 104) <= input(9);
output(4, 105) <= input(10);
output(4, 106) <= input(11);
output(4, 107) <= input(12);
output(4, 108) <= input(13);
output(4, 109) <= input(14);
output(4, 110) <= input(15);
output(4, 111) <= input(32);
output(4, 112) <= input(17);
output(4, 113) <= input(18);
output(4, 114) <= input(19);
output(4, 115) <= input(20);
output(4, 116) <= input(21);
output(4, 117) <= input(22);
output(4, 118) <= input(23);
output(4, 119) <= input(24);
output(4, 120) <= input(25);
output(4, 121) <= input(26);
output(4, 122) <= input(27);
output(4, 123) <= input(28);
output(4, 124) <= input(29);
output(4, 125) <= input(30);
output(4, 126) <= input(31);
output(4, 127) <= input(33);
output(4, 128) <= input(17);
output(4, 129) <= input(18);
output(4, 130) <= input(19);
output(4, 131) <= input(20);
output(4, 132) <= input(21);
output(4, 133) <= input(22);
output(4, 134) <= input(23);
output(4, 135) <= input(24);
output(4, 136) <= input(25);
output(4, 137) <= input(26);
output(4, 138) <= input(27);
output(4, 139) <= input(28);
output(4, 140) <= input(29);
output(4, 141) <= input(30);
output(4, 142) <= input(31);
output(4, 143) <= input(33);
output(4, 144) <= input(2);
output(4, 145) <= input(3);
output(4, 146) <= input(4);
output(4, 147) <= input(5);
output(4, 148) <= input(6);
output(4, 149) <= input(7);
output(4, 150) <= input(8);
output(4, 151) <= input(9);
output(4, 152) <= input(10);
output(4, 153) <= input(11);
output(4, 154) <= input(12);
output(4, 155) <= input(13);
output(4, 156) <= input(14);
output(4, 157) <= input(15);
output(4, 158) <= input(32);
output(4, 159) <= input(34);
output(4, 160) <= input(2);
output(4, 161) <= input(3);
output(4, 162) <= input(4);
output(4, 163) <= input(5);
output(4, 164) <= input(6);
output(4, 165) <= input(7);
output(4, 166) <= input(8);
output(4, 167) <= input(9);
output(4, 168) <= input(10);
output(4, 169) <= input(11);
output(4, 170) <= input(12);
output(4, 171) <= input(13);
output(4, 172) <= input(14);
output(4, 173) <= input(15);
output(4, 174) <= input(32);
output(4, 175) <= input(34);
output(4, 176) <= input(18);
output(4, 177) <= input(19);
output(4, 178) <= input(20);
output(4, 179) <= input(21);
output(4, 180) <= input(22);
output(4, 181) <= input(23);
output(4, 182) <= input(24);
output(4, 183) <= input(25);
output(4, 184) <= input(26);
output(4, 185) <= input(27);
output(4, 186) <= input(28);
output(4, 187) <= input(29);
output(4, 188) <= input(30);
output(4, 189) <= input(31);
output(4, 190) <= input(33);
output(4, 191) <= input(35);
output(4, 192) <= input(18);
output(4, 193) <= input(19);
output(4, 194) <= input(20);
output(4, 195) <= input(21);
output(4, 196) <= input(22);
output(4, 197) <= input(23);
output(4, 198) <= input(24);
output(4, 199) <= input(25);
output(4, 200) <= input(26);
output(4, 201) <= input(27);
output(4, 202) <= input(28);
output(4, 203) <= input(29);
output(4, 204) <= input(30);
output(4, 205) <= input(31);
output(4, 206) <= input(33);
output(4, 207) <= input(35);
output(4, 208) <= input(3);
output(4, 209) <= input(4);
output(4, 210) <= input(5);
output(4, 211) <= input(6);
output(4, 212) <= input(7);
output(4, 213) <= input(8);
output(4, 214) <= input(9);
output(4, 215) <= input(10);
output(4, 216) <= input(11);
output(4, 217) <= input(12);
output(4, 218) <= input(13);
output(4, 219) <= input(14);
output(4, 220) <= input(15);
output(4, 221) <= input(32);
output(4, 222) <= input(34);
output(4, 223) <= input(36);
output(4, 224) <= input(3);
output(4, 225) <= input(4);
output(4, 226) <= input(5);
output(4, 227) <= input(6);
output(4, 228) <= input(7);
output(4, 229) <= input(8);
output(4, 230) <= input(9);
output(4, 231) <= input(10);
output(4, 232) <= input(11);
output(4, 233) <= input(12);
output(4, 234) <= input(13);
output(4, 235) <= input(14);
output(4, 236) <= input(15);
output(4, 237) <= input(32);
output(4, 238) <= input(34);
output(4, 239) <= input(36);
output(4, 240) <= input(19);
output(4, 241) <= input(20);
output(4, 242) <= input(21);
output(4, 243) <= input(22);
output(4, 244) <= input(23);
output(4, 245) <= input(24);
output(4, 246) <= input(25);
output(4, 247) <= input(26);
output(4, 248) <= input(27);
output(4, 249) <= input(28);
output(4, 250) <= input(29);
output(4, 251) <= input(30);
output(4, 252) <= input(31);
output(4, 253) <= input(33);
output(4, 254) <= input(35);
output(4, 255) <= input(37);
output(5, 0) <= input(46);
output(5, 1) <= input(16);
output(5, 2) <= input(17);
output(5, 3) <= input(18);
output(5, 4) <= input(19);
output(5, 5) <= input(20);
output(5, 6) <= input(21);
output(5, 7) <= input(22);
output(5, 8) <= input(23);
output(5, 9) <= input(24);
output(5, 10) <= input(25);
output(5, 11) <= input(26);
output(5, 12) <= input(27);
output(5, 13) <= input(28);
output(5, 14) <= input(29);
output(5, 15) <= input(30);
output(5, 16) <= input(46);
output(5, 17) <= input(16);
output(5, 18) <= input(17);
output(5, 19) <= input(18);
output(5, 20) <= input(19);
output(5, 21) <= input(20);
output(5, 22) <= input(21);
output(5, 23) <= input(22);
output(5, 24) <= input(23);
output(5, 25) <= input(24);
output(5, 26) <= input(25);
output(5, 27) <= input(26);
output(5, 28) <= input(27);
output(5, 29) <= input(28);
output(5, 30) <= input(29);
output(5, 31) <= input(30);
output(5, 32) <= input(0);
output(5, 33) <= input(1);
output(5, 34) <= input(2);
output(5, 35) <= input(3);
output(5, 36) <= input(4);
output(5, 37) <= input(5);
output(5, 38) <= input(6);
output(5, 39) <= input(7);
output(5, 40) <= input(8);
output(5, 41) <= input(9);
output(5, 42) <= input(10);
output(5, 43) <= input(11);
output(5, 44) <= input(12);
output(5, 45) <= input(13);
output(5, 46) <= input(14);
output(5, 47) <= input(15);
output(5, 48) <= input(0);
output(5, 49) <= input(1);
output(5, 50) <= input(2);
output(5, 51) <= input(3);
output(5, 52) <= input(4);
output(5, 53) <= input(5);
output(5, 54) <= input(6);
output(5, 55) <= input(7);
output(5, 56) <= input(8);
output(5, 57) <= input(9);
output(5, 58) <= input(10);
output(5, 59) <= input(11);
output(5, 60) <= input(12);
output(5, 61) <= input(13);
output(5, 62) <= input(14);
output(5, 63) <= input(15);
output(5, 64) <= input(0);
output(5, 65) <= input(1);
output(5, 66) <= input(2);
output(5, 67) <= input(3);
output(5, 68) <= input(4);
output(5, 69) <= input(5);
output(5, 70) <= input(6);
output(5, 71) <= input(7);
output(5, 72) <= input(8);
output(5, 73) <= input(9);
output(5, 74) <= input(10);
output(5, 75) <= input(11);
output(5, 76) <= input(12);
output(5, 77) <= input(13);
output(5, 78) <= input(14);
output(5, 79) <= input(15);
output(5, 80) <= input(16);
output(5, 81) <= input(17);
output(5, 82) <= input(18);
output(5, 83) <= input(19);
output(5, 84) <= input(20);
output(5, 85) <= input(21);
output(5, 86) <= input(22);
output(5, 87) <= input(23);
output(5, 88) <= input(24);
output(5, 89) <= input(25);
output(5, 90) <= input(26);
output(5, 91) <= input(27);
output(5, 92) <= input(28);
output(5, 93) <= input(29);
output(5, 94) <= input(30);
output(5, 95) <= input(31);
output(5, 96) <= input(16);
output(5, 97) <= input(17);
output(5, 98) <= input(18);
output(5, 99) <= input(19);
output(5, 100) <= input(20);
output(5, 101) <= input(21);
output(5, 102) <= input(22);
output(5, 103) <= input(23);
output(5, 104) <= input(24);
output(5, 105) <= input(25);
output(5, 106) <= input(26);
output(5, 107) <= input(27);
output(5, 108) <= input(28);
output(5, 109) <= input(29);
output(5, 110) <= input(30);
output(5, 111) <= input(31);
output(5, 112) <= input(1);
output(5, 113) <= input(2);
output(5, 114) <= input(3);
output(5, 115) <= input(4);
output(5, 116) <= input(5);
output(5, 117) <= input(6);
output(5, 118) <= input(7);
output(5, 119) <= input(8);
output(5, 120) <= input(9);
output(5, 121) <= input(10);
output(5, 122) <= input(11);
output(5, 123) <= input(12);
output(5, 124) <= input(13);
output(5, 125) <= input(14);
output(5, 126) <= input(15);
output(5, 127) <= input(32);
output(5, 128) <= input(1);
output(5, 129) <= input(2);
output(5, 130) <= input(3);
output(5, 131) <= input(4);
output(5, 132) <= input(5);
output(5, 133) <= input(6);
output(5, 134) <= input(7);
output(5, 135) <= input(8);
output(5, 136) <= input(9);
output(5, 137) <= input(10);
output(5, 138) <= input(11);
output(5, 139) <= input(12);
output(5, 140) <= input(13);
output(5, 141) <= input(14);
output(5, 142) <= input(15);
output(5, 143) <= input(32);
output(5, 144) <= input(1);
output(5, 145) <= input(2);
output(5, 146) <= input(3);
output(5, 147) <= input(4);
output(5, 148) <= input(5);
output(5, 149) <= input(6);
output(5, 150) <= input(7);
output(5, 151) <= input(8);
output(5, 152) <= input(9);
output(5, 153) <= input(10);
output(5, 154) <= input(11);
output(5, 155) <= input(12);
output(5, 156) <= input(13);
output(5, 157) <= input(14);
output(5, 158) <= input(15);
output(5, 159) <= input(32);
output(5, 160) <= input(17);
output(5, 161) <= input(18);
output(5, 162) <= input(19);
output(5, 163) <= input(20);
output(5, 164) <= input(21);
output(5, 165) <= input(22);
output(5, 166) <= input(23);
output(5, 167) <= input(24);
output(5, 168) <= input(25);
output(5, 169) <= input(26);
output(5, 170) <= input(27);
output(5, 171) <= input(28);
output(5, 172) <= input(29);
output(5, 173) <= input(30);
output(5, 174) <= input(31);
output(5, 175) <= input(33);
output(5, 176) <= input(17);
output(5, 177) <= input(18);
output(5, 178) <= input(19);
output(5, 179) <= input(20);
output(5, 180) <= input(21);
output(5, 181) <= input(22);
output(5, 182) <= input(23);
output(5, 183) <= input(24);
output(5, 184) <= input(25);
output(5, 185) <= input(26);
output(5, 186) <= input(27);
output(5, 187) <= input(28);
output(5, 188) <= input(29);
output(5, 189) <= input(30);
output(5, 190) <= input(31);
output(5, 191) <= input(33);
output(5, 192) <= input(17);
output(5, 193) <= input(18);
output(5, 194) <= input(19);
output(5, 195) <= input(20);
output(5, 196) <= input(21);
output(5, 197) <= input(22);
output(5, 198) <= input(23);
output(5, 199) <= input(24);
output(5, 200) <= input(25);
output(5, 201) <= input(26);
output(5, 202) <= input(27);
output(5, 203) <= input(28);
output(5, 204) <= input(29);
output(5, 205) <= input(30);
output(5, 206) <= input(31);
output(5, 207) <= input(33);
output(5, 208) <= input(2);
output(5, 209) <= input(3);
output(5, 210) <= input(4);
output(5, 211) <= input(5);
output(5, 212) <= input(6);
output(5, 213) <= input(7);
output(5, 214) <= input(8);
output(5, 215) <= input(9);
output(5, 216) <= input(10);
output(5, 217) <= input(11);
output(5, 218) <= input(12);
output(5, 219) <= input(13);
output(5, 220) <= input(14);
output(5, 221) <= input(15);
output(5, 222) <= input(32);
output(5, 223) <= input(34);
output(5, 224) <= input(2);
output(5, 225) <= input(3);
output(5, 226) <= input(4);
output(5, 227) <= input(5);
output(5, 228) <= input(6);
output(5, 229) <= input(7);
output(5, 230) <= input(8);
output(5, 231) <= input(9);
output(5, 232) <= input(10);
output(5, 233) <= input(11);
output(5, 234) <= input(12);
output(5, 235) <= input(13);
output(5, 236) <= input(14);
output(5, 237) <= input(15);
output(5, 238) <= input(32);
output(5, 239) <= input(34);
output(5, 240) <= input(18);
output(5, 241) <= input(19);
output(5, 242) <= input(20);
output(5, 243) <= input(21);
output(5, 244) <= input(22);
output(5, 245) <= input(23);
output(5, 246) <= input(24);
output(5, 247) <= input(25);
output(5, 248) <= input(26);
output(5, 249) <= input(27);
output(5, 250) <= input(28);
output(5, 251) <= input(29);
output(5, 252) <= input(30);
output(5, 253) <= input(31);
output(5, 254) <= input(33);
output(5, 255) <= input(35);
when "0010" =>
output(0, 0) <= input(0);
output(0, 1) <= input(1);
output(0, 2) <= input(2);
output(0, 3) <= input(3);
output(0, 4) <= input(4);
output(0, 5) <= input(5);
output(0, 6) <= input(6);
output(0, 7) <= input(7);
output(0, 8) <= input(8);
output(0, 9) <= input(9);
output(0, 10) <= input(10);
output(0, 11) <= input(11);
output(0, 12) <= input(12);
output(0, 13) <= input(13);
output(0, 14) <= input(14);
output(0, 15) <= input(15);
output(0, 16) <= input(0);
output(0, 17) <= input(1);
output(0, 18) <= input(2);
output(0, 19) <= input(3);
output(0, 20) <= input(4);
output(0, 21) <= input(5);
output(0, 22) <= input(6);
output(0, 23) <= input(7);
output(0, 24) <= input(8);
output(0, 25) <= input(9);
output(0, 26) <= input(10);
output(0, 27) <= input(11);
output(0, 28) <= input(12);
output(0, 29) <= input(13);
output(0, 30) <= input(14);
output(0, 31) <= input(15);
output(0, 32) <= input(0);
output(0, 33) <= input(1);
output(0, 34) <= input(2);
output(0, 35) <= input(3);
output(0, 36) <= input(4);
output(0, 37) <= input(5);
output(0, 38) <= input(6);
output(0, 39) <= input(7);
output(0, 40) <= input(8);
output(0, 41) <= input(9);
output(0, 42) <= input(10);
output(0, 43) <= input(11);
output(0, 44) <= input(12);
output(0, 45) <= input(13);
output(0, 46) <= input(14);
output(0, 47) <= input(15);
output(0, 48) <= input(16);
output(0, 49) <= input(17);
output(0, 50) <= input(18);
output(0, 51) <= input(19);
output(0, 52) <= input(20);
output(0, 53) <= input(21);
output(0, 54) <= input(22);
output(0, 55) <= input(23);
output(0, 56) <= input(24);
output(0, 57) <= input(25);
output(0, 58) <= input(26);
output(0, 59) <= input(27);
output(0, 60) <= input(28);
output(0, 61) <= input(29);
output(0, 62) <= input(30);
output(0, 63) <= input(31);
output(0, 64) <= input(16);
output(0, 65) <= input(17);
output(0, 66) <= input(18);
output(0, 67) <= input(19);
output(0, 68) <= input(20);
output(0, 69) <= input(21);
output(0, 70) <= input(22);
output(0, 71) <= input(23);
output(0, 72) <= input(24);
output(0, 73) <= input(25);
output(0, 74) <= input(26);
output(0, 75) <= input(27);
output(0, 76) <= input(28);
output(0, 77) <= input(29);
output(0, 78) <= input(30);
output(0, 79) <= input(31);
output(0, 80) <= input(16);
output(0, 81) <= input(17);
output(0, 82) <= input(18);
output(0, 83) <= input(19);
output(0, 84) <= input(20);
output(0, 85) <= input(21);
output(0, 86) <= input(22);
output(0, 87) <= input(23);
output(0, 88) <= input(24);
output(0, 89) <= input(25);
output(0, 90) <= input(26);
output(0, 91) <= input(27);
output(0, 92) <= input(28);
output(0, 93) <= input(29);
output(0, 94) <= input(30);
output(0, 95) <= input(31);
output(0, 96) <= input(16);
output(0, 97) <= input(17);
output(0, 98) <= input(18);
output(0, 99) <= input(19);
output(0, 100) <= input(20);
output(0, 101) <= input(21);
output(0, 102) <= input(22);
output(0, 103) <= input(23);
output(0, 104) <= input(24);
output(0, 105) <= input(25);
output(0, 106) <= input(26);
output(0, 107) <= input(27);
output(0, 108) <= input(28);
output(0, 109) <= input(29);
output(0, 110) <= input(30);
output(0, 111) <= input(31);
output(0, 112) <= input(1);
output(0, 113) <= input(2);
output(0, 114) <= input(3);
output(0, 115) <= input(4);
output(0, 116) <= input(5);
output(0, 117) <= input(6);
output(0, 118) <= input(7);
output(0, 119) <= input(8);
output(0, 120) <= input(9);
output(0, 121) <= input(10);
output(0, 122) <= input(11);
output(0, 123) <= input(12);
output(0, 124) <= input(13);
output(0, 125) <= input(14);
output(0, 126) <= input(15);
output(0, 127) <= input(32);
output(0, 128) <= input(1);
output(0, 129) <= input(2);
output(0, 130) <= input(3);
output(0, 131) <= input(4);
output(0, 132) <= input(5);
output(0, 133) <= input(6);
output(0, 134) <= input(7);
output(0, 135) <= input(8);
output(0, 136) <= input(9);
output(0, 137) <= input(10);
output(0, 138) <= input(11);
output(0, 139) <= input(12);
output(0, 140) <= input(13);
output(0, 141) <= input(14);
output(0, 142) <= input(15);
output(0, 143) <= input(32);
output(0, 144) <= input(1);
output(0, 145) <= input(2);
output(0, 146) <= input(3);
output(0, 147) <= input(4);
output(0, 148) <= input(5);
output(0, 149) <= input(6);
output(0, 150) <= input(7);
output(0, 151) <= input(8);
output(0, 152) <= input(9);
output(0, 153) <= input(10);
output(0, 154) <= input(11);
output(0, 155) <= input(12);
output(0, 156) <= input(13);
output(0, 157) <= input(14);
output(0, 158) <= input(15);
output(0, 159) <= input(32);
output(0, 160) <= input(1);
output(0, 161) <= input(2);
output(0, 162) <= input(3);
output(0, 163) <= input(4);
output(0, 164) <= input(5);
output(0, 165) <= input(6);
output(0, 166) <= input(7);
output(0, 167) <= input(8);
output(0, 168) <= input(9);
output(0, 169) <= input(10);
output(0, 170) <= input(11);
output(0, 171) <= input(12);
output(0, 172) <= input(13);
output(0, 173) <= input(14);
output(0, 174) <= input(15);
output(0, 175) <= input(32);
output(0, 176) <= input(17);
output(0, 177) <= input(18);
output(0, 178) <= input(19);
output(0, 179) <= input(20);
output(0, 180) <= input(21);
output(0, 181) <= input(22);
output(0, 182) <= input(23);
output(0, 183) <= input(24);
output(0, 184) <= input(25);
output(0, 185) <= input(26);
output(0, 186) <= input(27);
output(0, 187) <= input(28);
output(0, 188) <= input(29);
output(0, 189) <= input(30);
output(0, 190) <= input(31);
output(0, 191) <= input(33);
output(0, 192) <= input(17);
output(0, 193) <= input(18);
output(0, 194) <= input(19);
output(0, 195) <= input(20);
output(0, 196) <= input(21);
output(0, 197) <= input(22);
output(0, 198) <= input(23);
output(0, 199) <= input(24);
output(0, 200) <= input(25);
output(0, 201) <= input(26);
output(0, 202) <= input(27);
output(0, 203) <= input(28);
output(0, 204) <= input(29);
output(0, 205) <= input(30);
output(0, 206) <= input(31);
output(0, 207) <= input(33);
output(0, 208) <= input(17);
output(0, 209) <= input(18);
output(0, 210) <= input(19);
output(0, 211) <= input(20);
output(0, 212) <= input(21);
output(0, 213) <= input(22);
output(0, 214) <= input(23);
output(0, 215) <= input(24);
output(0, 216) <= input(25);
output(0, 217) <= input(26);
output(0, 218) <= input(27);
output(0, 219) <= input(28);
output(0, 220) <= input(29);
output(0, 221) <= input(30);
output(0, 222) <= input(31);
output(0, 223) <= input(33);
output(0, 224) <= input(17);
output(0, 225) <= input(18);
output(0, 226) <= input(19);
output(0, 227) <= input(20);
output(0, 228) <= input(21);
output(0, 229) <= input(22);
output(0, 230) <= input(23);
output(0, 231) <= input(24);
output(0, 232) <= input(25);
output(0, 233) <= input(26);
output(0, 234) <= input(27);
output(0, 235) <= input(28);
output(0, 236) <= input(29);
output(0, 237) <= input(30);
output(0, 238) <= input(31);
output(0, 239) <= input(33);
output(0, 240) <= input(2);
output(0, 241) <= input(3);
output(0, 242) <= input(4);
output(0, 243) <= input(5);
output(0, 244) <= input(6);
output(0, 245) <= input(7);
output(0, 246) <= input(8);
output(0, 247) <= input(9);
output(0, 248) <= input(10);
output(0, 249) <= input(11);
output(0, 250) <= input(12);
output(0, 251) <= input(13);
output(0, 252) <= input(14);
output(0, 253) <= input(15);
output(0, 254) <= input(32);
output(0, 255) <= input(34);
output(1, 0) <= input(0);
output(1, 1) <= input(1);
output(1, 2) <= input(2);
output(1, 3) <= input(3);
output(1, 4) <= input(4);
output(1, 5) <= input(5);
output(1, 6) <= input(6);
output(1, 7) <= input(7);
output(1, 8) <= input(8);
output(1, 9) <= input(9);
output(1, 10) <= input(10);
output(1, 11) <= input(11);
output(1, 12) <= input(12);
output(1, 13) <= input(13);
output(1, 14) <= input(14);
output(1, 15) <= input(15);
output(1, 16) <= input(0);
output(1, 17) <= input(1);
output(1, 18) <= input(2);
output(1, 19) <= input(3);
output(1, 20) <= input(4);
output(1, 21) <= input(5);
output(1, 22) <= input(6);
output(1, 23) <= input(7);
output(1, 24) <= input(8);
output(1, 25) <= input(9);
output(1, 26) <= input(10);
output(1, 27) <= input(11);
output(1, 28) <= input(12);
output(1, 29) <= input(13);
output(1, 30) <= input(14);
output(1, 31) <= input(15);
output(1, 32) <= input(0);
output(1, 33) <= input(1);
output(1, 34) <= input(2);
output(1, 35) <= input(3);
output(1, 36) <= input(4);
output(1, 37) <= input(5);
output(1, 38) <= input(6);
output(1, 39) <= input(7);
output(1, 40) <= input(8);
output(1, 41) <= input(9);
output(1, 42) <= input(10);
output(1, 43) <= input(11);
output(1, 44) <= input(12);
output(1, 45) <= input(13);
output(1, 46) <= input(14);
output(1, 47) <= input(15);
output(1, 48) <= input(0);
output(1, 49) <= input(1);
output(1, 50) <= input(2);
output(1, 51) <= input(3);
output(1, 52) <= input(4);
output(1, 53) <= input(5);
output(1, 54) <= input(6);
output(1, 55) <= input(7);
output(1, 56) <= input(8);
output(1, 57) <= input(9);
output(1, 58) <= input(10);
output(1, 59) <= input(11);
output(1, 60) <= input(12);
output(1, 61) <= input(13);
output(1, 62) <= input(14);
output(1, 63) <= input(15);
output(1, 64) <= input(0);
output(1, 65) <= input(1);
output(1, 66) <= input(2);
output(1, 67) <= input(3);
output(1, 68) <= input(4);
output(1, 69) <= input(5);
output(1, 70) <= input(6);
output(1, 71) <= input(7);
output(1, 72) <= input(8);
output(1, 73) <= input(9);
output(1, 74) <= input(10);
output(1, 75) <= input(11);
output(1, 76) <= input(12);
output(1, 77) <= input(13);
output(1, 78) <= input(14);
output(1, 79) <= input(15);
output(1, 80) <= input(16);
output(1, 81) <= input(17);
output(1, 82) <= input(18);
output(1, 83) <= input(19);
output(1, 84) <= input(20);
output(1, 85) <= input(21);
output(1, 86) <= input(22);
output(1, 87) <= input(23);
output(1, 88) <= input(24);
output(1, 89) <= input(25);
output(1, 90) <= input(26);
output(1, 91) <= input(27);
output(1, 92) <= input(28);
output(1, 93) <= input(29);
output(1, 94) <= input(30);
output(1, 95) <= input(31);
output(1, 96) <= input(16);
output(1, 97) <= input(17);
output(1, 98) <= input(18);
output(1, 99) <= input(19);
output(1, 100) <= input(20);
output(1, 101) <= input(21);
output(1, 102) <= input(22);
output(1, 103) <= input(23);
output(1, 104) <= input(24);
output(1, 105) <= input(25);
output(1, 106) <= input(26);
output(1, 107) <= input(27);
output(1, 108) <= input(28);
output(1, 109) <= input(29);
output(1, 110) <= input(30);
output(1, 111) <= input(31);
output(1, 112) <= input(16);
output(1, 113) <= input(17);
output(1, 114) <= input(18);
output(1, 115) <= input(19);
output(1, 116) <= input(20);
output(1, 117) <= input(21);
output(1, 118) <= input(22);
output(1, 119) <= input(23);
output(1, 120) <= input(24);
output(1, 121) <= input(25);
output(1, 122) <= input(26);
output(1, 123) <= input(27);
output(1, 124) <= input(28);
output(1, 125) <= input(29);
output(1, 126) <= input(30);
output(1, 127) <= input(31);
output(1, 128) <= input(16);
output(1, 129) <= input(17);
output(1, 130) <= input(18);
output(1, 131) <= input(19);
output(1, 132) <= input(20);
output(1, 133) <= input(21);
output(1, 134) <= input(22);
output(1, 135) <= input(23);
output(1, 136) <= input(24);
output(1, 137) <= input(25);
output(1, 138) <= input(26);
output(1, 139) <= input(27);
output(1, 140) <= input(28);
output(1, 141) <= input(29);
output(1, 142) <= input(30);
output(1, 143) <= input(31);
output(1, 144) <= input(16);
output(1, 145) <= input(17);
output(1, 146) <= input(18);
output(1, 147) <= input(19);
output(1, 148) <= input(20);
output(1, 149) <= input(21);
output(1, 150) <= input(22);
output(1, 151) <= input(23);
output(1, 152) <= input(24);
output(1, 153) <= input(25);
output(1, 154) <= input(26);
output(1, 155) <= input(27);
output(1, 156) <= input(28);
output(1, 157) <= input(29);
output(1, 158) <= input(30);
output(1, 159) <= input(31);
output(1, 160) <= input(1);
output(1, 161) <= input(2);
output(1, 162) <= input(3);
output(1, 163) <= input(4);
output(1, 164) <= input(5);
output(1, 165) <= input(6);
output(1, 166) <= input(7);
output(1, 167) <= input(8);
output(1, 168) <= input(9);
output(1, 169) <= input(10);
output(1, 170) <= input(11);
output(1, 171) <= input(12);
output(1, 172) <= input(13);
output(1, 173) <= input(14);
output(1, 174) <= input(15);
output(1, 175) <= input(32);
output(1, 176) <= input(1);
output(1, 177) <= input(2);
output(1, 178) <= input(3);
output(1, 179) <= input(4);
output(1, 180) <= input(5);
output(1, 181) <= input(6);
output(1, 182) <= input(7);
output(1, 183) <= input(8);
output(1, 184) <= input(9);
output(1, 185) <= input(10);
output(1, 186) <= input(11);
output(1, 187) <= input(12);
output(1, 188) <= input(13);
output(1, 189) <= input(14);
output(1, 190) <= input(15);
output(1, 191) <= input(32);
output(1, 192) <= input(1);
output(1, 193) <= input(2);
output(1, 194) <= input(3);
output(1, 195) <= input(4);
output(1, 196) <= input(5);
output(1, 197) <= input(6);
output(1, 198) <= input(7);
output(1, 199) <= input(8);
output(1, 200) <= input(9);
output(1, 201) <= input(10);
output(1, 202) <= input(11);
output(1, 203) <= input(12);
output(1, 204) <= input(13);
output(1, 205) <= input(14);
output(1, 206) <= input(15);
output(1, 207) <= input(32);
output(1, 208) <= input(1);
output(1, 209) <= input(2);
output(1, 210) <= input(3);
output(1, 211) <= input(4);
output(1, 212) <= input(5);
output(1, 213) <= input(6);
output(1, 214) <= input(7);
output(1, 215) <= input(8);
output(1, 216) <= input(9);
output(1, 217) <= input(10);
output(1, 218) <= input(11);
output(1, 219) <= input(12);
output(1, 220) <= input(13);
output(1, 221) <= input(14);
output(1, 222) <= input(15);
output(1, 223) <= input(32);
output(1, 224) <= input(1);
output(1, 225) <= input(2);
output(1, 226) <= input(3);
output(1, 227) <= input(4);
output(1, 228) <= input(5);
output(1, 229) <= input(6);
output(1, 230) <= input(7);
output(1, 231) <= input(8);
output(1, 232) <= input(9);
output(1, 233) <= input(10);
output(1, 234) <= input(11);
output(1, 235) <= input(12);
output(1, 236) <= input(13);
output(1, 237) <= input(14);
output(1, 238) <= input(15);
output(1, 239) <= input(32);
output(1, 240) <= input(17);
output(1, 241) <= input(18);
output(1, 242) <= input(19);
output(1, 243) <= input(20);
output(1, 244) <= input(21);
output(1, 245) <= input(22);
output(1, 246) <= input(23);
output(1, 247) <= input(24);
output(1, 248) <= input(25);
output(1, 249) <= input(26);
output(1, 250) <= input(27);
output(1, 251) <= input(28);
output(1, 252) <= input(29);
output(1, 253) <= input(30);
output(1, 254) <= input(31);
output(1, 255) <= input(33);
output(2, 0) <= input(0);
output(2, 1) <= input(1);
output(2, 2) <= input(2);
output(2, 3) <= input(3);
output(2, 4) <= input(4);
output(2, 5) <= input(5);
output(2, 6) <= input(6);
output(2, 7) <= input(7);
output(2, 8) <= input(8);
output(2, 9) <= input(9);
output(2, 10) <= input(10);
output(2, 11) <= input(11);
output(2, 12) <= input(12);
output(2, 13) <= input(13);
output(2, 14) <= input(14);
output(2, 15) <= input(15);
output(2, 16) <= input(0);
output(2, 17) <= input(1);
output(2, 18) <= input(2);
output(2, 19) <= input(3);
output(2, 20) <= input(4);
output(2, 21) <= input(5);
output(2, 22) <= input(6);
output(2, 23) <= input(7);
output(2, 24) <= input(8);
output(2, 25) <= input(9);
output(2, 26) <= input(10);
output(2, 27) <= input(11);
output(2, 28) <= input(12);
output(2, 29) <= input(13);
output(2, 30) <= input(14);
output(2, 31) <= input(15);
output(2, 32) <= input(0);
output(2, 33) <= input(1);
output(2, 34) <= input(2);
output(2, 35) <= input(3);
output(2, 36) <= input(4);
output(2, 37) <= input(5);
output(2, 38) <= input(6);
output(2, 39) <= input(7);
output(2, 40) <= input(8);
output(2, 41) <= input(9);
output(2, 42) <= input(10);
output(2, 43) <= input(11);
output(2, 44) <= input(12);
output(2, 45) <= input(13);
output(2, 46) <= input(14);
output(2, 47) <= input(15);
output(2, 48) <= input(0);
output(2, 49) <= input(1);
output(2, 50) <= input(2);
output(2, 51) <= input(3);
output(2, 52) <= input(4);
output(2, 53) <= input(5);
output(2, 54) <= input(6);
output(2, 55) <= input(7);
output(2, 56) <= input(8);
output(2, 57) <= input(9);
output(2, 58) <= input(10);
output(2, 59) <= input(11);
output(2, 60) <= input(12);
output(2, 61) <= input(13);
output(2, 62) <= input(14);
output(2, 63) <= input(15);
output(2, 64) <= input(0);
output(2, 65) <= input(1);
output(2, 66) <= input(2);
output(2, 67) <= input(3);
output(2, 68) <= input(4);
output(2, 69) <= input(5);
output(2, 70) <= input(6);
output(2, 71) <= input(7);
output(2, 72) <= input(8);
output(2, 73) <= input(9);
output(2, 74) <= input(10);
output(2, 75) <= input(11);
output(2, 76) <= input(12);
output(2, 77) <= input(13);
output(2, 78) <= input(14);
output(2, 79) <= input(15);
output(2, 80) <= input(0);
output(2, 81) <= input(1);
output(2, 82) <= input(2);
output(2, 83) <= input(3);
output(2, 84) <= input(4);
output(2, 85) <= input(5);
output(2, 86) <= input(6);
output(2, 87) <= input(7);
output(2, 88) <= input(8);
output(2, 89) <= input(9);
output(2, 90) <= input(10);
output(2, 91) <= input(11);
output(2, 92) <= input(12);
output(2, 93) <= input(13);
output(2, 94) <= input(14);
output(2, 95) <= input(15);
output(2, 96) <= input(0);
output(2, 97) <= input(1);
output(2, 98) <= input(2);
output(2, 99) <= input(3);
output(2, 100) <= input(4);
output(2, 101) <= input(5);
output(2, 102) <= input(6);
output(2, 103) <= input(7);
output(2, 104) <= input(8);
output(2, 105) <= input(9);
output(2, 106) <= input(10);
output(2, 107) <= input(11);
output(2, 108) <= input(12);
output(2, 109) <= input(13);
output(2, 110) <= input(14);
output(2, 111) <= input(15);
output(2, 112) <= input(16);
output(2, 113) <= input(17);
output(2, 114) <= input(18);
output(2, 115) <= input(19);
output(2, 116) <= input(20);
output(2, 117) <= input(21);
output(2, 118) <= input(22);
output(2, 119) <= input(23);
output(2, 120) <= input(24);
output(2, 121) <= input(25);
output(2, 122) <= input(26);
output(2, 123) <= input(27);
output(2, 124) <= input(28);
output(2, 125) <= input(29);
output(2, 126) <= input(30);
output(2, 127) <= input(31);
output(2, 128) <= input(16);
output(2, 129) <= input(17);
output(2, 130) <= input(18);
output(2, 131) <= input(19);
output(2, 132) <= input(20);
output(2, 133) <= input(21);
output(2, 134) <= input(22);
output(2, 135) <= input(23);
output(2, 136) <= input(24);
output(2, 137) <= input(25);
output(2, 138) <= input(26);
output(2, 139) <= input(27);
output(2, 140) <= input(28);
output(2, 141) <= input(29);
output(2, 142) <= input(30);
output(2, 143) <= input(31);
output(2, 144) <= input(16);
output(2, 145) <= input(17);
output(2, 146) <= input(18);
output(2, 147) <= input(19);
output(2, 148) <= input(20);
output(2, 149) <= input(21);
output(2, 150) <= input(22);
output(2, 151) <= input(23);
output(2, 152) <= input(24);
output(2, 153) <= input(25);
output(2, 154) <= input(26);
output(2, 155) <= input(27);
output(2, 156) <= input(28);
output(2, 157) <= input(29);
output(2, 158) <= input(30);
output(2, 159) <= input(31);
output(2, 160) <= input(16);
output(2, 161) <= input(17);
output(2, 162) <= input(18);
output(2, 163) <= input(19);
output(2, 164) <= input(20);
output(2, 165) <= input(21);
output(2, 166) <= input(22);
output(2, 167) <= input(23);
output(2, 168) <= input(24);
output(2, 169) <= input(25);
output(2, 170) <= input(26);
output(2, 171) <= input(27);
output(2, 172) <= input(28);
output(2, 173) <= input(29);
output(2, 174) <= input(30);
output(2, 175) <= input(31);
output(2, 176) <= input(16);
output(2, 177) <= input(17);
output(2, 178) <= input(18);
output(2, 179) <= input(19);
output(2, 180) <= input(20);
output(2, 181) <= input(21);
output(2, 182) <= input(22);
output(2, 183) <= input(23);
output(2, 184) <= input(24);
output(2, 185) <= input(25);
output(2, 186) <= input(26);
output(2, 187) <= input(27);
output(2, 188) <= input(28);
output(2, 189) <= input(29);
output(2, 190) <= input(30);
output(2, 191) <= input(31);
output(2, 192) <= input(16);
output(2, 193) <= input(17);
output(2, 194) <= input(18);
output(2, 195) <= input(19);
output(2, 196) <= input(20);
output(2, 197) <= input(21);
output(2, 198) <= input(22);
output(2, 199) <= input(23);
output(2, 200) <= input(24);
output(2, 201) <= input(25);
output(2, 202) <= input(26);
output(2, 203) <= input(27);
output(2, 204) <= input(28);
output(2, 205) <= input(29);
output(2, 206) <= input(30);
output(2, 207) <= input(31);
output(2, 208) <= input(16);
output(2, 209) <= input(17);
output(2, 210) <= input(18);
output(2, 211) <= input(19);
output(2, 212) <= input(20);
output(2, 213) <= input(21);
output(2, 214) <= input(22);
output(2, 215) <= input(23);
output(2, 216) <= input(24);
output(2, 217) <= input(25);
output(2, 218) <= input(26);
output(2, 219) <= input(27);
output(2, 220) <= input(28);
output(2, 221) <= input(29);
output(2, 222) <= input(30);
output(2, 223) <= input(31);
output(2, 224) <= input(16);
output(2, 225) <= input(17);
output(2, 226) <= input(18);
output(2, 227) <= input(19);
output(2, 228) <= input(20);
output(2, 229) <= input(21);
output(2, 230) <= input(22);
output(2, 231) <= input(23);
output(2, 232) <= input(24);
output(2, 233) <= input(25);
output(2, 234) <= input(26);
output(2, 235) <= input(27);
output(2, 236) <= input(28);
output(2, 237) <= input(29);
output(2, 238) <= input(30);
output(2, 239) <= input(31);
output(2, 240) <= input(1);
output(2, 241) <= input(2);
output(2, 242) <= input(3);
output(2, 243) <= input(4);
output(2, 244) <= input(5);
output(2, 245) <= input(6);
output(2, 246) <= input(7);
output(2, 247) <= input(8);
output(2, 248) <= input(9);
output(2, 249) <= input(10);
output(2, 250) <= input(11);
output(2, 251) <= input(12);
output(2, 252) <= input(13);
output(2, 253) <= input(14);
output(2, 254) <= input(15);
output(2, 255) <= input(32);
output(3, 0) <= input(0);
output(3, 1) <= input(1);
output(3, 2) <= input(2);
output(3, 3) <= input(3);
output(3, 4) <= input(4);
output(3, 5) <= input(5);
output(3, 6) <= input(6);
output(3, 7) <= input(7);
output(3, 8) <= input(8);
output(3, 9) <= input(9);
output(3, 10) <= input(10);
output(3, 11) <= input(11);
output(3, 12) <= input(12);
output(3, 13) <= input(13);
output(3, 14) <= input(14);
output(3, 15) <= input(15);
output(3, 16) <= input(0);
output(3, 17) <= input(1);
output(3, 18) <= input(2);
output(3, 19) <= input(3);
output(3, 20) <= input(4);
output(3, 21) <= input(5);
output(3, 22) <= input(6);
output(3, 23) <= input(7);
output(3, 24) <= input(8);
output(3, 25) <= input(9);
output(3, 26) <= input(10);
output(3, 27) <= input(11);
output(3, 28) <= input(12);
output(3, 29) <= input(13);
output(3, 30) <= input(14);
output(3, 31) <= input(15);
output(3, 32) <= input(0);
output(3, 33) <= input(1);
output(3, 34) <= input(2);
output(3, 35) <= input(3);
output(3, 36) <= input(4);
output(3, 37) <= input(5);
output(3, 38) <= input(6);
output(3, 39) <= input(7);
output(3, 40) <= input(8);
output(3, 41) <= input(9);
output(3, 42) <= input(10);
output(3, 43) <= input(11);
output(3, 44) <= input(12);
output(3, 45) <= input(13);
output(3, 46) <= input(14);
output(3, 47) <= input(15);
output(3, 48) <= input(0);
output(3, 49) <= input(1);
output(3, 50) <= input(2);
output(3, 51) <= input(3);
output(3, 52) <= input(4);
output(3, 53) <= input(5);
output(3, 54) <= input(6);
output(3, 55) <= input(7);
output(3, 56) <= input(8);
output(3, 57) <= input(9);
output(3, 58) <= input(10);
output(3, 59) <= input(11);
output(3, 60) <= input(12);
output(3, 61) <= input(13);
output(3, 62) <= input(14);
output(3, 63) <= input(15);
output(3, 64) <= input(0);
output(3, 65) <= input(1);
output(3, 66) <= input(2);
output(3, 67) <= input(3);
output(3, 68) <= input(4);
output(3, 69) <= input(5);
output(3, 70) <= input(6);
output(3, 71) <= input(7);
output(3, 72) <= input(8);
output(3, 73) <= input(9);
output(3, 74) <= input(10);
output(3, 75) <= input(11);
output(3, 76) <= input(12);
output(3, 77) <= input(13);
output(3, 78) <= input(14);
output(3, 79) <= input(15);
output(3, 80) <= input(0);
output(3, 81) <= input(1);
output(3, 82) <= input(2);
output(3, 83) <= input(3);
output(3, 84) <= input(4);
output(3, 85) <= input(5);
output(3, 86) <= input(6);
output(3, 87) <= input(7);
output(3, 88) <= input(8);
output(3, 89) <= input(9);
output(3, 90) <= input(10);
output(3, 91) <= input(11);
output(3, 92) <= input(12);
output(3, 93) <= input(13);
output(3, 94) <= input(14);
output(3, 95) <= input(15);
output(3, 96) <= input(0);
output(3, 97) <= input(1);
output(3, 98) <= input(2);
output(3, 99) <= input(3);
output(3, 100) <= input(4);
output(3, 101) <= input(5);
output(3, 102) <= input(6);
output(3, 103) <= input(7);
output(3, 104) <= input(8);
output(3, 105) <= input(9);
output(3, 106) <= input(10);
output(3, 107) <= input(11);
output(3, 108) <= input(12);
output(3, 109) <= input(13);
output(3, 110) <= input(14);
output(3, 111) <= input(15);
output(3, 112) <= input(0);
output(3, 113) <= input(1);
output(3, 114) <= input(2);
output(3, 115) <= input(3);
output(3, 116) <= input(4);
output(3, 117) <= input(5);
output(3, 118) <= input(6);
output(3, 119) <= input(7);
output(3, 120) <= input(8);
output(3, 121) <= input(9);
output(3, 122) <= input(10);
output(3, 123) <= input(11);
output(3, 124) <= input(12);
output(3, 125) <= input(13);
output(3, 126) <= input(14);
output(3, 127) <= input(15);
output(3, 128) <= input(0);
output(3, 129) <= input(1);
output(3, 130) <= input(2);
output(3, 131) <= input(3);
output(3, 132) <= input(4);
output(3, 133) <= input(5);
output(3, 134) <= input(6);
output(3, 135) <= input(7);
output(3, 136) <= input(8);
output(3, 137) <= input(9);
output(3, 138) <= input(10);
output(3, 139) <= input(11);
output(3, 140) <= input(12);
output(3, 141) <= input(13);
output(3, 142) <= input(14);
output(3, 143) <= input(15);
output(3, 144) <= input(0);
output(3, 145) <= input(1);
output(3, 146) <= input(2);
output(3, 147) <= input(3);
output(3, 148) <= input(4);
output(3, 149) <= input(5);
output(3, 150) <= input(6);
output(3, 151) <= input(7);
output(3, 152) <= input(8);
output(3, 153) <= input(9);
output(3, 154) <= input(10);
output(3, 155) <= input(11);
output(3, 156) <= input(12);
output(3, 157) <= input(13);
output(3, 158) <= input(14);
output(3, 159) <= input(15);
output(3, 160) <= input(0);
output(3, 161) <= input(1);
output(3, 162) <= input(2);
output(3, 163) <= input(3);
output(3, 164) <= input(4);
output(3, 165) <= input(5);
output(3, 166) <= input(6);
output(3, 167) <= input(7);
output(3, 168) <= input(8);
output(3, 169) <= input(9);
output(3, 170) <= input(10);
output(3, 171) <= input(11);
output(3, 172) <= input(12);
output(3, 173) <= input(13);
output(3, 174) <= input(14);
output(3, 175) <= input(15);
output(3, 176) <= input(0);
output(3, 177) <= input(1);
output(3, 178) <= input(2);
output(3, 179) <= input(3);
output(3, 180) <= input(4);
output(3, 181) <= input(5);
output(3, 182) <= input(6);
output(3, 183) <= input(7);
output(3, 184) <= input(8);
output(3, 185) <= input(9);
output(3, 186) <= input(10);
output(3, 187) <= input(11);
output(3, 188) <= input(12);
output(3, 189) <= input(13);
output(3, 190) <= input(14);
output(3, 191) <= input(15);
output(3, 192) <= input(0);
output(3, 193) <= input(1);
output(3, 194) <= input(2);
output(3, 195) <= input(3);
output(3, 196) <= input(4);
output(3, 197) <= input(5);
output(3, 198) <= input(6);
output(3, 199) <= input(7);
output(3, 200) <= input(8);
output(3, 201) <= input(9);
output(3, 202) <= input(10);
output(3, 203) <= input(11);
output(3, 204) <= input(12);
output(3, 205) <= input(13);
output(3, 206) <= input(14);
output(3, 207) <= input(15);
output(3, 208) <= input(0);
output(3, 209) <= input(1);
output(3, 210) <= input(2);
output(3, 211) <= input(3);
output(3, 212) <= input(4);
output(3, 213) <= input(5);
output(3, 214) <= input(6);
output(3, 215) <= input(7);
output(3, 216) <= input(8);
output(3, 217) <= input(9);
output(3, 218) <= input(10);
output(3, 219) <= input(11);
output(3, 220) <= input(12);
output(3, 221) <= input(13);
output(3, 222) <= input(14);
output(3, 223) <= input(15);
output(3, 224) <= input(0);
output(3, 225) <= input(1);
output(3, 226) <= input(2);
output(3, 227) <= input(3);
output(3, 228) <= input(4);
output(3, 229) <= input(5);
output(3, 230) <= input(6);
output(3, 231) <= input(7);
output(3, 232) <= input(8);
output(3, 233) <= input(9);
output(3, 234) <= input(10);
output(3, 235) <= input(11);
output(3, 236) <= input(12);
output(3, 237) <= input(13);
output(3, 238) <= input(14);
output(3, 239) <= input(15);
output(3, 240) <= input(16);
output(3, 241) <= input(17);
output(3, 242) <= input(18);
output(3, 243) <= input(19);
output(3, 244) <= input(20);
output(3, 245) <= input(21);
output(3, 246) <= input(22);
output(3, 247) <= input(23);
output(3, 248) <= input(24);
output(3, 249) <= input(25);
output(3, 250) <= input(26);
output(3, 251) <= input(27);
output(3, 252) <= input(28);
output(3, 253) <= input(29);
output(3, 254) <= input(30);
output(3, 255) <= input(31);
output(4, 0) <= input(0);
output(4, 1) <= input(1);
output(4, 2) <= input(2);
output(4, 3) <= input(3);
output(4, 4) <= input(4);
output(4, 5) <= input(5);
output(4, 6) <= input(6);
output(4, 7) <= input(7);
output(4, 8) <= input(8);
output(4, 9) <= input(9);
output(4, 10) <= input(10);
output(4, 11) <= input(11);
output(4, 12) <= input(12);
output(4, 13) <= input(13);
output(4, 14) <= input(14);
output(4, 15) <= input(15);
output(4, 16) <= input(0);
output(4, 17) <= input(1);
output(4, 18) <= input(2);
output(4, 19) <= input(3);
output(4, 20) <= input(4);
output(4, 21) <= input(5);
output(4, 22) <= input(6);
output(4, 23) <= input(7);
output(4, 24) <= input(8);
output(4, 25) <= input(9);
output(4, 26) <= input(10);
output(4, 27) <= input(11);
output(4, 28) <= input(12);
output(4, 29) <= input(13);
output(4, 30) <= input(14);
output(4, 31) <= input(15);
output(4, 32) <= input(0);
output(4, 33) <= input(1);
output(4, 34) <= input(2);
output(4, 35) <= input(3);
output(4, 36) <= input(4);
output(4, 37) <= input(5);
output(4, 38) <= input(6);
output(4, 39) <= input(7);
output(4, 40) <= input(8);
output(4, 41) <= input(9);
output(4, 42) <= input(10);
output(4, 43) <= input(11);
output(4, 44) <= input(12);
output(4, 45) <= input(13);
output(4, 46) <= input(14);
output(4, 47) <= input(15);
output(4, 48) <= input(0);
output(4, 49) <= input(1);
output(4, 50) <= input(2);
output(4, 51) <= input(3);
output(4, 52) <= input(4);
output(4, 53) <= input(5);
output(4, 54) <= input(6);
output(4, 55) <= input(7);
output(4, 56) <= input(8);
output(4, 57) <= input(9);
output(4, 58) <= input(10);
output(4, 59) <= input(11);
output(4, 60) <= input(12);
output(4, 61) <= input(13);
output(4, 62) <= input(14);
output(4, 63) <= input(15);
output(4, 64) <= input(0);
output(4, 65) <= input(1);
output(4, 66) <= input(2);
output(4, 67) <= input(3);
output(4, 68) <= input(4);
output(4, 69) <= input(5);
output(4, 70) <= input(6);
output(4, 71) <= input(7);
output(4, 72) <= input(8);
output(4, 73) <= input(9);
output(4, 74) <= input(10);
output(4, 75) <= input(11);
output(4, 76) <= input(12);
output(4, 77) <= input(13);
output(4, 78) <= input(14);
output(4, 79) <= input(15);
output(4, 80) <= input(0);
output(4, 81) <= input(1);
output(4, 82) <= input(2);
output(4, 83) <= input(3);
output(4, 84) <= input(4);
output(4, 85) <= input(5);
output(4, 86) <= input(6);
output(4, 87) <= input(7);
output(4, 88) <= input(8);
output(4, 89) <= input(9);
output(4, 90) <= input(10);
output(4, 91) <= input(11);
output(4, 92) <= input(12);
output(4, 93) <= input(13);
output(4, 94) <= input(14);
output(4, 95) <= input(15);
output(4, 96) <= input(0);
output(4, 97) <= input(1);
output(4, 98) <= input(2);
output(4, 99) <= input(3);
output(4, 100) <= input(4);
output(4, 101) <= input(5);
output(4, 102) <= input(6);
output(4, 103) <= input(7);
output(4, 104) <= input(8);
output(4, 105) <= input(9);
output(4, 106) <= input(10);
output(4, 107) <= input(11);
output(4, 108) <= input(12);
output(4, 109) <= input(13);
output(4, 110) <= input(14);
output(4, 111) <= input(15);
output(4, 112) <= input(0);
output(4, 113) <= input(1);
output(4, 114) <= input(2);
output(4, 115) <= input(3);
output(4, 116) <= input(4);
output(4, 117) <= input(5);
output(4, 118) <= input(6);
output(4, 119) <= input(7);
output(4, 120) <= input(8);
output(4, 121) <= input(9);
output(4, 122) <= input(10);
output(4, 123) <= input(11);
output(4, 124) <= input(12);
output(4, 125) <= input(13);
output(4, 126) <= input(14);
output(4, 127) <= input(15);
output(4, 128) <= input(0);
output(4, 129) <= input(1);
output(4, 130) <= input(2);
output(4, 131) <= input(3);
output(4, 132) <= input(4);
output(4, 133) <= input(5);
output(4, 134) <= input(6);
output(4, 135) <= input(7);
output(4, 136) <= input(8);
output(4, 137) <= input(9);
output(4, 138) <= input(10);
output(4, 139) <= input(11);
output(4, 140) <= input(12);
output(4, 141) <= input(13);
output(4, 142) <= input(14);
output(4, 143) <= input(15);
output(4, 144) <= input(0);
output(4, 145) <= input(1);
output(4, 146) <= input(2);
output(4, 147) <= input(3);
output(4, 148) <= input(4);
output(4, 149) <= input(5);
output(4, 150) <= input(6);
output(4, 151) <= input(7);
output(4, 152) <= input(8);
output(4, 153) <= input(9);
output(4, 154) <= input(10);
output(4, 155) <= input(11);
output(4, 156) <= input(12);
output(4, 157) <= input(13);
output(4, 158) <= input(14);
output(4, 159) <= input(15);
output(4, 160) <= input(0);
output(4, 161) <= input(1);
output(4, 162) <= input(2);
output(4, 163) <= input(3);
output(4, 164) <= input(4);
output(4, 165) <= input(5);
output(4, 166) <= input(6);
output(4, 167) <= input(7);
output(4, 168) <= input(8);
output(4, 169) <= input(9);
output(4, 170) <= input(10);
output(4, 171) <= input(11);
output(4, 172) <= input(12);
output(4, 173) <= input(13);
output(4, 174) <= input(14);
output(4, 175) <= input(15);
output(4, 176) <= input(0);
output(4, 177) <= input(1);
output(4, 178) <= input(2);
output(4, 179) <= input(3);
output(4, 180) <= input(4);
output(4, 181) <= input(5);
output(4, 182) <= input(6);
output(4, 183) <= input(7);
output(4, 184) <= input(8);
output(4, 185) <= input(9);
output(4, 186) <= input(10);
output(4, 187) <= input(11);
output(4, 188) <= input(12);
output(4, 189) <= input(13);
output(4, 190) <= input(14);
output(4, 191) <= input(15);
output(4, 192) <= input(0);
output(4, 193) <= input(1);
output(4, 194) <= input(2);
output(4, 195) <= input(3);
output(4, 196) <= input(4);
output(4, 197) <= input(5);
output(4, 198) <= input(6);
output(4, 199) <= input(7);
output(4, 200) <= input(8);
output(4, 201) <= input(9);
output(4, 202) <= input(10);
output(4, 203) <= input(11);
output(4, 204) <= input(12);
output(4, 205) <= input(13);
output(4, 206) <= input(14);
output(4, 207) <= input(15);
output(4, 208) <= input(0);
output(4, 209) <= input(1);
output(4, 210) <= input(2);
output(4, 211) <= input(3);
output(4, 212) <= input(4);
output(4, 213) <= input(5);
output(4, 214) <= input(6);
output(4, 215) <= input(7);
output(4, 216) <= input(8);
output(4, 217) <= input(9);
output(4, 218) <= input(10);
output(4, 219) <= input(11);
output(4, 220) <= input(12);
output(4, 221) <= input(13);
output(4, 222) <= input(14);
output(4, 223) <= input(15);
output(4, 224) <= input(0);
output(4, 225) <= input(1);
output(4, 226) <= input(2);
output(4, 227) <= input(3);
output(4, 228) <= input(4);
output(4, 229) <= input(5);
output(4, 230) <= input(6);
output(4, 231) <= input(7);
output(4, 232) <= input(8);
output(4, 233) <= input(9);
output(4, 234) <= input(10);
output(4, 235) <= input(11);
output(4, 236) <= input(12);
output(4, 237) <= input(13);
output(4, 238) <= input(14);
output(4, 239) <= input(15);
output(4, 240) <= input(0);
output(4, 241) <= input(1);
output(4, 242) <= input(2);
output(4, 243) <= input(3);
output(4, 244) <= input(4);
output(4, 245) <= input(5);
output(4, 246) <= input(6);
output(4, 247) <= input(7);
output(4, 248) <= input(8);
output(4, 249) <= input(9);
output(4, 250) <= input(10);
output(4, 251) <= input(11);
output(4, 252) <= input(12);
output(4, 253) <= input(13);
output(4, 254) <= input(14);
output(4, 255) <= input(15);
output(5, 0) <= input(35);
output(5, 1) <= input(16);
output(5, 2) <= input(17);
output(5, 3) <= input(18);
output(5, 4) <= input(19);
output(5, 5) <= input(20);
output(5, 6) <= input(21);
output(5, 7) <= input(22);
output(5, 8) <= input(23);
output(5, 9) <= input(24);
output(5, 10) <= input(25);
output(5, 11) <= input(26);
output(5, 12) <= input(27);
output(5, 13) <= input(28);
output(5, 14) <= input(29);
output(5, 15) <= input(30);
output(5, 16) <= input(35);
output(5, 17) <= input(16);
output(5, 18) <= input(17);
output(5, 19) <= input(18);
output(5, 20) <= input(19);
output(5, 21) <= input(20);
output(5, 22) <= input(21);
output(5, 23) <= input(22);
output(5, 24) <= input(23);
output(5, 25) <= input(24);
output(5, 26) <= input(25);
output(5, 27) <= input(26);
output(5, 28) <= input(27);
output(5, 29) <= input(28);
output(5, 30) <= input(29);
output(5, 31) <= input(30);
output(5, 32) <= input(35);
output(5, 33) <= input(16);
output(5, 34) <= input(17);
output(5, 35) <= input(18);
output(5, 36) <= input(19);
output(5, 37) <= input(20);
output(5, 38) <= input(21);
output(5, 39) <= input(22);
output(5, 40) <= input(23);
output(5, 41) <= input(24);
output(5, 42) <= input(25);
output(5, 43) <= input(26);
output(5, 44) <= input(27);
output(5, 45) <= input(28);
output(5, 46) <= input(29);
output(5, 47) <= input(30);
output(5, 48) <= input(35);
output(5, 49) <= input(16);
output(5, 50) <= input(17);
output(5, 51) <= input(18);
output(5, 52) <= input(19);
output(5, 53) <= input(20);
output(5, 54) <= input(21);
output(5, 55) <= input(22);
output(5, 56) <= input(23);
output(5, 57) <= input(24);
output(5, 58) <= input(25);
output(5, 59) <= input(26);
output(5, 60) <= input(27);
output(5, 61) <= input(28);
output(5, 62) <= input(29);
output(5, 63) <= input(30);
output(5, 64) <= input(35);
output(5, 65) <= input(16);
output(5, 66) <= input(17);
output(5, 67) <= input(18);
output(5, 68) <= input(19);
output(5, 69) <= input(20);
output(5, 70) <= input(21);
output(5, 71) <= input(22);
output(5, 72) <= input(23);
output(5, 73) <= input(24);
output(5, 74) <= input(25);
output(5, 75) <= input(26);
output(5, 76) <= input(27);
output(5, 77) <= input(28);
output(5, 78) <= input(29);
output(5, 79) <= input(30);
output(5, 80) <= input(35);
output(5, 81) <= input(16);
output(5, 82) <= input(17);
output(5, 83) <= input(18);
output(5, 84) <= input(19);
output(5, 85) <= input(20);
output(5, 86) <= input(21);
output(5, 87) <= input(22);
output(5, 88) <= input(23);
output(5, 89) <= input(24);
output(5, 90) <= input(25);
output(5, 91) <= input(26);
output(5, 92) <= input(27);
output(5, 93) <= input(28);
output(5, 94) <= input(29);
output(5, 95) <= input(30);
output(5, 96) <= input(35);
output(5, 97) <= input(16);
output(5, 98) <= input(17);
output(5, 99) <= input(18);
output(5, 100) <= input(19);
output(5, 101) <= input(20);
output(5, 102) <= input(21);
output(5, 103) <= input(22);
output(5, 104) <= input(23);
output(5, 105) <= input(24);
output(5, 106) <= input(25);
output(5, 107) <= input(26);
output(5, 108) <= input(27);
output(5, 109) <= input(28);
output(5, 110) <= input(29);
output(5, 111) <= input(30);
output(5, 112) <= input(35);
output(5, 113) <= input(16);
output(5, 114) <= input(17);
output(5, 115) <= input(18);
output(5, 116) <= input(19);
output(5, 117) <= input(20);
output(5, 118) <= input(21);
output(5, 119) <= input(22);
output(5, 120) <= input(23);
output(5, 121) <= input(24);
output(5, 122) <= input(25);
output(5, 123) <= input(26);
output(5, 124) <= input(27);
output(5, 125) <= input(28);
output(5, 126) <= input(29);
output(5, 127) <= input(30);
output(5, 128) <= input(35);
output(5, 129) <= input(16);
output(5, 130) <= input(17);
output(5, 131) <= input(18);
output(5, 132) <= input(19);
output(5, 133) <= input(20);
output(5, 134) <= input(21);
output(5, 135) <= input(22);
output(5, 136) <= input(23);
output(5, 137) <= input(24);
output(5, 138) <= input(25);
output(5, 139) <= input(26);
output(5, 140) <= input(27);
output(5, 141) <= input(28);
output(5, 142) <= input(29);
output(5, 143) <= input(30);
output(5, 144) <= input(35);
output(5, 145) <= input(16);
output(5, 146) <= input(17);
output(5, 147) <= input(18);
output(5, 148) <= input(19);
output(5, 149) <= input(20);
output(5, 150) <= input(21);
output(5, 151) <= input(22);
output(5, 152) <= input(23);
output(5, 153) <= input(24);
output(5, 154) <= input(25);
output(5, 155) <= input(26);
output(5, 156) <= input(27);
output(5, 157) <= input(28);
output(5, 158) <= input(29);
output(5, 159) <= input(30);
output(5, 160) <= input(35);
output(5, 161) <= input(16);
output(5, 162) <= input(17);
output(5, 163) <= input(18);
output(5, 164) <= input(19);
output(5, 165) <= input(20);
output(5, 166) <= input(21);
output(5, 167) <= input(22);
output(5, 168) <= input(23);
output(5, 169) <= input(24);
output(5, 170) <= input(25);
output(5, 171) <= input(26);
output(5, 172) <= input(27);
output(5, 173) <= input(28);
output(5, 174) <= input(29);
output(5, 175) <= input(30);
output(5, 176) <= input(35);
output(5, 177) <= input(16);
output(5, 178) <= input(17);
output(5, 179) <= input(18);
output(5, 180) <= input(19);
output(5, 181) <= input(20);
output(5, 182) <= input(21);
output(5, 183) <= input(22);
output(5, 184) <= input(23);
output(5, 185) <= input(24);
output(5, 186) <= input(25);
output(5, 187) <= input(26);
output(5, 188) <= input(27);
output(5, 189) <= input(28);
output(5, 190) <= input(29);
output(5, 191) <= input(30);
output(5, 192) <= input(35);
output(5, 193) <= input(16);
output(5, 194) <= input(17);
output(5, 195) <= input(18);
output(5, 196) <= input(19);
output(5, 197) <= input(20);
output(5, 198) <= input(21);
output(5, 199) <= input(22);
output(5, 200) <= input(23);
output(5, 201) <= input(24);
output(5, 202) <= input(25);
output(5, 203) <= input(26);
output(5, 204) <= input(27);
output(5, 205) <= input(28);
output(5, 206) <= input(29);
output(5, 207) <= input(30);
output(5, 208) <= input(35);
output(5, 209) <= input(16);
output(5, 210) <= input(17);
output(5, 211) <= input(18);
output(5, 212) <= input(19);
output(5, 213) <= input(20);
output(5, 214) <= input(21);
output(5, 215) <= input(22);
output(5, 216) <= input(23);
output(5, 217) <= input(24);
output(5, 218) <= input(25);
output(5, 219) <= input(26);
output(5, 220) <= input(27);
output(5, 221) <= input(28);
output(5, 222) <= input(29);
output(5, 223) <= input(30);
output(5, 224) <= input(35);
output(5, 225) <= input(16);
output(5, 226) <= input(17);
output(5, 227) <= input(18);
output(5, 228) <= input(19);
output(5, 229) <= input(20);
output(5, 230) <= input(21);
output(5, 231) <= input(22);
output(5, 232) <= input(23);
output(5, 233) <= input(24);
output(5, 234) <= input(25);
output(5, 235) <= input(26);
output(5, 236) <= input(27);
output(5, 237) <= input(28);
output(5, 238) <= input(29);
output(5, 239) <= input(30);
output(5, 240) <= input(35);
output(5, 241) <= input(16);
output(5, 242) <= input(17);
output(5, 243) <= input(18);
output(5, 244) <= input(19);
output(5, 245) <= input(20);
output(5, 246) <= input(21);
output(5, 247) <= input(22);
output(5, 248) <= input(23);
output(5, 249) <= input(24);
output(5, 250) <= input(25);
output(5, 251) <= input(26);
output(5, 252) <= input(27);
output(5, 253) <= input(28);
output(5, 254) <= input(29);
output(5, 255) <= input(30);
output(6, 0) <= input(35);
output(6, 1) <= input(16);
output(6, 2) <= input(17);
output(6, 3) <= input(18);
output(6, 4) <= input(19);
output(6, 5) <= input(20);
output(6, 6) <= input(21);
output(6, 7) <= input(22);
output(6, 8) <= input(23);
output(6, 9) <= input(24);
output(6, 10) <= input(25);
output(6, 11) <= input(26);
output(6, 12) <= input(27);
output(6, 13) <= input(28);
output(6, 14) <= input(29);
output(6, 15) <= input(30);
output(6, 16) <= input(35);
output(6, 17) <= input(16);
output(6, 18) <= input(17);
output(6, 19) <= input(18);
output(6, 20) <= input(19);
output(6, 21) <= input(20);
output(6, 22) <= input(21);
output(6, 23) <= input(22);
output(6, 24) <= input(23);
output(6, 25) <= input(24);
output(6, 26) <= input(25);
output(6, 27) <= input(26);
output(6, 28) <= input(27);
output(6, 29) <= input(28);
output(6, 30) <= input(29);
output(6, 31) <= input(30);
output(6, 32) <= input(35);
output(6, 33) <= input(16);
output(6, 34) <= input(17);
output(6, 35) <= input(18);
output(6, 36) <= input(19);
output(6, 37) <= input(20);
output(6, 38) <= input(21);
output(6, 39) <= input(22);
output(6, 40) <= input(23);
output(6, 41) <= input(24);
output(6, 42) <= input(25);
output(6, 43) <= input(26);
output(6, 44) <= input(27);
output(6, 45) <= input(28);
output(6, 46) <= input(29);
output(6, 47) <= input(30);
output(6, 48) <= input(35);
output(6, 49) <= input(16);
output(6, 50) <= input(17);
output(6, 51) <= input(18);
output(6, 52) <= input(19);
output(6, 53) <= input(20);
output(6, 54) <= input(21);
output(6, 55) <= input(22);
output(6, 56) <= input(23);
output(6, 57) <= input(24);
output(6, 58) <= input(25);
output(6, 59) <= input(26);
output(6, 60) <= input(27);
output(6, 61) <= input(28);
output(6, 62) <= input(29);
output(6, 63) <= input(30);
output(6, 64) <= input(35);
output(6, 65) <= input(16);
output(6, 66) <= input(17);
output(6, 67) <= input(18);
output(6, 68) <= input(19);
output(6, 69) <= input(20);
output(6, 70) <= input(21);
output(6, 71) <= input(22);
output(6, 72) <= input(23);
output(6, 73) <= input(24);
output(6, 74) <= input(25);
output(6, 75) <= input(26);
output(6, 76) <= input(27);
output(6, 77) <= input(28);
output(6, 78) <= input(29);
output(6, 79) <= input(30);
output(6, 80) <= input(35);
output(6, 81) <= input(16);
output(6, 82) <= input(17);
output(6, 83) <= input(18);
output(6, 84) <= input(19);
output(6, 85) <= input(20);
output(6, 86) <= input(21);
output(6, 87) <= input(22);
output(6, 88) <= input(23);
output(6, 89) <= input(24);
output(6, 90) <= input(25);
output(6, 91) <= input(26);
output(6, 92) <= input(27);
output(6, 93) <= input(28);
output(6, 94) <= input(29);
output(6, 95) <= input(30);
output(6, 96) <= input(35);
output(6, 97) <= input(16);
output(6, 98) <= input(17);
output(6, 99) <= input(18);
output(6, 100) <= input(19);
output(6, 101) <= input(20);
output(6, 102) <= input(21);
output(6, 103) <= input(22);
output(6, 104) <= input(23);
output(6, 105) <= input(24);
output(6, 106) <= input(25);
output(6, 107) <= input(26);
output(6, 108) <= input(27);
output(6, 109) <= input(28);
output(6, 110) <= input(29);
output(6, 111) <= input(30);
output(6, 112) <= input(35);
output(6, 113) <= input(16);
output(6, 114) <= input(17);
output(6, 115) <= input(18);
output(6, 116) <= input(19);
output(6, 117) <= input(20);
output(6, 118) <= input(21);
output(6, 119) <= input(22);
output(6, 120) <= input(23);
output(6, 121) <= input(24);
output(6, 122) <= input(25);
output(6, 123) <= input(26);
output(6, 124) <= input(27);
output(6, 125) <= input(28);
output(6, 126) <= input(29);
output(6, 127) <= input(30);
output(6, 128) <= input(36);
output(6, 129) <= input(0);
output(6, 130) <= input(1);
output(6, 131) <= input(2);
output(6, 132) <= input(3);
output(6, 133) <= input(4);
output(6, 134) <= input(5);
output(6, 135) <= input(6);
output(6, 136) <= input(7);
output(6, 137) <= input(8);
output(6, 138) <= input(9);
output(6, 139) <= input(10);
output(6, 140) <= input(11);
output(6, 141) <= input(12);
output(6, 142) <= input(13);
output(6, 143) <= input(14);
output(6, 144) <= input(36);
output(6, 145) <= input(0);
output(6, 146) <= input(1);
output(6, 147) <= input(2);
output(6, 148) <= input(3);
output(6, 149) <= input(4);
output(6, 150) <= input(5);
output(6, 151) <= input(6);
output(6, 152) <= input(7);
output(6, 153) <= input(8);
output(6, 154) <= input(9);
output(6, 155) <= input(10);
output(6, 156) <= input(11);
output(6, 157) <= input(12);
output(6, 158) <= input(13);
output(6, 159) <= input(14);
output(6, 160) <= input(36);
output(6, 161) <= input(0);
output(6, 162) <= input(1);
output(6, 163) <= input(2);
output(6, 164) <= input(3);
output(6, 165) <= input(4);
output(6, 166) <= input(5);
output(6, 167) <= input(6);
output(6, 168) <= input(7);
output(6, 169) <= input(8);
output(6, 170) <= input(9);
output(6, 171) <= input(10);
output(6, 172) <= input(11);
output(6, 173) <= input(12);
output(6, 174) <= input(13);
output(6, 175) <= input(14);
output(6, 176) <= input(36);
output(6, 177) <= input(0);
output(6, 178) <= input(1);
output(6, 179) <= input(2);
output(6, 180) <= input(3);
output(6, 181) <= input(4);
output(6, 182) <= input(5);
output(6, 183) <= input(6);
output(6, 184) <= input(7);
output(6, 185) <= input(8);
output(6, 186) <= input(9);
output(6, 187) <= input(10);
output(6, 188) <= input(11);
output(6, 189) <= input(12);
output(6, 190) <= input(13);
output(6, 191) <= input(14);
output(6, 192) <= input(36);
output(6, 193) <= input(0);
output(6, 194) <= input(1);
output(6, 195) <= input(2);
output(6, 196) <= input(3);
output(6, 197) <= input(4);
output(6, 198) <= input(5);
output(6, 199) <= input(6);
output(6, 200) <= input(7);
output(6, 201) <= input(8);
output(6, 202) <= input(9);
output(6, 203) <= input(10);
output(6, 204) <= input(11);
output(6, 205) <= input(12);
output(6, 206) <= input(13);
output(6, 207) <= input(14);
output(6, 208) <= input(36);
output(6, 209) <= input(0);
output(6, 210) <= input(1);
output(6, 211) <= input(2);
output(6, 212) <= input(3);
output(6, 213) <= input(4);
output(6, 214) <= input(5);
output(6, 215) <= input(6);
output(6, 216) <= input(7);
output(6, 217) <= input(8);
output(6, 218) <= input(9);
output(6, 219) <= input(10);
output(6, 220) <= input(11);
output(6, 221) <= input(12);
output(6, 222) <= input(13);
output(6, 223) <= input(14);
output(6, 224) <= input(36);
output(6, 225) <= input(0);
output(6, 226) <= input(1);
output(6, 227) <= input(2);
output(6, 228) <= input(3);
output(6, 229) <= input(4);
output(6, 230) <= input(5);
output(6, 231) <= input(6);
output(6, 232) <= input(7);
output(6, 233) <= input(8);
output(6, 234) <= input(9);
output(6, 235) <= input(10);
output(6, 236) <= input(11);
output(6, 237) <= input(12);
output(6, 238) <= input(13);
output(6, 239) <= input(14);
output(6, 240) <= input(36);
output(6, 241) <= input(0);
output(6, 242) <= input(1);
output(6, 243) <= input(2);
output(6, 244) <= input(3);
output(6, 245) <= input(4);
output(6, 246) <= input(5);
output(6, 247) <= input(6);
output(6, 248) <= input(7);
output(6, 249) <= input(8);
output(6, 250) <= input(9);
output(6, 251) <= input(10);
output(6, 252) <= input(11);
output(6, 253) <= input(12);
output(6, 254) <= input(13);
output(6, 255) <= input(14);
output(7, 0) <= input(35);
output(7, 1) <= input(16);
output(7, 2) <= input(17);
output(7, 3) <= input(18);
output(7, 4) <= input(19);
output(7, 5) <= input(20);
output(7, 6) <= input(21);
output(7, 7) <= input(22);
output(7, 8) <= input(23);
output(7, 9) <= input(24);
output(7, 10) <= input(25);
output(7, 11) <= input(26);
output(7, 12) <= input(27);
output(7, 13) <= input(28);
output(7, 14) <= input(29);
output(7, 15) <= input(30);
output(7, 16) <= input(35);
output(7, 17) <= input(16);
output(7, 18) <= input(17);
output(7, 19) <= input(18);
output(7, 20) <= input(19);
output(7, 21) <= input(20);
output(7, 22) <= input(21);
output(7, 23) <= input(22);
output(7, 24) <= input(23);
output(7, 25) <= input(24);
output(7, 26) <= input(25);
output(7, 27) <= input(26);
output(7, 28) <= input(27);
output(7, 29) <= input(28);
output(7, 30) <= input(29);
output(7, 31) <= input(30);
output(7, 32) <= input(35);
output(7, 33) <= input(16);
output(7, 34) <= input(17);
output(7, 35) <= input(18);
output(7, 36) <= input(19);
output(7, 37) <= input(20);
output(7, 38) <= input(21);
output(7, 39) <= input(22);
output(7, 40) <= input(23);
output(7, 41) <= input(24);
output(7, 42) <= input(25);
output(7, 43) <= input(26);
output(7, 44) <= input(27);
output(7, 45) <= input(28);
output(7, 46) <= input(29);
output(7, 47) <= input(30);
output(7, 48) <= input(35);
output(7, 49) <= input(16);
output(7, 50) <= input(17);
output(7, 51) <= input(18);
output(7, 52) <= input(19);
output(7, 53) <= input(20);
output(7, 54) <= input(21);
output(7, 55) <= input(22);
output(7, 56) <= input(23);
output(7, 57) <= input(24);
output(7, 58) <= input(25);
output(7, 59) <= input(26);
output(7, 60) <= input(27);
output(7, 61) <= input(28);
output(7, 62) <= input(29);
output(7, 63) <= input(30);
output(7, 64) <= input(35);
output(7, 65) <= input(16);
output(7, 66) <= input(17);
output(7, 67) <= input(18);
output(7, 68) <= input(19);
output(7, 69) <= input(20);
output(7, 70) <= input(21);
output(7, 71) <= input(22);
output(7, 72) <= input(23);
output(7, 73) <= input(24);
output(7, 74) <= input(25);
output(7, 75) <= input(26);
output(7, 76) <= input(27);
output(7, 77) <= input(28);
output(7, 78) <= input(29);
output(7, 79) <= input(30);
output(7, 80) <= input(36);
output(7, 81) <= input(0);
output(7, 82) <= input(1);
output(7, 83) <= input(2);
output(7, 84) <= input(3);
output(7, 85) <= input(4);
output(7, 86) <= input(5);
output(7, 87) <= input(6);
output(7, 88) <= input(7);
output(7, 89) <= input(8);
output(7, 90) <= input(9);
output(7, 91) <= input(10);
output(7, 92) <= input(11);
output(7, 93) <= input(12);
output(7, 94) <= input(13);
output(7, 95) <= input(14);
output(7, 96) <= input(36);
output(7, 97) <= input(0);
output(7, 98) <= input(1);
output(7, 99) <= input(2);
output(7, 100) <= input(3);
output(7, 101) <= input(4);
output(7, 102) <= input(5);
output(7, 103) <= input(6);
output(7, 104) <= input(7);
output(7, 105) <= input(8);
output(7, 106) <= input(9);
output(7, 107) <= input(10);
output(7, 108) <= input(11);
output(7, 109) <= input(12);
output(7, 110) <= input(13);
output(7, 111) <= input(14);
output(7, 112) <= input(36);
output(7, 113) <= input(0);
output(7, 114) <= input(1);
output(7, 115) <= input(2);
output(7, 116) <= input(3);
output(7, 117) <= input(4);
output(7, 118) <= input(5);
output(7, 119) <= input(6);
output(7, 120) <= input(7);
output(7, 121) <= input(8);
output(7, 122) <= input(9);
output(7, 123) <= input(10);
output(7, 124) <= input(11);
output(7, 125) <= input(12);
output(7, 126) <= input(13);
output(7, 127) <= input(14);
output(7, 128) <= input(36);
output(7, 129) <= input(0);
output(7, 130) <= input(1);
output(7, 131) <= input(2);
output(7, 132) <= input(3);
output(7, 133) <= input(4);
output(7, 134) <= input(5);
output(7, 135) <= input(6);
output(7, 136) <= input(7);
output(7, 137) <= input(8);
output(7, 138) <= input(9);
output(7, 139) <= input(10);
output(7, 140) <= input(11);
output(7, 141) <= input(12);
output(7, 142) <= input(13);
output(7, 143) <= input(14);
output(7, 144) <= input(36);
output(7, 145) <= input(0);
output(7, 146) <= input(1);
output(7, 147) <= input(2);
output(7, 148) <= input(3);
output(7, 149) <= input(4);
output(7, 150) <= input(5);
output(7, 151) <= input(6);
output(7, 152) <= input(7);
output(7, 153) <= input(8);
output(7, 154) <= input(9);
output(7, 155) <= input(10);
output(7, 156) <= input(11);
output(7, 157) <= input(12);
output(7, 158) <= input(13);
output(7, 159) <= input(14);
output(7, 160) <= input(37);
output(7, 161) <= input(35);
output(7, 162) <= input(16);
output(7, 163) <= input(17);
output(7, 164) <= input(18);
output(7, 165) <= input(19);
output(7, 166) <= input(20);
output(7, 167) <= input(21);
output(7, 168) <= input(22);
output(7, 169) <= input(23);
output(7, 170) <= input(24);
output(7, 171) <= input(25);
output(7, 172) <= input(26);
output(7, 173) <= input(27);
output(7, 174) <= input(28);
output(7, 175) <= input(29);
output(7, 176) <= input(37);
output(7, 177) <= input(35);
output(7, 178) <= input(16);
output(7, 179) <= input(17);
output(7, 180) <= input(18);
output(7, 181) <= input(19);
output(7, 182) <= input(20);
output(7, 183) <= input(21);
output(7, 184) <= input(22);
output(7, 185) <= input(23);
output(7, 186) <= input(24);
output(7, 187) <= input(25);
output(7, 188) <= input(26);
output(7, 189) <= input(27);
output(7, 190) <= input(28);
output(7, 191) <= input(29);
output(7, 192) <= input(37);
output(7, 193) <= input(35);
output(7, 194) <= input(16);
output(7, 195) <= input(17);
output(7, 196) <= input(18);
output(7, 197) <= input(19);
output(7, 198) <= input(20);
output(7, 199) <= input(21);
output(7, 200) <= input(22);
output(7, 201) <= input(23);
output(7, 202) <= input(24);
output(7, 203) <= input(25);
output(7, 204) <= input(26);
output(7, 205) <= input(27);
output(7, 206) <= input(28);
output(7, 207) <= input(29);
output(7, 208) <= input(37);
output(7, 209) <= input(35);
output(7, 210) <= input(16);
output(7, 211) <= input(17);
output(7, 212) <= input(18);
output(7, 213) <= input(19);
output(7, 214) <= input(20);
output(7, 215) <= input(21);
output(7, 216) <= input(22);
output(7, 217) <= input(23);
output(7, 218) <= input(24);
output(7, 219) <= input(25);
output(7, 220) <= input(26);
output(7, 221) <= input(27);
output(7, 222) <= input(28);
output(7, 223) <= input(29);
output(7, 224) <= input(37);
output(7, 225) <= input(35);
output(7, 226) <= input(16);
output(7, 227) <= input(17);
output(7, 228) <= input(18);
output(7, 229) <= input(19);
output(7, 230) <= input(20);
output(7, 231) <= input(21);
output(7, 232) <= input(22);
output(7, 233) <= input(23);
output(7, 234) <= input(24);
output(7, 235) <= input(25);
output(7, 236) <= input(26);
output(7, 237) <= input(27);
output(7, 238) <= input(28);
output(7, 239) <= input(29);
output(7, 240) <= input(37);
output(7, 241) <= input(35);
output(7, 242) <= input(16);
output(7, 243) <= input(17);
output(7, 244) <= input(18);
output(7, 245) <= input(19);
output(7, 246) <= input(20);
output(7, 247) <= input(21);
output(7, 248) <= input(22);
output(7, 249) <= input(23);
output(7, 250) <= input(24);
output(7, 251) <= input(25);
output(7, 252) <= input(26);
output(7, 253) <= input(27);
output(7, 254) <= input(28);
output(7, 255) <= input(29);
when "0011" =>
output(0, 0) <= input(0);
output(0, 1) <= input(1);
output(0, 2) <= input(2);
output(0, 3) <= input(3);
output(0, 4) <= input(4);
output(0, 5) <= input(5);
output(0, 6) <= input(6);
output(0, 7) <= input(7);
output(0, 8) <= input(8);
output(0, 9) <= input(9);
output(0, 10) <= input(10);
output(0, 11) <= input(11);
output(0, 12) <= input(12);
output(0, 13) <= input(13);
output(0, 14) <= input(14);
output(0, 15) <= input(15);
output(0, 16) <= input(0);
output(0, 17) <= input(1);
output(0, 18) <= input(2);
output(0, 19) <= input(3);
output(0, 20) <= input(4);
output(0, 21) <= input(5);
output(0, 22) <= input(6);
output(0, 23) <= input(7);
output(0, 24) <= input(8);
output(0, 25) <= input(9);
output(0, 26) <= input(10);
output(0, 27) <= input(11);
output(0, 28) <= input(12);
output(0, 29) <= input(13);
output(0, 30) <= input(14);
output(0, 31) <= input(15);
output(0, 32) <= input(0);
output(0, 33) <= input(1);
output(0, 34) <= input(2);
output(0, 35) <= input(3);
output(0, 36) <= input(4);
output(0, 37) <= input(5);
output(0, 38) <= input(6);
output(0, 39) <= input(7);
output(0, 40) <= input(8);
output(0, 41) <= input(9);
output(0, 42) <= input(10);
output(0, 43) <= input(11);
output(0, 44) <= input(12);
output(0, 45) <= input(13);
output(0, 46) <= input(14);
output(0, 47) <= input(15);
output(0, 48) <= input(0);
output(0, 49) <= input(1);
output(0, 50) <= input(2);
output(0, 51) <= input(3);
output(0, 52) <= input(4);
output(0, 53) <= input(5);
output(0, 54) <= input(6);
output(0, 55) <= input(7);
output(0, 56) <= input(8);
output(0, 57) <= input(9);
output(0, 58) <= input(10);
output(0, 59) <= input(11);
output(0, 60) <= input(12);
output(0, 61) <= input(13);
output(0, 62) <= input(14);
output(0, 63) <= input(15);
output(0, 64) <= input(16);
output(0, 65) <= input(17);
output(0, 66) <= input(18);
output(0, 67) <= input(19);
output(0, 68) <= input(20);
output(0, 69) <= input(21);
output(0, 70) <= input(22);
output(0, 71) <= input(23);
output(0, 72) <= input(24);
output(0, 73) <= input(25);
output(0, 74) <= input(26);
output(0, 75) <= input(27);
output(0, 76) <= input(28);
output(0, 77) <= input(29);
output(0, 78) <= input(30);
output(0, 79) <= input(31);
output(0, 80) <= input(16);
output(0, 81) <= input(17);
output(0, 82) <= input(18);
output(0, 83) <= input(19);
output(0, 84) <= input(20);
output(0, 85) <= input(21);
output(0, 86) <= input(22);
output(0, 87) <= input(23);
output(0, 88) <= input(24);
output(0, 89) <= input(25);
output(0, 90) <= input(26);
output(0, 91) <= input(27);
output(0, 92) <= input(28);
output(0, 93) <= input(29);
output(0, 94) <= input(30);
output(0, 95) <= input(31);
output(0, 96) <= input(16);
output(0, 97) <= input(17);
output(0, 98) <= input(18);
output(0, 99) <= input(19);
output(0, 100) <= input(20);
output(0, 101) <= input(21);
output(0, 102) <= input(22);
output(0, 103) <= input(23);
output(0, 104) <= input(24);
output(0, 105) <= input(25);
output(0, 106) <= input(26);
output(0, 107) <= input(27);
output(0, 108) <= input(28);
output(0, 109) <= input(29);
output(0, 110) <= input(30);
output(0, 111) <= input(31);
output(0, 112) <= input(16);
output(0, 113) <= input(17);
output(0, 114) <= input(18);
output(0, 115) <= input(19);
output(0, 116) <= input(20);
output(0, 117) <= input(21);
output(0, 118) <= input(22);
output(0, 119) <= input(23);
output(0, 120) <= input(24);
output(0, 121) <= input(25);
output(0, 122) <= input(26);
output(0, 123) <= input(27);
output(0, 124) <= input(28);
output(0, 125) <= input(29);
output(0, 126) <= input(30);
output(0, 127) <= input(31);
output(0, 128) <= input(32);
output(0, 129) <= input(0);
output(0, 130) <= input(1);
output(0, 131) <= input(2);
output(0, 132) <= input(3);
output(0, 133) <= input(4);
output(0, 134) <= input(5);
output(0, 135) <= input(6);
output(0, 136) <= input(7);
output(0, 137) <= input(8);
output(0, 138) <= input(9);
output(0, 139) <= input(10);
output(0, 140) <= input(11);
output(0, 141) <= input(12);
output(0, 142) <= input(13);
output(0, 143) <= input(14);
output(0, 144) <= input(32);
output(0, 145) <= input(0);
output(0, 146) <= input(1);
output(0, 147) <= input(2);
output(0, 148) <= input(3);
output(0, 149) <= input(4);
output(0, 150) <= input(5);
output(0, 151) <= input(6);
output(0, 152) <= input(7);
output(0, 153) <= input(8);
output(0, 154) <= input(9);
output(0, 155) <= input(10);
output(0, 156) <= input(11);
output(0, 157) <= input(12);
output(0, 158) <= input(13);
output(0, 159) <= input(14);
output(0, 160) <= input(32);
output(0, 161) <= input(0);
output(0, 162) <= input(1);
output(0, 163) <= input(2);
output(0, 164) <= input(3);
output(0, 165) <= input(4);
output(0, 166) <= input(5);
output(0, 167) <= input(6);
output(0, 168) <= input(7);
output(0, 169) <= input(8);
output(0, 170) <= input(9);
output(0, 171) <= input(10);
output(0, 172) <= input(11);
output(0, 173) <= input(12);
output(0, 174) <= input(13);
output(0, 175) <= input(14);
output(0, 176) <= input(32);
output(0, 177) <= input(0);
output(0, 178) <= input(1);
output(0, 179) <= input(2);
output(0, 180) <= input(3);
output(0, 181) <= input(4);
output(0, 182) <= input(5);
output(0, 183) <= input(6);
output(0, 184) <= input(7);
output(0, 185) <= input(8);
output(0, 186) <= input(9);
output(0, 187) <= input(10);
output(0, 188) <= input(11);
output(0, 189) <= input(12);
output(0, 190) <= input(13);
output(0, 191) <= input(14);
output(0, 192) <= input(33);
output(0, 193) <= input(16);
output(0, 194) <= input(17);
output(0, 195) <= input(18);
output(0, 196) <= input(19);
output(0, 197) <= input(20);
output(0, 198) <= input(21);
output(0, 199) <= input(22);
output(0, 200) <= input(23);
output(0, 201) <= input(24);
output(0, 202) <= input(25);
output(0, 203) <= input(26);
output(0, 204) <= input(27);
output(0, 205) <= input(28);
output(0, 206) <= input(29);
output(0, 207) <= input(30);
output(0, 208) <= input(33);
output(0, 209) <= input(16);
output(0, 210) <= input(17);
output(0, 211) <= input(18);
output(0, 212) <= input(19);
output(0, 213) <= input(20);
output(0, 214) <= input(21);
output(0, 215) <= input(22);
output(0, 216) <= input(23);
output(0, 217) <= input(24);
output(0, 218) <= input(25);
output(0, 219) <= input(26);
output(0, 220) <= input(27);
output(0, 221) <= input(28);
output(0, 222) <= input(29);
output(0, 223) <= input(30);
output(0, 224) <= input(33);
output(0, 225) <= input(16);
output(0, 226) <= input(17);
output(0, 227) <= input(18);
output(0, 228) <= input(19);
output(0, 229) <= input(20);
output(0, 230) <= input(21);
output(0, 231) <= input(22);
output(0, 232) <= input(23);
output(0, 233) <= input(24);
output(0, 234) <= input(25);
output(0, 235) <= input(26);
output(0, 236) <= input(27);
output(0, 237) <= input(28);
output(0, 238) <= input(29);
output(0, 239) <= input(30);
output(0, 240) <= input(33);
output(0, 241) <= input(16);
output(0, 242) <= input(17);
output(0, 243) <= input(18);
output(0, 244) <= input(19);
output(0, 245) <= input(20);
output(0, 246) <= input(21);
output(0, 247) <= input(22);
output(0, 248) <= input(23);
output(0, 249) <= input(24);
output(0, 250) <= input(25);
output(0, 251) <= input(26);
output(0, 252) <= input(27);
output(0, 253) <= input(28);
output(0, 254) <= input(29);
output(0, 255) <= input(30);
output(1, 0) <= input(0);
output(1, 1) <= input(1);
output(1, 2) <= input(2);
output(1, 3) <= input(3);
output(1, 4) <= input(4);
output(1, 5) <= input(5);
output(1, 6) <= input(6);
output(1, 7) <= input(7);
output(1, 8) <= input(8);
output(1, 9) <= input(9);
output(1, 10) <= input(10);
output(1, 11) <= input(11);
output(1, 12) <= input(12);
output(1, 13) <= input(13);
output(1, 14) <= input(14);
output(1, 15) <= input(15);
output(1, 16) <= input(0);
output(1, 17) <= input(1);
output(1, 18) <= input(2);
output(1, 19) <= input(3);
output(1, 20) <= input(4);
output(1, 21) <= input(5);
output(1, 22) <= input(6);
output(1, 23) <= input(7);
output(1, 24) <= input(8);
output(1, 25) <= input(9);
output(1, 26) <= input(10);
output(1, 27) <= input(11);
output(1, 28) <= input(12);
output(1, 29) <= input(13);
output(1, 30) <= input(14);
output(1, 31) <= input(15);
output(1, 32) <= input(16);
output(1, 33) <= input(17);
output(1, 34) <= input(18);
output(1, 35) <= input(19);
output(1, 36) <= input(20);
output(1, 37) <= input(21);
output(1, 38) <= input(22);
output(1, 39) <= input(23);
output(1, 40) <= input(24);
output(1, 41) <= input(25);
output(1, 42) <= input(26);
output(1, 43) <= input(27);
output(1, 44) <= input(28);
output(1, 45) <= input(29);
output(1, 46) <= input(30);
output(1, 47) <= input(31);
output(1, 48) <= input(16);
output(1, 49) <= input(17);
output(1, 50) <= input(18);
output(1, 51) <= input(19);
output(1, 52) <= input(20);
output(1, 53) <= input(21);
output(1, 54) <= input(22);
output(1, 55) <= input(23);
output(1, 56) <= input(24);
output(1, 57) <= input(25);
output(1, 58) <= input(26);
output(1, 59) <= input(27);
output(1, 60) <= input(28);
output(1, 61) <= input(29);
output(1, 62) <= input(30);
output(1, 63) <= input(31);
output(1, 64) <= input(16);
output(1, 65) <= input(17);
output(1, 66) <= input(18);
output(1, 67) <= input(19);
output(1, 68) <= input(20);
output(1, 69) <= input(21);
output(1, 70) <= input(22);
output(1, 71) <= input(23);
output(1, 72) <= input(24);
output(1, 73) <= input(25);
output(1, 74) <= input(26);
output(1, 75) <= input(27);
output(1, 76) <= input(28);
output(1, 77) <= input(29);
output(1, 78) <= input(30);
output(1, 79) <= input(31);
output(1, 80) <= input(32);
output(1, 81) <= input(0);
output(1, 82) <= input(1);
output(1, 83) <= input(2);
output(1, 84) <= input(3);
output(1, 85) <= input(4);
output(1, 86) <= input(5);
output(1, 87) <= input(6);
output(1, 88) <= input(7);
output(1, 89) <= input(8);
output(1, 90) <= input(9);
output(1, 91) <= input(10);
output(1, 92) <= input(11);
output(1, 93) <= input(12);
output(1, 94) <= input(13);
output(1, 95) <= input(14);
output(1, 96) <= input(32);
output(1, 97) <= input(0);
output(1, 98) <= input(1);
output(1, 99) <= input(2);
output(1, 100) <= input(3);
output(1, 101) <= input(4);
output(1, 102) <= input(5);
output(1, 103) <= input(6);
output(1, 104) <= input(7);
output(1, 105) <= input(8);
output(1, 106) <= input(9);
output(1, 107) <= input(10);
output(1, 108) <= input(11);
output(1, 109) <= input(12);
output(1, 110) <= input(13);
output(1, 111) <= input(14);
output(1, 112) <= input(32);
output(1, 113) <= input(0);
output(1, 114) <= input(1);
output(1, 115) <= input(2);
output(1, 116) <= input(3);
output(1, 117) <= input(4);
output(1, 118) <= input(5);
output(1, 119) <= input(6);
output(1, 120) <= input(7);
output(1, 121) <= input(8);
output(1, 122) <= input(9);
output(1, 123) <= input(10);
output(1, 124) <= input(11);
output(1, 125) <= input(12);
output(1, 126) <= input(13);
output(1, 127) <= input(14);
output(1, 128) <= input(33);
output(1, 129) <= input(16);
output(1, 130) <= input(17);
output(1, 131) <= input(18);
output(1, 132) <= input(19);
output(1, 133) <= input(20);
output(1, 134) <= input(21);
output(1, 135) <= input(22);
output(1, 136) <= input(23);
output(1, 137) <= input(24);
output(1, 138) <= input(25);
output(1, 139) <= input(26);
output(1, 140) <= input(27);
output(1, 141) <= input(28);
output(1, 142) <= input(29);
output(1, 143) <= input(30);
output(1, 144) <= input(33);
output(1, 145) <= input(16);
output(1, 146) <= input(17);
output(1, 147) <= input(18);
output(1, 148) <= input(19);
output(1, 149) <= input(20);
output(1, 150) <= input(21);
output(1, 151) <= input(22);
output(1, 152) <= input(23);
output(1, 153) <= input(24);
output(1, 154) <= input(25);
output(1, 155) <= input(26);
output(1, 156) <= input(27);
output(1, 157) <= input(28);
output(1, 158) <= input(29);
output(1, 159) <= input(30);
output(1, 160) <= input(34);
output(1, 161) <= input(32);
output(1, 162) <= input(0);
output(1, 163) <= input(1);
output(1, 164) <= input(2);
output(1, 165) <= input(3);
output(1, 166) <= input(4);
output(1, 167) <= input(5);
output(1, 168) <= input(6);
output(1, 169) <= input(7);
output(1, 170) <= input(8);
output(1, 171) <= input(9);
output(1, 172) <= input(10);
output(1, 173) <= input(11);
output(1, 174) <= input(12);
output(1, 175) <= input(13);
output(1, 176) <= input(34);
output(1, 177) <= input(32);
output(1, 178) <= input(0);
output(1, 179) <= input(1);
output(1, 180) <= input(2);
output(1, 181) <= input(3);
output(1, 182) <= input(4);
output(1, 183) <= input(5);
output(1, 184) <= input(6);
output(1, 185) <= input(7);
output(1, 186) <= input(8);
output(1, 187) <= input(9);
output(1, 188) <= input(10);
output(1, 189) <= input(11);
output(1, 190) <= input(12);
output(1, 191) <= input(13);
output(1, 192) <= input(34);
output(1, 193) <= input(32);
output(1, 194) <= input(0);
output(1, 195) <= input(1);
output(1, 196) <= input(2);
output(1, 197) <= input(3);
output(1, 198) <= input(4);
output(1, 199) <= input(5);
output(1, 200) <= input(6);
output(1, 201) <= input(7);
output(1, 202) <= input(8);
output(1, 203) <= input(9);
output(1, 204) <= input(10);
output(1, 205) <= input(11);
output(1, 206) <= input(12);
output(1, 207) <= input(13);
output(1, 208) <= input(35);
output(1, 209) <= input(33);
output(1, 210) <= input(16);
output(1, 211) <= input(17);
output(1, 212) <= input(18);
output(1, 213) <= input(19);
output(1, 214) <= input(20);
output(1, 215) <= input(21);
output(1, 216) <= input(22);
output(1, 217) <= input(23);
output(1, 218) <= input(24);
output(1, 219) <= input(25);
output(1, 220) <= input(26);
output(1, 221) <= input(27);
output(1, 222) <= input(28);
output(1, 223) <= input(29);
output(1, 224) <= input(35);
output(1, 225) <= input(33);
output(1, 226) <= input(16);
output(1, 227) <= input(17);
output(1, 228) <= input(18);
output(1, 229) <= input(19);
output(1, 230) <= input(20);
output(1, 231) <= input(21);
output(1, 232) <= input(22);
output(1, 233) <= input(23);
output(1, 234) <= input(24);
output(1, 235) <= input(25);
output(1, 236) <= input(26);
output(1, 237) <= input(27);
output(1, 238) <= input(28);
output(1, 239) <= input(29);
output(1, 240) <= input(35);
output(1, 241) <= input(33);
output(1, 242) <= input(16);
output(1, 243) <= input(17);
output(1, 244) <= input(18);
output(1, 245) <= input(19);
output(1, 246) <= input(20);
output(1, 247) <= input(21);
output(1, 248) <= input(22);
output(1, 249) <= input(23);
output(1, 250) <= input(24);
output(1, 251) <= input(25);
output(1, 252) <= input(26);
output(1, 253) <= input(27);
output(1, 254) <= input(28);
output(1, 255) <= input(29);
output(2, 0) <= input(0);
output(2, 1) <= input(1);
output(2, 2) <= input(2);
output(2, 3) <= input(3);
output(2, 4) <= input(4);
output(2, 5) <= input(5);
output(2, 6) <= input(6);
output(2, 7) <= input(7);
output(2, 8) <= input(8);
output(2, 9) <= input(9);
output(2, 10) <= input(10);
output(2, 11) <= input(11);
output(2, 12) <= input(12);
output(2, 13) <= input(13);
output(2, 14) <= input(14);
output(2, 15) <= input(15);
output(2, 16) <= input(0);
output(2, 17) <= input(1);
output(2, 18) <= input(2);
output(2, 19) <= input(3);
output(2, 20) <= input(4);
output(2, 21) <= input(5);
output(2, 22) <= input(6);
output(2, 23) <= input(7);
output(2, 24) <= input(8);
output(2, 25) <= input(9);
output(2, 26) <= input(10);
output(2, 27) <= input(11);
output(2, 28) <= input(12);
output(2, 29) <= input(13);
output(2, 30) <= input(14);
output(2, 31) <= input(15);
output(2, 32) <= input(16);
output(2, 33) <= input(17);
output(2, 34) <= input(18);
output(2, 35) <= input(19);
output(2, 36) <= input(20);
output(2, 37) <= input(21);
output(2, 38) <= input(22);
output(2, 39) <= input(23);
output(2, 40) <= input(24);
output(2, 41) <= input(25);
output(2, 42) <= input(26);
output(2, 43) <= input(27);
output(2, 44) <= input(28);
output(2, 45) <= input(29);
output(2, 46) <= input(30);
output(2, 47) <= input(31);
output(2, 48) <= input(16);
output(2, 49) <= input(17);
output(2, 50) <= input(18);
output(2, 51) <= input(19);
output(2, 52) <= input(20);
output(2, 53) <= input(21);
output(2, 54) <= input(22);
output(2, 55) <= input(23);
output(2, 56) <= input(24);
output(2, 57) <= input(25);
output(2, 58) <= input(26);
output(2, 59) <= input(27);
output(2, 60) <= input(28);
output(2, 61) <= input(29);
output(2, 62) <= input(30);
output(2, 63) <= input(31);
output(2, 64) <= input(32);
output(2, 65) <= input(0);
output(2, 66) <= input(1);
output(2, 67) <= input(2);
output(2, 68) <= input(3);
output(2, 69) <= input(4);
output(2, 70) <= input(5);
output(2, 71) <= input(6);
output(2, 72) <= input(7);
output(2, 73) <= input(8);
output(2, 74) <= input(9);
output(2, 75) <= input(10);
output(2, 76) <= input(11);
output(2, 77) <= input(12);
output(2, 78) <= input(13);
output(2, 79) <= input(14);
output(2, 80) <= input(32);
output(2, 81) <= input(0);
output(2, 82) <= input(1);
output(2, 83) <= input(2);
output(2, 84) <= input(3);
output(2, 85) <= input(4);
output(2, 86) <= input(5);
output(2, 87) <= input(6);
output(2, 88) <= input(7);
output(2, 89) <= input(8);
output(2, 90) <= input(9);
output(2, 91) <= input(10);
output(2, 92) <= input(11);
output(2, 93) <= input(12);
output(2, 94) <= input(13);
output(2, 95) <= input(14);
output(2, 96) <= input(33);
output(2, 97) <= input(16);
output(2, 98) <= input(17);
output(2, 99) <= input(18);
output(2, 100) <= input(19);
output(2, 101) <= input(20);
output(2, 102) <= input(21);
output(2, 103) <= input(22);
output(2, 104) <= input(23);
output(2, 105) <= input(24);
output(2, 106) <= input(25);
output(2, 107) <= input(26);
output(2, 108) <= input(27);
output(2, 109) <= input(28);
output(2, 110) <= input(29);
output(2, 111) <= input(30);
output(2, 112) <= input(33);
output(2, 113) <= input(16);
output(2, 114) <= input(17);
output(2, 115) <= input(18);
output(2, 116) <= input(19);
output(2, 117) <= input(20);
output(2, 118) <= input(21);
output(2, 119) <= input(22);
output(2, 120) <= input(23);
output(2, 121) <= input(24);
output(2, 122) <= input(25);
output(2, 123) <= input(26);
output(2, 124) <= input(27);
output(2, 125) <= input(28);
output(2, 126) <= input(29);
output(2, 127) <= input(30);
output(2, 128) <= input(34);
output(2, 129) <= input(32);
output(2, 130) <= input(0);
output(2, 131) <= input(1);
output(2, 132) <= input(2);
output(2, 133) <= input(3);
output(2, 134) <= input(4);
output(2, 135) <= input(5);
output(2, 136) <= input(6);
output(2, 137) <= input(7);
output(2, 138) <= input(8);
output(2, 139) <= input(9);
output(2, 140) <= input(10);
output(2, 141) <= input(11);
output(2, 142) <= input(12);
output(2, 143) <= input(13);
output(2, 144) <= input(34);
output(2, 145) <= input(32);
output(2, 146) <= input(0);
output(2, 147) <= input(1);
output(2, 148) <= input(2);
output(2, 149) <= input(3);
output(2, 150) <= input(4);
output(2, 151) <= input(5);
output(2, 152) <= input(6);
output(2, 153) <= input(7);
output(2, 154) <= input(8);
output(2, 155) <= input(9);
output(2, 156) <= input(10);
output(2, 157) <= input(11);
output(2, 158) <= input(12);
output(2, 159) <= input(13);
output(2, 160) <= input(35);
output(2, 161) <= input(33);
output(2, 162) <= input(16);
output(2, 163) <= input(17);
output(2, 164) <= input(18);
output(2, 165) <= input(19);
output(2, 166) <= input(20);
output(2, 167) <= input(21);
output(2, 168) <= input(22);
output(2, 169) <= input(23);
output(2, 170) <= input(24);
output(2, 171) <= input(25);
output(2, 172) <= input(26);
output(2, 173) <= input(27);
output(2, 174) <= input(28);
output(2, 175) <= input(29);
output(2, 176) <= input(35);
output(2, 177) <= input(33);
output(2, 178) <= input(16);
output(2, 179) <= input(17);
output(2, 180) <= input(18);
output(2, 181) <= input(19);
output(2, 182) <= input(20);
output(2, 183) <= input(21);
output(2, 184) <= input(22);
output(2, 185) <= input(23);
output(2, 186) <= input(24);
output(2, 187) <= input(25);
output(2, 188) <= input(26);
output(2, 189) <= input(27);
output(2, 190) <= input(28);
output(2, 191) <= input(29);
output(2, 192) <= input(36);
output(2, 193) <= input(34);
output(2, 194) <= input(32);
output(2, 195) <= input(0);
output(2, 196) <= input(1);
output(2, 197) <= input(2);
output(2, 198) <= input(3);
output(2, 199) <= input(4);
output(2, 200) <= input(5);
output(2, 201) <= input(6);
output(2, 202) <= input(7);
output(2, 203) <= input(8);
output(2, 204) <= input(9);
output(2, 205) <= input(10);
output(2, 206) <= input(11);
output(2, 207) <= input(12);
output(2, 208) <= input(36);
output(2, 209) <= input(34);
output(2, 210) <= input(32);
output(2, 211) <= input(0);
output(2, 212) <= input(1);
output(2, 213) <= input(2);
output(2, 214) <= input(3);
output(2, 215) <= input(4);
output(2, 216) <= input(5);
output(2, 217) <= input(6);
output(2, 218) <= input(7);
output(2, 219) <= input(8);
output(2, 220) <= input(9);
output(2, 221) <= input(10);
output(2, 222) <= input(11);
output(2, 223) <= input(12);
output(2, 224) <= input(37);
output(2, 225) <= input(35);
output(2, 226) <= input(33);
output(2, 227) <= input(16);
output(2, 228) <= input(17);
output(2, 229) <= input(18);
output(2, 230) <= input(19);
output(2, 231) <= input(20);
output(2, 232) <= input(21);
output(2, 233) <= input(22);
output(2, 234) <= input(23);
output(2, 235) <= input(24);
output(2, 236) <= input(25);
output(2, 237) <= input(26);
output(2, 238) <= input(27);
output(2, 239) <= input(28);
output(2, 240) <= input(37);
output(2, 241) <= input(35);
output(2, 242) <= input(33);
output(2, 243) <= input(16);
output(2, 244) <= input(17);
output(2, 245) <= input(18);
output(2, 246) <= input(19);
output(2, 247) <= input(20);
output(2, 248) <= input(21);
output(2, 249) <= input(22);
output(2, 250) <= input(23);
output(2, 251) <= input(24);
output(2, 252) <= input(25);
output(2, 253) <= input(26);
output(2, 254) <= input(27);
output(2, 255) <= input(28);
when "0100" =>
output(0, 0) <= input(0);
output(0, 1) <= input(1);
output(0, 2) <= input(2);
output(0, 3) <= input(3);
output(0, 4) <= input(4);
output(0, 5) <= input(5);
output(0, 6) <= input(6);
output(0, 7) <= input(7);
output(0, 8) <= input(8);
output(0, 9) <= input(9);
output(0, 10) <= input(10);
output(0, 11) <= input(11);
output(0, 12) <= input(12);
output(0, 13) <= input(13);
output(0, 14) <= input(14);
output(0, 15) <= input(15);
output(0, 16) <= input(16);
output(0, 17) <= input(17);
output(0, 18) <= input(18);
output(0, 19) <= input(19);
output(0, 20) <= input(20);
output(0, 21) <= input(21);
output(0, 22) <= input(22);
output(0, 23) <= input(23);
output(0, 24) <= input(24);
output(0, 25) <= input(25);
output(0, 26) <= input(26);
output(0, 27) <= input(27);
output(0, 28) <= input(28);
output(0, 29) <= input(29);
output(0, 30) <= input(30);
output(0, 31) <= input(31);
output(0, 32) <= input(16);
output(0, 33) <= input(17);
output(0, 34) <= input(18);
output(0, 35) <= input(19);
output(0, 36) <= input(20);
output(0, 37) <= input(21);
output(0, 38) <= input(22);
output(0, 39) <= input(23);
output(0, 40) <= input(24);
output(0, 41) <= input(25);
output(0, 42) <= input(26);
output(0, 43) <= input(27);
output(0, 44) <= input(28);
output(0, 45) <= input(29);
output(0, 46) <= input(30);
output(0, 47) <= input(31);
output(0, 48) <= input(32);
output(0, 49) <= input(0);
output(0, 50) <= input(1);
output(0, 51) <= input(2);
output(0, 52) <= input(3);
output(0, 53) <= input(4);
output(0, 54) <= input(5);
output(0, 55) <= input(6);
output(0, 56) <= input(7);
output(0, 57) <= input(8);
output(0, 58) <= input(9);
output(0, 59) <= input(10);
output(0, 60) <= input(11);
output(0, 61) <= input(12);
output(0, 62) <= input(13);
output(0, 63) <= input(14);
output(0, 64) <= input(33);
output(0, 65) <= input(16);
output(0, 66) <= input(17);
output(0, 67) <= input(18);
output(0, 68) <= input(19);
output(0, 69) <= input(20);
output(0, 70) <= input(21);
output(0, 71) <= input(22);
output(0, 72) <= input(23);
output(0, 73) <= input(24);
output(0, 74) <= input(25);
output(0, 75) <= input(26);
output(0, 76) <= input(27);
output(0, 77) <= input(28);
output(0, 78) <= input(29);
output(0, 79) <= input(30);
output(0, 80) <= input(33);
output(0, 81) <= input(16);
output(0, 82) <= input(17);
output(0, 83) <= input(18);
output(0, 84) <= input(19);
output(0, 85) <= input(20);
output(0, 86) <= input(21);
output(0, 87) <= input(22);
output(0, 88) <= input(23);
output(0, 89) <= input(24);
output(0, 90) <= input(25);
output(0, 91) <= input(26);
output(0, 92) <= input(27);
output(0, 93) <= input(28);
output(0, 94) <= input(29);
output(0, 95) <= input(30);
output(0, 96) <= input(34);
output(0, 97) <= input(32);
output(0, 98) <= input(0);
output(0, 99) <= input(1);
output(0, 100) <= input(2);
output(0, 101) <= input(3);
output(0, 102) <= input(4);
output(0, 103) <= input(5);
output(0, 104) <= input(6);
output(0, 105) <= input(7);
output(0, 106) <= input(8);
output(0, 107) <= input(9);
output(0, 108) <= input(10);
output(0, 109) <= input(11);
output(0, 110) <= input(12);
output(0, 111) <= input(13);
output(0, 112) <= input(34);
output(0, 113) <= input(32);
output(0, 114) <= input(0);
output(0, 115) <= input(1);
output(0, 116) <= input(2);
output(0, 117) <= input(3);
output(0, 118) <= input(4);
output(0, 119) <= input(5);
output(0, 120) <= input(6);
output(0, 121) <= input(7);
output(0, 122) <= input(8);
output(0, 123) <= input(9);
output(0, 124) <= input(10);
output(0, 125) <= input(11);
output(0, 126) <= input(12);
output(0, 127) <= input(13);
output(0, 128) <= input(35);
output(0, 129) <= input(33);
output(0, 130) <= input(16);
output(0, 131) <= input(17);
output(0, 132) <= input(18);
output(0, 133) <= input(19);
output(0, 134) <= input(20);
output(0, 135) <= input(21);
output(0, 136) <= input(22);
output(0, 137) <= input(23);
output(0, 138) <= input(24);
output(0, 139) <= input(25);
output(0, 140) <= input(26);
output(0, 141) <= input(27);
output(0, 142) <= input(28);
output(0, 143) <= input(29);
output(0, 144) <= input(36);
output(0, 145) <= input(34);
output(0, 146) <= input(32);
output(0, 147) <= input(0);
output(0, 148) <= input(1);
output(0, 149) <= input(2);
output(0, 150) <= input(3);
output(0, 151) <= input(4);
output(0, 152) <= input(5);
output(0, 153) <= input(6);
output(0, 154) <= input(7);
output(0, 155) <= input(8);
output(0, 156) <= input(9);
output(0, 157) <= input(10);
output(0, 158) <= input(11);
output(0, 159) <= input(12);
output(0, 160) <= input(36);
output(0, 161) <= input(34);
output(0, 162) <= input(32);
output(0, 163) <= input(0);
output(0, 164) <= input(1);
output(0, 165) <= input(2);
output(0, 166) <= input(3);
output(0, 167) <= input(4);
output(0, 168) <= input(5);
output(0, 169) <= input(6);
output(0, 170) <= input(7);
output(0, 171) <= input(8);
output(0, 172) <= input(9);
output(0, 173) <= input(10);
output(0, 174) <= input(11);
output(0, 175) <= input(12);
output(0, 176) <= input(37);
output(0, 177) <= input(35);
output(0, 178) <= input(33);
output(0, 179) <= input(16);
output(0, 180) <= input(17);
output(0, 181) <= input(18);
output(0, 182) <= input(19);
output(0, 183) <= input(20);
output(0, 184) <= input(21);
output(0, 185) <= input(22);
output(0, 186) <= input(23);
output(0, 187) <= input(24);
output(0, 188) <= input(25);
output(0, 189) <= input(26);
output(0, 190) <= input(27);
output(0, 191) <= input(28);
output(0, 192) <= input(38);
output(0, 193) <= input(36);
output(0, 194) <= input(34);
output(0, 195) <= input(32);
output(0, 196) <= input(0);
output(0, 197) <= input(1);
output(0, 198) <= input(2);
output(0, 199) <= input(3);
output(0, 200) <= input(4);
output(0, 201) <= input(5);
output(0, 202) <= input(6);
output(0, 203) <= input(7);
output(0, 204) <= input(8);
output(0, 205) <= input(9);
output(0, 206) <= input(10);
output(0, 207) <= input(11);
output(0, 208) <= input(38);
output(0, 209) <= input(36);
output(0, 210) <= input(34);
output(0, 211) <= input(32);
output(0, 212) <= input(0);
output(0, 213) <= input(1);
output(0, 214) <= input(2);
output(0, 215) <= input(3);
output(0, 216) <= input(4);
output(0, 217) <= input(5);
output(0, 218) <= input(6);
output(0, 219) <= input(7);
output(0, 220) <= input(8);
output(0, 221) <= input(9);
output(0, 222) <= input(10);
output(0, 223) <= input(11);
output(0, 224) <= input(39);
output(0, 225) <= input(37);
output(0, 226) <= input(35);
output(0, 227) <= input(33);
output(0, 228) <= input(16);
output(0, 229) <= input(17);
output(0, 230) <= input(18);
output(0, 231) <= input(19);
output(0, 232) <= input(20);
output(0, 233) <= input(21);
output(0, 234) <= input(22);
output(0, 235) <= input(23);
output(0, 236) <= input(24);
output(0, 237) <= input(25);
output(0, 238) <= input(26);
output(0, 239) <= input(27);
output(0, 240) <= input(39);
output(0, 241) <= input(37);
output(0, 242) <= input(35);
output(0, 243) <= input(33);
output(0, 244) <= input(16);
output(0, 245) <= input(17);
output(0, 246) <= input(18);
output(0, 247) <= input(19);
output(0, 248) <= input(20);
output(0, 249) <= input(21);
output(0, 250) <= input(22);
output(0, 251) <= input(23);
output(0, 252) <= input(24);
output(0, 253) <= input(25);
output(0, 254) <= input(26);
output(0, 255) <= input(27);
output(1, 0) <= input(0);
output(1, 1) <= input(1);
output(1, 2) <= input(2);
output(1, 3) <= input(3);
output(1, 4) <= input(4);
output(1, 5) <= input(5);
output(1, 6) <= input(6);
output(1, 7) <= input(7);
output(1, 8) <= input(8);
output(1, 9) <= input(9);
output(1, 10) <= input(10);
output(1, 11) <= input(11);
output(1, 12) <= input(12);
output(1, 13) <= input(13);
output(1, 14) <= input(14);
output(1, 15) <= input(15);
output(1, 16) <= input(16);
output(1, 17) <= input(17);
output(1, 18) <= input(18);
output(1, 19) <= input(19);
output(1, 20) <= input(20);
output(1, 21) <= input(21);
output(1, 22) <= input(22);
output(1, 23) <= input(23);
output(1, 24) <= input(24);
output(1, 25) <= input(25);
output(1, 26) <= input(26);
output(1, 27) <= input(27);
output(1, 28) <= input(28);
output(1, 29) <= input(29);
output(1, 30) <= input(30);
output(1, 31) <= input(31);
output(1, 32) <= input(32);
output(1, 33) <= input(0);
output(1, 34) <= input(1);
output(1, 35) <= input(2);
output(1, 36) <= input(3);
output(1, 37) <= input(4);
output(1, 38) <= input(5);
output(1, 39) <= input(6);
output(1, 40) <= input(7);
output(1, 41) <= input(8);
output(1, 42) <= input(9);
output(1, 43) <= input(10);
output(1, 44) <= input(11);
output(1, 45) <= input(12);
output(1, 46) <= input(13);
output(1, 47) <= input(14);
output(1, 48) <= input(32);
output(1, 49) <= input(0);
output(1, 50) <= input(1);
output(1, 51) <= input(2);
output(1, 52) <= input(3);
output(1, 53) <= input(4);
output(1, 54) <= input(5);
output(1, 55) <= input(6);
output(1, 56) <= input(7);
output(1, 57) <= input(8);
output(1, 58) <= input(9);
output(1, 59) <= input(10);
output(1, 60) <= input(11);
output(1, 61) <= input(12);
output(1, 62) <= input(13);
output(1, 63) <= input(14);
output(1, 64) <= input(33);
output(1, 65) <= input(16);
output(1, 66) <= input(17);
output(1, 67) <= input(18);
output(1, 68) <= input(19);
output(1, 69) <= input(20);
output(1, 70) <= input(21);
output(1, 71) <= input(22);
output(1, 72) <= input(23);
output(1, 73) <= input(24);
output(1, 74) <= input(25);
output(1, 75) <= input(26);
output(1, 76) <= input(27);
output(1, 77) <= input(28);
output(1, 78) <= input(29);
output(1, 79) <= input(30);
output(1, 80) <= input(34);
output(1, 81) <= input(32);
output(1, 82) <= input(0);
output(1, 83) <= input(1);
output(1, 84) <= input(2);
output(1, 85) <= input(3);
output(1, 86) <= input(4);
output(1, 87) <= input(5);
output(1, 88) <= input(6);
output(1, 89) <= input(7);
output(1, 90) <= input(8);
output(1, 91) <= input(9);
output(1, 92) <= input(10);
output(1, 93) <= input(11);
output(1, 94) <= input(12);
output(1, 95) <= input(13);
output(1, 96) <= input(35);
output(1, 97) <= input(33);
output(1, 98) <= input(16);
output(1, 99) <= input(17);
output(1, 100) <= input(18);
output(1, 101) <= input(19);
output(1, 102) <= input(20);
output(1, 103) <= input(21);
output(1, 104) <= input(22);
output(1, 105) <= input(23);
output(1, 106) <= input(24);
output(1, 107) <= input(25);
output(1, 108) <= input(26);
output(1, 109) <= input(27);
output(1, 110) <= input(28);
output(1, 111) <= input(29);
output(1, 112) <= input(35);
output(1, 113) <= input(33);
output(1, 114) <= input(16);
output(1, 115) <= input(17);
output(1, 116) <= input(18);
output(1, 117) <= input(19);
output(1, 118) <= input(20);
output(1, 119) <= input(21);
output(1, 120) <= input(22);
output(1, 121) <= input(23);
output(1, 122) <= input(24);
output(1, 123) <= input(25);
output(1, 124) <= input(26);
output(1, 125) <= input(27);
output(1, 126) <= input(28);
output(1, 127) <= input(29);
output(1, 128) <= input(36);
output(1, 129) <= input(34);
output(1, 130) <= input(32);
output(1, 131) <= input(0);
output(1, 132) <= input(1);
output(1, 133) <= input(2);
output(1, 134) <= input(3);
output(1, 135) <= input(4);
output(1, 136) <= input(5);
output(1, 137) <= input(6);
output(1, 138) <= input(7);
output(1, 139) <= input(8);
output(1, 140) <= input(9);
output(1, 141) <= input(10);
output(1, 142) <= input(11);
output(1, 143) <= input(12);
output(1, 144) <= input(37);
output(1, 145) <= input(35);
output(1, 146) <= input(33);
output(1, 147) <= input(16);
output(1, 148) <= input(17);
output(1, 149) <= input(18);
output(1, 150) <= input(19);
output(1, 151) <= input(20);
output(1, 152) <= input(21);
output(1, 153) <= input(22);
output(1, 154) <= input(23);
output(1, 155) <= input(24);
output(1, 156) <= input(25);
output(1, 157) <= input(26);
output(1, 158) <= input(27);
output(1, 159) <= input(28);
output(1, 160) <= input(38);
output(1, 161) <= input(36);
output(1, 162) <= input(34);
output(1, 163) <= input(32);
output(1, 164) <= input(0);
output(1, 165) <= input(1);
output(1, 166) <= input(2);
output(1, 167) <= input(3);
output(1, 168) <= input(4);
output(1, 169) <= input(5);
output(1, 170) <= input(6);
output(1, 171) <= input(7);
output(1, 172) <= input(8);
output(1, 173) <= input(9);
output(1, 174) <= input(10);
output(1, 175) <= input(11);
output(1, 176) <= input(38);
output(1, 177) <= input(36);
output(1, 178) <= input(34);
output(1, 179) <= input(32);
output(1, 180) <= input(0);
output(1, 181) <= input(1);
output(1, 182) <= input(2);
output(1, 183) <= input(3);
output(1, 184) <= input(4);
output(1, 185) <= input(5);
output(1, 186) <= input(6);
output(1, 187) <= input(7);
output(1, 188) <= input(8);
output(1, 189) <= input(9);
output(1, 190) <= input(10);
output(1, 191) <= input(11);
output(1, 192) <= input(39);
output(1, 193) <= input(37);
output(1, 194) <= input(35);
output(1, 195) <= input(33);
output(1, 196) <= input(16);
output(1, 197) <= input(17);
output(1, 198) <= input(18);
output(1, 199) <= input(19);
output(1, 200) <= input(20);
output(1, 201) <= input(21);
output(1, 202) <= input(22);
output(1, 203) <= input(23);
output(1, 204) <= input(24);
output(1, 205) <= input(25);
output(1, 206) <= input(26);
output(1, 207) <= input(27);
output(1, 208) <= input(40);
output(1, 209) <= input(38);
output(1, 210) <= input(36);
output(1, 211) <= input(34);
output(1, 212) <= input(32);
output(1, 213) <= input(0);
output(1, 214) <= input(1);
output(1, 215) <= input(2);
output(1, 216) <= input(3);
output(1, 217) <= input(4);
output(1, 218) <= input(5);
output(1, 219) <= input(6);
output(1, 220) <= input(7);
output(1, 221) <= input(8);
output(1, 222) <= input(9);
output(1, 223) <= input(10);
output(1, 224) <= input(41);
output(1, 225) <= input(39);
output(1, 226) <= input(37);
output(1, 227) <= input(35);
output(1, 228) <= input(33);
output(1, 229) <= input(16);
output(1, 230) <= input(17);
output(1, 231) <= input(18);
output(1, 232) <= input(19);
output(1, 233) <= input(20);
output(1, 234) <= input(21);
output(1, 235) <= input(22);
output(1, 236) <= input(23);
output(1, 237) <= input(24);
output(1, 238) <= input(25);
output(1, 239) <= input(26);
output(1, 240) <= input(41);
output(1, 241) <= input(39);
output(1, 242) <= input(37);
output(1, 243) <= input(35);
output(1, 244) <= input(33);
output(1, 245) <= input(16);
output(1, 246) <= input(17);
output(1, 247) <= input(18);
output(1, 248) <= input(19);
output(1, 249) <= input(20);
output(1, 250) <= input(21);
output(1, 251) <= input(22);
output(1, 252) <= input(23);
output(1, 253) <= input(24);
output(1, 254) <= input(25);
output(1, 255) <= input(26);
output(2, 0) <= input(0);
output(2, 1) <= input(1);
output(2, 2) <= input(2);
output(2, 3) <= input(3);
output(2, 4) <= input(4);
output(2, 5) <= input(5);
output(2, 6) <= input(6);
output(2, 7) <= input(7);
output(2, 8) <= input(8);
output(2, 9) <= input(9);
output(2, 10) <= input(10);
output(2, 11) <= input(11);
output(2, 12) <= input(12);
output(2, 13) <= input(13);
output(2, 14) <= input(14);
output(2, 15) <= input(15);
output(2, 16) <= input(16);
output(2, 17) <= input(17);
output(2, 18) <= input(18);
output(2, 19) <= input(19);
output(2, 20) <= input(20);
output(2, 21) <= input(21);
output(2, 22) <= input(22);
output(2, 23) <= input(23);
output(2, 24) <= input(24);
output(2, 25) <= input(25);
output(2, 26) <= input(26);
output(2, 27) <= input(27);
output(2, 28) <= input(28);
output(2, 29) <= input(29);
output(2, 30) <= input(30);
output(2, 31) <= input(31);
output(2, 32) <= input(32);
output(2, 33) <= input(0);
output(2, 34) <= input(1);
output(2, 35) <= input(2);
output(2, 36) <= input(3);
output(2, 37) <= input(4);
output(2, 38) <= input(5);
output(2, 39) <= input(6);
output(2, 40) <= input(7);
output(2, 41) <= input(8);
output(2, 42) <= input(9);
output(2, 43) <= input(10);
output(2, 44) <= input(11);
output(2, 45) <= input(12);
output(2, 46) <= input(13);
output(2, 47) <= input(14);
output(2, 48) <= input(33);
output(2, 49) <= input(16);
output(2, 50) <= input(17);
output(2, 51) <= input(18);
output(2, 52) <= input(19);
output(2, 53) <= input(20);
output(2, 54) <= input(21);
output(2, 55) <= input(22);
output(2, 56) <= input(23);
output(2, 57) <= input(24);
output(2, 58) <= input(25);
output(2, 59) <= input(26);
output(2, 60) <= input(27);
output(2, 61) <= input(28);
output(2, 62) <= input(29);
output(2, 63) <= input(30);
output(2, 64) <= input(34);
output(2, 65) <= input(32);
output(2, 66) <= input(0);
output(2, 67) <= input(1);
output(2, 68) <= input(2);
output(2, 69) <= input(3);
output(2, 70) <= input(4);
output(2, 71) <= input(5);
output(2, 72) <= input(6);
output(2, 73) <= input(7);
output(2, 74) <= input(8);
output(2, 75) <= input(9);
output(2, 76) <= input(10);
output(2, 77) <= input(11);
output(2, 78) <= input(12);
output(2, 79) <= input(13);
output(2, 80) <= input(35);
output(2, 81) <= input(33);
output(2, 82) <= input(16);
output(2, 83) <= input(17);
output(2, 84) <= input(18);
output(2, 85) <= input(19);
output(2, 86) <= input(20);
output(2, 87) <= input(21);
output(2, 88) <= input(22);
output(2, 89) <= input(23);
output(2, 90) <= input(24);
output(2, 91) <= input(25);
output(2, 92) <= input(26);
output(2, 93) <= input(27);
output(2, 94) <= input(28);
output(2, 95) <= input(29);
output(2, 96) <= input(36);
output(2, 97) <= input(34);
output(2, 98) <= input(32);
output(2, 99) <= input(0);
output(2, 100) <= input(1);
output(2, 101) <= input(2);
output(2, 102) <= input(3);
output(2, 103) <= input(4);
output(2, 104) <= input(5);
output(2, 105) <= input(6);
output(2, 106) <= input(7);
output(2, 107) <= input(8);
output(2, 108) <= input(9);
output(2, 109) <= input(10);
output(2, 110) <= input(11);
output(2, 111) <= input(12);
output(2, 112) <= input(36);
output(2, 113) <= input(34);
output(2, 114) <= input(32);
output(2, 115) <= input(0);
output(2, 116) <= input(1);
output(2, 117) <= input(2);
output(2, 118) <= input(3);
output(2, 119) <= input(4);
output(2, 120) <= input(5);
output(2, 121) <= input(6);
output(2, 122) <= input(7);
output(2, 123) <= input(8);
output(2, 124) <= input(9);
output(2, 125) <= input(10);
output(2, 126) <= input(11);
output(2, 127) <= input(12);
output(2, 128) <= input(37);
output(2, 129) <= input(35);
output(2, 130) <= input(33);
output(2, 131) <= input(16);
output(2, 132) <= input(17);
output(2, 133) <= input(18);
output(2, 134) <= input(19);
output(2, 135) <= input(20);
output(2, 136) <= input(21);
output(2, 137) <= input(22);
output(2, 138) <= input(23);
output(2, 139) <= input(24);
output(2, 140) <= input(25);
output(2, 141) <= input(26);
output(2, 142) <= input(27);
output(2, 143) <= input(28);
output(2, 144) <= input(38);
output(2, 145) <= input(36);
output(2, 146) <= input(34);
output(2, 147) <= input(32);
output(2, 148) <= input(0);
output(2, 149) <= input(1);
output(2, 150) <= input(2);
output(2, 151) <= input(3);
output(2, 152) <= input(4);
output(2, 153) <= input(5);
output(2, 154) <= input(6);
output(2, 155) <= input(7);
output(2, 156) <= input(8);
output(2, 157) <= input(9);
output(2, 158) <= input(10);
output(2, 159) <= input(11);
output(2, 160) <= input(39);
output(2, 161) <= input(37);
output(2, 162) <= input(35);
output(2, 163) <= input(33);
output(2, 164) <= input(16);
output(2, 165) <= input(17);
output(2, 166) <= input(18);
output(2, 167) <= input(19);
output(2, 168) <= input(20);
output(2, 169) <= input(21);
output(2, 170) <= input(22);
output(2, 171) <= input(23);
output(2, 172) <= input(24);
output(2, 173) <= input(25);
output(2, 174) <= input(26);
output(2, 175) <= input(27);
output(2, 176) <= input(40);
output(2, 177) <= input(38);
output(2, 178) <= input(36);
output(2, 179) <= input(34);
output(2, 180) <= input(32);
output(2, 181) <= input(0);
output(2, 182) <= input(1);
output(2, 183) <= input(2);
output(2, 184) <= input(3);
output(2, 185) <= input(4);
output(2, 186) <= input(5);
output(2, 187) <= input(6);
output(2, 188) <= input(7);
output(2, 189) <= input(8);
output(2, 190) <= input(9);
output(2, 191) <= input(10);
output(2, 192) <= input(41);
output(2, 193) <= input(39);
output(2, 194) <= input(37);
output(2, 195) <= input(35);
output(2, 196) <= input(33);
output(2, 197) <= input(16);
output(2, 198) <= input(17);
output(2, 199) <= input(18);
output(2, 200) <= input(19);
output(2, 201) <= input(20);
output(2, 202) <= input(21);
output(2, 203) <= input(22);
output(2, 204) <= input(23);
output(2, 205) <= input(24);
output(2, 206) <= input(25);
output(2, 207) <= input(26);
output(2, 208) <= input(42);
output(2, 209) <= input(40);
output(2, 210) <= input(38);
output(2, 211) <= input(36);
output(2, 212) <= input(34);
output(2, 213) <= input(32);
output(2, 214) <= input(0);
output(2, 215) <= input(1);
output(2, 216) <= input(2);
output(2, 217) <= input(3);
output(2, 218) <= input(4);
output(2, 219) <= input(5);
output(2, 220) <= input(6);
output(2, 221) <= input(7);
output(2, 222) <= input(8);
output(2, 223) <= input(9);
output(2, 224) <= input(43);
output(2, 225) <= input(41);
output(2, 226) <= input(39);
output(2, 227) <= input(37);
output(2, 228) <= input(35);
output(2, 229) <= input(33);
output(2, 230) <= input(16);
output(2, 231) <= input(17);
output(2, 232) <= input(18);
output(2, 233) <= input(19);
output(2, 234) <= input(20);
output(2, 235) <= input(21);
output(2, 236) <= input(22);
output(2, 237) <= input(23);
output(2, 238) <= input(24);
output(2, 239) <= input(25);
output(2, 240) <= input(43);
output(2, 241) <= input(41);
output(2, 242) <= input(39);
output(2, 243) <= input(37);
output(2, 244) <= input(35);
output(2, 245) <= input(33);
output(2, 246) <= input(16);
output(2, 247) <= input(17);
output(2, 248) <= input(18);
output(2, 249) <= input(19);
output(2, 250) <= input(20);
output(2, 251) <= input(21);
output(2, 252) <= input(22);
output(2, 253) <= input(23);
output(2, 254) <= input(24);
output(2, 255) <= input(25);
when "0101" =>
output(0, 0) <= input(0);
output(0, 1) <= input(1);
output(0, 2) <= input(2);
output(0, 3) <= input(3);
output(0, 4) <= input(4);
output(0, 5) <= input(5);
output(0, 6) <= input(6);
output(0, 7) <= input(7);
output(0, 8) <= input(8);
output(0, 9) <= input(9);
output(0, 10) <= input(10);
output(0, 11) <= input(11);
output(0, 12) <= input(12);
output(0, 13) <= input(13);
output(0, 14) <= input(14);
output(0, 15) <= input(15);
output(0, 16) <= input(16);
output(0, 17) <= input(17);
output(0, 18) <= input(18);
output(0, 19) <= input(19);
output(0, 20) <= input(20);
output(0, 21) <= input(21);
output(0, 22) <= input(22);
output(0, 23) <= input(23);
output(0, 24) <= input(24);
output(0, 25) <= input(25);
output(0, 26) <= input(26);
output(0, 27) <= input(27);
output(0, 28) <= input(28);
output(0, 29) <= input(29);
output(0, 30) <= input(30);
output(0, 31) <= input(31);
output(0, 32) <= input(32);
output(0, 33) <= input(0);
output(0, 34) <= input(1);
output(0, 35) <= input(2);
output(0, 36) <= input(3);
output(0, 37) <= input(4);
output(0, 38) <= input(5);
output(0, 39) <= input(6);
output(0, 40) <= input(7);
output(0, 41) <= input(8);
output(0, 42) <= input(9);
output(0, 43) <= input(10);
output(0, 44) <= input(11);
output(0, 45) <= input(12);
output(0, 46) <= input(13);
output(0, 47) <= input(14);
output(0, 48) <= input(33);
output(0, 49) <= input(16);
output(0, 50) <= input(17);
output(0, 51) <= input(18);
output(0, 52) <= input(19);
output(0, 53) <= input(20);
output(0, 54) <= input(21);
output(0, 55) <= input(22);
output(0, 56) <= input(23);
output(0, 57) <= input(24);
output(0, 58) <= input(25);
output(0, 59) <= input(26);
output(0, 60) <= input(27);
output(0, 61) <= input(28);
output(0, 62) <= input(29);
output(0, 63) <= input(30);
output(0, 64) <= input(34);
output(0, 65) <= input(32);
output(0, 66) <= input(0);
output(0, 67) <= input(1);
output(0, 68) <= input(2);
output(0, 69) <= input(3);
output(0, 70) <= input(4);
output(0, 71) <= input(5);
output(0, 72) <= input(6);
output(0, 73) <= input(7);
output(0, 74) <= input(8);
output(0, 75) <= input(9);
output(0, 76) <= input(10);
output(0, 77) <= input(11);
output(0, 78) <= input(12);
output(0, 79) <= input(13);
output(0, 80) <= input(35);
output(0, 81) <= input(33);
output(0, 82) <= input(16);
output(0, 83) <= input(17);
output(0, 84) <= input(18);
output(0, 85) <= input(19);
output(0, 86) <= input(20);
output(0, 87) <= input(21);
output(0, 88) <= input(22);
output(0, 89) <= input(23);
output(0, 90) <= input(24);
output(0, 91) <= input(25);
output(0, 92) <= input(26);
output(0, 93) <= input(27);
output(0, 94) <= input(28);
output(0, 95) <= input(29);
output(0, 96) <= input(36);
output(0, 97) <= input(34);
output(0, 98) <= input(32);
output(0, 99) <= input(0);
output(0, 100) <= input(1);
output(0, 101) <= input(2);
output(0, 102) <= input(3);
output(0, 103) <= input(4);
output(0, 104) <= input(5);
output(0, 105) <= input(6);
output(0, 106) <= input(7);
output(0, 107) <= input(8);
output(0, 108) <= input(9);
output(0, 109) <= input(10);
output(0, 110) <= input(11);
output(0, 111) <= input(12);
output(0, 112) <= input(37);
output(0, 113) <= input(35);
output(0, 114) <= input(33);
output(0, 115) <= input(16);
output(0, 116) <= input(17);
output(0, 117) <= input(18);
output(0, 118) <= input(19);
output(0, 119) <= input(20);
output(0, 120) <= input(21);
output(0, 121) <= input(22);
output(0, 122) <= input(23);
output(0, 123) <= input(24);
output(0, 124) <= input(25);
output(0, 125) <= input(26);
output(0, 126) <= input(27);
output(0, 127) <= input(28);
output(0, 128) <= input(38);
output(0, 129) <= input(36);
output(0, 130) <= input(34);
output(0, 131) <= input(32);
output(0, 132) <= input(0);
output(0, 133) <= input(1);
output(0, 134) <= input(2);
output(0, 135) <= input(3);
output(0, 136) <= input(4);
output(0, 137) <= input(5);
output(0, 138) <= input(6);
output(0, 139) <= input(7);
output(0, 140) <= input(8);
output(0, 141) <= input(9);
output(0, 142) <= input(10);
output(0, 143) <= input(11);
output(0, 144) <= input(39);
output(0, 145) <= input(37);
output(0, 146) <= input(35);
output(0, 147) <= input(33);
output(0, 148) <= input(16);
output(0, 149) <= input(17);
output(0, 150) <= input(18);
output(0, 151) <= input(19);
output(0, 152) <= input(20);
output(0, 153) <= input(21);
output(0, 154) <= input(22);
output(0, 155) <= input(23);
output(0, 156) <= input(24);
output(0, 157) <= input(25);
output(0, 158) <= input(26);
output(0, 159) <= input(27);
output(0, 160) <= input(40);
output(0, 161) <= input(38);
output(0, 162) <= input(36);
output(0, 163) <= input(34);
output(0, 164) <= input(32);
output(0, 165) <= input(0);
output(0, 166) <= input(1);
output(0, 167) <= input(2);
output(0, 168) <= input(3);
output(0, 169) <= input(4);
output(0, 170) <= input(5);
output(0, 171) <= input(6);
output(0, 172) <= input(7);
output(0, 173) <= input(8);
output(0, 174) <= input(9);
output(0, 175) <= input(10);
output(0, 176) <= input(41);
output(0, 177) <= input(39);
output(0, 178) <= input(37);
output(0, 179) <= input(35);
output(0, 180) <= input(33);
output(0, 181) <= input(16);
output(0, 182) <= input(17);
output(0, 183) <= input(18);
output(0, 184) <= input(19);
output(0, 185) <= input(20);
output(0, 186) <= input(21);
output(0, 187) <= input(22);
output(0, 188) <= input(23);
output(0, 189) <= input(24);
output(0, 190) <= input(25);
output(0, 191) <= input(26);
output(0, 192) <= input(42);
output(0, 193) <= input(40);
output(0, 194) <= input(38);
output(0, 195) <= input(36);
output(0, 196) <= input(34);
output(0, 197) <= input(32);
output(0, 198) <= input(0);
output(0, 199) <= input(1);
output(0, 200) <= input(2);
output(0, 201) <= input(3);
output(0, 202) <= input(4);
output(0, 203) <= input(5);
output(0, 204) <= input(6);
output(0, 205) <= input(7);
output(0, 206) <= input(8);
output(0, 207) <= input(9);
output(0, 208) <= input(43);
output(0, 209) <= input(41);
output(0, 210) <= input(39);
output(0, 211) <= input(37);
output(0, 212) <= input(35);
output(0, 213) <= input(33);
output(0, 214) <= input(16);
output(0, 215) <= input(17);
output(0, 216) <= input(18);
output(0, 217) <= input(19);
output(0, 218) <= input(20);
output(0, 219) <= input(21);
output(0, 220) <= input(22);
output(0, 221) <= input(23);
output(0, 222) <= input(24);
output(0, 223) <= input(25);
output(0, 224) <= input(44);
output(0, 225) <= input(42);
output(0, 226) <= input(40);
output(0, 227) <= input(38);
output(0, 228) <= input(36);
output(0, 229) <= input(34);
output(0, 230) <= input(32);
output(0, 231) <= input(0);
output(0, 232) <= input(1);
output(0, 233) <= input(2);
output(0, 234) <= input(3);
output(0, 235) <= input(4);
output(0, 236) <= input(5);
output(0, 237) <= input(6);
output(0, 238) <= input(7);
output(0, 239) <= input(8);
output(0, 240) <= input(45);
output(0, 241) <= input(43);
output(0, 242) <= input(41);
output(0, 243) <= input(39);
output(0, 244) <= input(37);
output(0, 245) <= input(35);
output(0, 246) <= input(33);
output(0, 247) <= input(16);
output(0, 248) <= input(17);
output(0, 249) <= input(18);
output(0, 250) <= input(19);
output(0, 251) <= input(20);
output(0, 252) <= input(21);
output(0, 253) <= input(22);
output(0, 254) <= input(23);
output(0, 255) <= input(24);
output(1, 0) <= input(16);
output(1, 1) <= input(17);
output(1, 2) <= input(18);
output(1, 3) <= input(19);
output(1, 4) <= input(20);
output(1, 5) <= input(21);
output(1, 6) <= input(22);
output(1, 7) <= input(23);
output(1, 8) <= input(24);
output(1, 9) <= input(25);
output(1, 10) <= input(26);
output(1, 11) <= input(27);
output(1, 12) <= input(28);
output(1, 13) <= input(29);
output(1, 14) <= input(30);
output(1, 15) <= input(31);
output(1, 16) <= input(32);
output(1, 17) <= input(0);
output(1, 18) <= input(1);
output(1, 19) <= input(2);
output(1, 20) <= input(3);
output(1, 21) <= input(4);
output(1, 22) <= input(5);
output(1, 23) <= input(6);
output(1, 24) <= input(7);
output(1, 25) <= input(8);
output(1, 26) <= input(9);
output(1, 27) <= input(10);
output(1, 28) <= input(11);
output(1, 29) <= input(12);
output(1, 30) <= input(13);
output(1, 31) <= input(14);
output(1, 32) <= input(33);
output(1, 33) <= input(16);
output(1, 34) <= input(17);
output(1, 35) <= input(18);
output(1, 36) <= input(19);
output(1, 37) <= input(20);
output(1, 38) <= input(21);
output(1, 39) <= input(22);
output(1, 40) <= input(23);
output(1, 41) <= input(24);
output(1, 42) <= input(25);
output(1, 43) <= input(26);
output(1, 44) <= input(27);
output(1, 45) <= input(28);
output(1, 46) <= input(29);
output(1, 47) <= input(30);
output(1, 48) <= input(34);
output(1, 49) <= input(32);
output(1, 50) <= input(0);
output(1, 51) <= input(1);
output(1, 52) <= input(2);
output(1, 53) <= input(3);
output(1, 54) <= input(4);
output(1, 55) <= input(5);
output(1, 56) <= input(6);
output(1, 57) <= input(7);
output(1, 58) <= input(8);
output(1, 59) <= input(9);
output(1, 60) <= input(10);
output(1, 61) <= input(11);
output(1, 62) <= input(12);
output(1, 63) <= input(13);
output(1, 64) <= input(35);
output(1, 65) <= input(33);
output(1, 66) <= input(16);
output(1, 67) <= input(17);
output(1, 68) <= input(18);
output(1, 69) <= input(19);
output(1, 70) <= input(20);
output(1, 71) <= input(21);
output(1, 72) <= input(22);
output(1, 73) <= input(23);
output(1, 74) <= input(24);
output(1, 75) <= input(25);
output(1, 76) <= input(26);
output(1, 77) <= input(27);
output(1, 78) <= input(28);
output(1, 79) <= input(29);
output(1, 80) <= input(36);
output(1, 81) <= input(34);
output(1, 82) <= input(32);
output(1, 83) <= input(0);
output(1, 84) <= input(1);
output(1, 85) <= input(2);
output(1, 86) <= input(3);
output(1, 87) <= input(4);
output(1, 88) <= input(5);
output(1, 89) <= input(6);
output(1, 90) <= input(7);
output(1, 91) <= input(8);
output(1, 92) <= input(9);
output(1, 93) <= input(10);
output(1, 94) <= input(11);
output(1, 95) <= input(12);
output(1, 96) <= input(37);
output(1, 97) <= input(35);
output(1, 98) <= input(33);
output(1, 99) <= input(16);
output(1, 100) <= input(17);
output(1, 101) <= input(18);
output(1, 102) <= input(19);
output(1, 103) <= input(20);
output(1, 104) <= input(21);
output(1, 105) <= input(22);
output(1, 106) <= input(23);
output(1, 107) <= input(24);
output(1, 108) <= input(25);
output(1, 109) <= input(26);
output(1, 110) <= input(27);
output(1, 111) <= input(28);
output(1, 112) <= input(38);
output(1, 113) <= input(36);
output(1, 114) <= input(34);
output(1, 115) <= input(32);
output(1, 116) <= input(0);
output(1, 117) <= input(1);
output(1, 118) <= input(2);
output(1, 119) <= input(3);
output(1, 120) <= input(4);
output(1, 121) <= input(5);
output(1, 122) <= input(6);
output(1, 123) <= input(7);
output(1, 124) <= input(8);
output(1, 125) <= input(9);
output(1, 126) <= input(10);
output(1, 127) <= input(11);
output(1, 128) <= input(40);
output(1, 129) <= input(38);
output(1, 130) <= input(36);
output(1, 131) <= input(34);
output(1, 132) <= input(32);
output(1, 133) <= input(0);
output(1, 134) <= input(1);
output(1, 135) <= input(2);
output(1, 136) <= input(3);
output(1, 137) <= input(4);
output(1, 138) <= input(5);
output(1, 139) <= input(6);
output(1, 140) <= input(7);
output(1, 141) <= input(8);
output(1, 142) <= input(9);
output(1, 143) <= input(10);
output(1, 144) <= input(41);
output(1, 145) <= input(39);
output(1, 146) <= input(37);
output(1, 147) <= input(35);
output(1, 148) <= input(33);
output(1, 149) <= input(16);
output(1, 150) <= input(17);
output(1, 151) <= input(18);
output(1, 152) <= input(19);
output(1, 153) <= input(20);
output(1, 154) <= input(21);
output(1, 155) <= input(22);
output(1, 156) <= input(23);
output(1, 157) <= input(24);
output(1, 158) <= input(25);
output(1, 159) <= input(26);
output(1, 160) <= input(42);
output(1, 161) <= input(40);
output(1, 162) <= input(38);
output(1, 163) <= input(36);
output(1, 164) <= input(34);
output(1, 165) <= input(32);
output(1, 166) <= input(0);
output(1, 167) <= input(1);
output(1, 168) <= input(2);
output(1, 169) <= input(3);
output(1, 170) <= input(4);
output(1, 171) <= input(5);
output(1, 172) <= input(6);
output(1, 173) <= input(7);
output(1, 174) <= input(8);
output(1, 175) <= input(9);
output(1, 176) <= input(43);
output(1, 177) <= input(41);
output(1, 178) <= input(39);
output(1, 179) <= input(37);
output(1, 180) <= input(35);
output(1, 181) <= input(33);
output(1, 182) <= input(16);
output(1, 183) <= input(17);
output(1, 184) <= input(18);
output(1, 185) <= input(19);
output(1, 186) <= input(20);
output(1, 187) <= input(21);
output(1, 188) <= input(22);
output(1, 189) <= input(23);
output(1, 190) <= input(24);
output(1, 191) <= input(25);
output(1, 192) <= input(44);
output(1, 193) <= input(42);
output(1, 194) <= input(40);
output(1, 195) <= input(38);
output(1, 196) <= input(36);
output(1, 197) <= input(34);
output(1, 198) <= input(32);
output(1, 199) <= input(0);
output(1, 200) <= input(1);
output(1, 201) <= input(2);
output(1, 202) <= input(3);
output(1, 203) <= input(4);
output(1, 204) <= input(5);
output(1, 205) <= input(6);
output(1, 206) <= input(7);
output(1, 207) <= input(8);
output(1, 208) <= input(45);
output(1, 209) <= input(43);
output(1, 210) <= input(41);
output(1, 211) <= input(39);
output(1, 212) <= input(37);
output(1, 213) <= input(35);
output(1, 214) <= input(33);
output(1, 215) <= input(16);
output(1, 216) <= input(17);
output(1, 217) <= input(18);
output(1, 218) <= input(19);
output(1, 219) <= input(20);
output(1, 220) <= input(21);
output(1, 221) <= input(22);
output(1, 222) <= input(23);
output(1, 223) <= input(24);
output(1, 224) <= input(46);
output(1, 225) <= input(44);
output(1, 226) <= input(42);
output(1, 227) <= input(40);
output(1, 228) <= input(38);
output(1, 229) <= input(36);
output(1, 230) <= input(34);
output(1, 231) <= input(32);
output(1, 232) <= input(0);
output(1, 233) <= input(1);
output(1, 234) <= input(2);
output(1, 235) <= input(3);
output(1, 236) <= input(4);
output(1, 237) <= input(5);
output(1, 238) <= input(6);
output(1, 239) <= input(7);
output(1, 240) <= input(47);
output(1, 241) <= input(45);
output(1, 242) <= input(43);
output(1, 243) <= input(41);
output(1, 244) <= input(39);
output(1, 245) <= input(37);
output(1, 246) <= input(35);
output(1, 247) <= input(33);
output(1, 248) <= input(16);
output(1, 249) <= input(17);
output(1, 250) <= input(18);
output(1, 251) <= input(19);
output(1, 252) <= input(20);
output(1, 253) <= input(21);
output(1, 254) <= input(22);
output(1, 255) <= input(23);
when "0110" =>
output(0, 0) <= input(0);
output(0, 1) <= input(1);
output(0, 2) <= input(2);
output(0, 3) <= input(3);
output(0, 4) <= input(4);
output(0, 5) <= input(5);
output(0, 6) <= input(6);
output(0, 7) <= input(7);
output(0, 8) <= input(8);
output(0, 9) <= input(9);
output(0, 10) <= input(10);
output(0, 11) <= input(11);
output(0, 12) <= input(12);
output(0, 13) <= input(13);
output(0, 14) <= input(14);
output(0, 15) <= input(15);
output(0, 16) <= input(16);
output(0, 17) <= input(17);
output(0, 18) <= input(18);
output(0, 19) <= input(19);
output(0, 20) <= input(20);
output(0, 21) <= input(21);
output(0, 22) <= input(22);
output(0, 23) <= input(23);
output(0, 24) <= input(24);
output(0, 25) <= input(25);
output(0, 26) <= input(26);
output(0, 27) <= input(27);
output(0, 28) <= input(28);
output(0, 29) <= input(29);
output(0, 30) <= input(30);
output(0, 31) <= input(31);
output(0, 32) <= input(32);
output(0, 33) <= input(0);
output(0, 34) <= input(1);
output(0, 35) <= input(2);
output(0, 36) <= input(3);
output(0, 37) <= input(4);
output(0, 38) <= input(5);
output(0, 39) <= input(6);
output(0, 40) <= input(7);
output(0, 41) <= input(8);
output(0, 42) <= input(9);
output(0, 43) <= input(10);
output(0, 44) <= input(11);
output(0, 45) <= input(12);
output(0, 46) <= input(13);
output(0, 47) <= input(14);
output(0, 48) <= input(33);
output(0, 49) <= input(16);
output(0, 50) <= input(17);
output(0, 51) <= input(18);
output(0, 52) <= input(19);
output(0, 53) <= input(20);
output(0, 54) <= input(21);
output(0, 55) <= input(22);
output(0, 56) <= input(23);
output(0, 57) <= input(24);
output(0, 58) <= input(25);
output(0, 59) <= input(26);
output(0, 60) <= input(27);
output(0, 61) <= input(28);
output(0, 62) <= input(29);
output(0, 63) <= input(30);
output(0, 64) <= input(34);
output(0, 65) <= input(33);
output(0, 66) <= input(16);
output(0, 67) <= input(17);
output(0, 68) <= input(18);
output(0, 69) <= input(19);
output(0, 70) <= input(20);
output(0, 71) <= input(21);
output(0, 72) <= input(22);
output(0, 73) <= input(23);
output(0, 74) <= input(24);
output(0, 75) <= input(25);
output(0, 76) <= input(26);
output(0, 77) <= input(27);
output(0, 78) <= input(28);
output(0, 79) <= input(29);
output(0, 80) <= input(35);
output(0, 81) <= input(36);
output(0, 82) <= input(32);
output(0, 83) <= input(0);
output(0, 84) <= input(1);
output(0, 85) <= input(2);
output(0, 86) <= input(3);
output(0, 87) <= input(4);
output(0, 88) <= input(5);
output(0, 89) <= input(6);
output(0, 90) <= input(7);
output(0, 91) <= input(8);
output(0, 92) <= input(9);
output(0, 93) <= input(10);
output(0, 94) <= input(11);
output(0, 95) <= input(12);
output(0, 96) <= input(37);
output(0, 97) <= input(34);
output(0, 98) <= input(33);
output(0, 99) <= input(16);
output(0, 100) <= input(17);
output(0, 101) <= input(18);
output(0, 102) <= input(19);
output(0, 103) <= input(20);
output(0, 104) <= input(21);
output(0, 105) <= input(22);
output(0, 106) <= input(23);
output(0, 107) <= input(24);
output(0, 108) <= input(25);
output(0, 109) <= input(26);
output(0, 110) <= input(27);
output(0, 111) <= input(28);
output(0, 112) <= input(38);
output(0, 113) <= input(35);
output(0, 114) <= input(36);
output(0, 115) <= input(32);
output(0, 116) <= input(0);
output(0, 117) <= input(1);
output(0, 118) <= input(2);
output(0, 119) <= input(3);
output(0, 120) <= input(4);
output(0, 121) <= input(5);
output(0, 122) <= input(6);
output(0, 123) <= input(7);
output(0, 124) <= input(8);
output(0, 125) <= input(9);
output(0, 126) <= input(10);
output(0, 127) <= input(11);
output(0, 128) <= input(39);
output(0, 129) <= input(38);
output(0, 130) <= input(35);
output(0, 131) <= input(36);
output(0, 132) <= input(32);
output(0, 133) <= input(0);
output(0, 134) <= input(1);
output(0, 135) <= input(2);
output(0, 136) <= input(3);
output(0, 137) <= input(4);
output(0, 138) <= input(5);
output(0, 139) <= input(6);
output(0, 140) <= input(7);
output(0, 141) <= input(8);
output(0, 142) <= input(9);
output(0, 143) <= input(10);
output(0, 144) <= input(40);
output(0, 145) <= input(41);
output(0, 146) <= input(37);
output(0, 147) <= input(34);
output(0, 148) <= input(33);
output(0, 149) <= input(16);
output(0, 150) <= input(17);
output(0, 151) <= input(18);
output(0, 152) <= input(19);
output(0, 153) <= input(20);
output(0, 154) <= input(21);
output(0, 155) <= input(22);
output(0, 156) <= input(23);
output(0, 157) <= input(24);
output(0, 158) <= input(25);
output(0, 159) <= input(26);
output(0, 160) <= input(42);
output(0, 161) <= input(39);
output(0, 162) <= input(38);
output(0, 163) <= input(35);
output(0, 164) <= input(36);
output(0, 165) <= input(32);
output(0, 166) <= input(0);
output(0, 167) <= input(1);
output(0, 168) <= input(2);
output(0, 169) <= input(3);
output(0, 170) <= input(4);
output(0, 171) <= input(5);
output(0, 172) <= input(6);
output(0, 173) <= input(7);
output(0, 174) <= input(8);
output(0, 175) <= input(9);
output(0, 176) <= input(43);
output(0, 177) <= input(40);
output(0, 178) <= input(41);
output(0, 179) <= input(37);
output(0, 180) <= input(34);
output(0, 181) <= input(33);
output(0, 182) <= input(16);
output(0, 183) <= input(17);
output(0, 184) <= input(18);
output(0, 185) <= input(19);
output(0, 186) <= input(20);
output(0, 187) <= input(21);
output(0, 188) <= input(22);
output(0, 189) <= input(23);
output(0, 190) <= input(24);
output(0, 191) <= input(25);
output(0, 192) <= input(44);
output(0, 193) <= input(43);
output(0, 194) <= input(40);
output(0, 195) <= input(41);
output(0, 196) <= input(37);
output(0, 197) <= input(34);
output(0, 198) <= input(33);
output(0, 199) <= input(16);
output(0, 200) <= input(17);
output(0, 201) <= input(18);
output(0, 202) <= input(19);
output(0, 203) <= input(20);
output(0, 204) <= input(21);
output(0, 205) <= input(22);
output(0, 206) <= input(23);
output(0, 207) <= input(24);
output(0, 208) <= input(45);
output(0, 209) <= input(46);
output(0, 210) <= input(42);
output(0, 211) <= input(39);
output(0, 212) <= input(38);
output(0, 213) <= input(35);
output(0, 214) <= input(36);
output(0, 215) <= input(32);
output(0, 216) <= input(0);
output(0, 217) <= input(1);
output(0, 218) <= input(2);
output(0, 219) <= input(3);
output(0, 220) <= input(4);
output(0, 221) <= input(5);
output(0, 222) <= input(6);
output(0, 223) <= input(7);
output(0, 224) <= input(47);
output(0, 225) <= input(44);
output(0, 226) <= input(43);
output(0, 227) <= input(40);
output(0, 228) <= input(41);
output(0, 229) <= input(37);
output(0, 230) <= input(34);
output(0, 231) <= input(33);
output(0, 232) <= input(16);
output(0, 233) <= input(17);
output(0, 234) <= input(18);
output(0, 235) <= input(19);
output(0, 236) <= input(20);
output(0, 237) <= input(21);
output(0, 238) <= input(22);
output(0, 239) <= input(23);
output(0, 240) <= input(48);
output(0, 241) <= input(45);
output(0, 242) <= input(46);
output(0, 243) <= input(42);
output(0, 244) <= input(39);
output(0, 245) <= input(38);
output(0, 246) <= input(35);
output(0, 247) <= input(36);
output(0, 248) <= input(32);
output(0, 249) <= input(0);
output(0, 250) <= input(1);
output(0, 251) <= input(2);
output(0, 252) <= input(3);
output(0, 253) <= input(4);
output(0, 254) <= input(5);
output(0, 255) <= input(6);
output(1, 0) <= input(0);
output(1, 1) <= input(1);
output(1, 2) <= input(2);
output(1, 3) <= input(3);
output(1, 4) <= input(4);
output(1, 5) <= input(5);
output(1, 6) <= input(6);
output(1, 7) <= input(7);
output(1, 8) <= input(8);
output(1, 9) <= input(9);
output(1, 10) <= input(10);
output(1, 11) <= input(11);
output(1, 12) <= input(12);
output(1, 13) <= input(13);
output(1, 14) <= input(14);
output(1, 15) <= input(15);
output(1, 16) <= input(16);
output(1, 17) <= input(17);
output(1, 18) <= input(18);
output(1, 19) <= input(19);
output(1, 20) <= input(20);
output(1, 21) <= input(21);
output(1, 22) <= input(22);
output(1, 23) <= input(23);
output(1, 24) <= input(24);
output(1, 25) <= input(25);
output(1, 26) <= input(26);
output(1, 27) <= input(27);
output(1, 28) <= input(28);
output(1, 29) <= input(29);
output(1, 30) <= input(30);
output(1, 31) <= input(31);
output(1, 32) <= input(33);
output(1, 33) <= input(16);
output(1, 34) <= input(17);
output(1, 35) <= input(18);
output(1, 36) <= input(19);
output(1, 37) <= input(20);
output(1, 38) <= input(21);
output(1, 39) <= input(22);
output(1, 40) <= input(23);
output(1, 41) <= input(24);
output(1, 42) <= input(25);
output(1, 43) <= input(26);
output(1, 44) <= input(27);
output(1, 45) <= input(28);
output(1, 46) <= input(29);
output(1, 47) <= input(30);
output(1, 48) <= input(36);
output(1, 49) <= input(32);
output(1, 50) <= input(0);
output(1, 51) <= input(1);
output(1, 52) <= input(2);
output(1, 53) <= input(3);
output(1, 54) <= input(4);
output(1, 55) <= input(5);
output(1, 56) <= input(6);
output(1, 57) <= input(7);
output(1, 58) <= input(8);
output(1, 59) <= input(9);
output(1, 60) <= input(10);
output(1, 61) <= input(11);
output(1, 62) <= input(12);
output(1, 63) <= input(13);
output(1, 64) <= input(35);
output(1, 65) <= input(36);
output(1, 66) <= input(32);
output(1, 67) <= input(0);
output(1, 68) <= input(1);
output(1, 69) <= input(2);
output(1, 70) <= input(3);
output(1, 71) <= input(4);
output(1, 72) <= input(5);
output(1, 73) <= input(6);
output(1, 74) <= input(7);
output(1, 75) <= input(8);
output(1, 76) <= input(9);
output(1, 77) <= input(10);
output(1, 78) <= input(11);
output(1, 79) <= input(12);
output(1, 80) <= input(37);
output(1, 81) <= input(34);
output(1, 82) <= input(33);
output(1, 83) <= input(16);
output(1, 84) <= input(17);
output(1, 85) <= input(18);
output(1, 86) <= input(19);
output(1, 87) <= input(20);
output(1, 88) <= input(21);
output(1, 89) <= input(22);
output(1, 90) <= input(23);
output(1, 91) <= input(24);
output(1, 92) <= input(25);
output(1, 93) <= input(26);
output(1, 94) <= input(27);
output(1, 95) <= input(28);
output(1, 96) <= input(41);
output(1, 97) <= input(37);
output(1, 98) <= input(34);
output(1, 99) <= input(33);
output(1, 100) <= input(16);
output(1, 101) <= input(17);
output(1, 102) <= input(18);
output(1, 103) <= input(19);
output(1, 104) <= input(20);
output(1, 105) <= input(21);
output(1, 106) <= input(22);
output(1, 107) <= input(23);
output(1, 108) <= input(24);
output(1, 109) <= input(25);
output(1, 110) <= input(26);
output(1, 111) <= input(27);
output(1, 112) <= input(39);
output(1, 113) <= input(38);
output(1, 114) <= input(35);
output(1, 115) <= input(36);
output(1, 116) <= input(32);
output(1, 117) <= input(0);
output(1, 118) <= input(1);
output(1, 119) <= input(2);
output(1, 120) <= input(3);
output(1, 121) <= input(4);
output(1, 122) <= input(5);
output(1, 123) <= input(6);
output(1, 124) <= input(7);
output(1, 125) <= input(8);
output(1, 126) <= input(9);
output(1, 127) <= input(10);
output(1, 128) <= input(40);
output(1, 129) <= input(41);
output(1, 130) <= input(37);
output(1, 131) <= input(34);
output(1, 132) <= input(33);
output(1, 133) <= input(16);
output(1, 134) <= input(17);
output(1, 135) <= input(18);
output(1, 136) <= input(19);
output(1, 137) <= input(20);
output(1, 138) <= input(21);
output(1, 139) <= input(22);
output(1, 140) <= input(23);
output(1, 141) <= input(24);
output(1, 142) <= input(25);
output(1, 143) <= input(26);
output(1, 144) <= input(43);
output(1, 145) <= input(40);
output(1, 146) <= input(41);
output(1, 147) <= input(37);
output(1, 148) <= input(34);
output(1, 149) <= input(33);
output(1, 150) <= input(16);
output(1, 151) <= input(17);
output(1, 152) <= input(18);
output(1, 153) <= input(19);
output(1, 154) <= input(20);
output(1, 155) <= input(21);
output(1, 156) <= input(22);
output(1, 157) <= input(23);
output(1, 158) <= input(24);
output(1, 159) <= input(25);
output(1, 160) <= input(46);
output(1, 161) <= input(42);
output(1, 162) <= input(39);
output(1, 163) <= input(38);
output(1, 164) <= input(35);
output(1, 165) <= input(36);
output(1, 166) <= input(32);
output(1, 167) <= input(0);
output(1, 168) <= input(1);
output(1, 169) <= input(2);
output(1, 170) <= input(3);
output(1, 171) <= input(4);
output(1, 172) <= input(5);
output(1, 173) <= input(6);
output(1, 174) <= input(7);
output(1, 175) <= input(8);
output(1, 176) <= input(45);
output(1, 177) <= input(46);
output(1, 178) <= input(42);
output(1, 179) <= input(39);
output(1, 180) <= input(38);
output(1, 181) <= input(35);
output(1, 182) <= input(36);
output(1, 183) <= input(32);
output(1, 184) <= input(0);
output(1, 185) <= input(1);
output(1, 186) <= input(2);
output(1, 187) <= input(3);
output(1, 188) <= input(4);
output(1, 189) <= input(5);
output(1, 190) <= input(6);
output(1, 191) <= input(7);
output(1, 192) <= input(47);
output(1, 193) <= input(44);
output(1, 194) <= input(43);
output(1, 195) <= input(40);
output(1, 196) <= input(41);
output(1, 197) <= input(37);
output(1, 198) <= input(34);
output(1, 199) <= input(33);
output(1, 200) <= input(16);
output(1, 201) <= input(17);
output(1, 202) <= input(18);
output(1, 203) <= input(19);
output(1, 204) <= input(20);
output(1, 205) <= input(21);
output(1, 206) <= input(22);
output(1, 207) <= input(23);
output(1, 208) <= input(49);
output(1, 209) <= input(47);
output(1, 210) <= input(44);
output(1, 211) <= input(43);
output(1, 212) <= input(40);
output(1, 213) <= input(41);
output(1, 214) <= input(37);
output(1, 215) <= input(34);
output(1, 216) <= input(33);
output(1, 217) <= input(16);
output(1, 218) <= input(17);
output(1, 219) <= input(18);
output(1, 220) <= input(19);
output(1, 221) <= input(20);
output(1, 222) <= input(21);
output(1, 223) <= input(22);
output(1, 224) <= input(50);
output(1, 225) <= input(48);
output(1, 226) <= input(45);
output(1, 227) <= input(46);
output(1, 228) <= input(42);
output(1, 229) <= input(39);
output(1, 230) <= input(38);
output(1, 231) <= input(35);
output(1, 232) <= input(36);
output(1, 233) <= input(32);
output(1, 234) <= input(0);
output(1, 235) <= input(1);
output(1, 236) <= input(2);
output(1, 237) <= input(3);
output(1, 238) <= input(4);
output(1, 239) <= input(5);
output(1, 240) <= input(51);
output(1, 241) <= input(49);
output(1, 242) <= input(47);
output(1, 243) <= input(44);
output(1, 244) <= input(43);
output(1, 245) <= input(40);
output(1, 246) <= input(41);
output(1, 247) <= input(37);
output(1, 248) <= input(34);
output(1, 249) <= input(33);
output(1, 250) <= input(16);
output(1, 251) <= input(17);
output(1, 252) <= input(18);
output(1, 253) <= input(19);
output(1, 254) <= input(20);
output(1, 255) <= input(21);
output(2, 0) <= input(0);
output(2, 1) <= input(1);
output(2, 2) <= input(2);
output(2, 3) <= input(3);
output(2, 4) <= input(4);
output(2, 5) <= input(5);
output(2, 6) <= input(6);
output(2, 7) <= input(7);
output(2, 8) <= input(8);
output(2, 9) <= input(9);
output(2, 10) <= input(10);
output(2, 11) <= input(11);
output(2, 12) <= input(12);
output(2, 13) <= input(13);
output(2, 14) <= input(14);
output(2, 15) <= input(15);
output(2, 16) <= input(32);
output(2, 17) <= input(0);
output(2, 18) <= input(1);
output(2, 19) <= input(2);
output(2, 20) <= input(3);
output(2, 21) <= input(4);
output(2, 22) <= input(5);
output(2, 23) <= input(6);
output(2, 24) <= input(7);
output(2, 25) <= input(8);
output(2, 26) <= input(9);
output(2, 27) <= input(10);
output(2, 28) <= input(11);
output(2, 29) <= input(12);
output(2, 30) <= input(13);
output(2, 31) <= input(14);
output(2, 32) <= input(33);
output(2, 33) <= input(16);
output(2, 34) <= input(17);
output(2, 35) <= input(18);
output(2, 36) <= input(19);
output(2, 37) <= input(20);
output(2, 38) <= input(21);
output(2, 39) <= input(22);
output(2, 40) <= input(23);
output(2, 41) <= input(24);
output(2, 42) <= input(25);
output(2, 43) <= input(26);
output(2, 44) <= input(27);
output(2, 45) <= input(28);
output(2, 46) <= input(29);
output(2, 47) <= input(30);
output(2, 48) <= input(34);
output(2, 49) <= input(33);
output(2, 50) <= input(16);
output(2, 51) <= input(17);
output(2, 52) <= input(18);
output(2, 53) <= input(19);
output(2, 54) <= input(20);
output(2, 55) <= input(21);
output(2, 56) <= input(22);
output(2, 57) <= input(23);
output(2, 58) <= input(24);
output(2, 59) <= input(25);
output(2, 60) <= input(26);
output(2, 61) <= input(27);
output(2, 62) <= input(28);
output(2, 63) <= input(29);
output(2, 64) <= input(37);
output(2, 65) <= input(34);
output(2, 66) <= input(33);
output(2, 67) <= input(16);
output(2, 68) <= input(17);
output(2, 69) <= input(18);
output(2, 70) <= input(19);
output(2, 71) <= input(20);
output(2, 72) <= input(21);
output(2, 73) <= input(22);
output(2, 74) <= input(23);
output(2, 75) <= input(24);
output(2, 76) <= input(25);
output(2, 77) <= input(26);
output(2, 78) <= input(27);
output(2, 79) <= input(28);
output(2, 80) <= input(38);
output(2, 81) <= input(35);
output(2, 82) <= input(36);
output(2, 83) <= input(32);
output(2, 84) <= input(0);
output(2, 85) <= input(1);
output(2, 86) <= input(2);
output(2, 87) <= input(3);
output(2, 88) <= input(4);
output(2, 89) <= input(5);
output(2, 90) <= input(6);
output(2, 91) <= input(7);
output(2, 92) <= input(8);
output(2, 93) <= input(9);
output(2, 94) <= input(10);
output(2, 95) <= input(11);
output(2, 96) <= input(39);
output(2, 97) <= input(38);
output(2, 98) <= input(35);
output(2, 99) <= input(36);
output(2, 100) <= input(32);
output(2, 101) <= input(0);
output(2, 102) <= input(1);
output(2, 103) <= input(2);
output(2, 104) <= input(3);
output(2, 105) <= input(4);
output(2, 106) <= input(5);
output(2, 107) <= input(6);
output(2, 108) <= input(7);
output(2, 109) <= input(8);
output(2, 110) <= input(9);
output(2, 111) <= input(10);
output(2, 112) <= input(40);
output(2, 113) <= input(41);
output(2, 114) <= input(37);
output(2, 115) <= input(34);
output(2, 116) <= input(33);
output(2, 117) <= input(16);
output(2, 118) <= input(17);
output(2, 119) <= input(18);
output(2, 120) <= input(19);
output(2, 121) <= input(20);
output(2, 122) <= input(21);
output(2, 123) <= input(22);
output(2, 124) <= input(23);
output(2, 125) <= input(24);
output(2, 126) <= input(25);
output(2, 127) <= input(26);
output(2, 128) <= input(43);
output(2, 129) <= input(40);
output(2, 130) <= input(41);
output(2, 131) <= input(37);
output(2, 132) <= input(34);
output(2, 133) <= input(33);
output(2, 134) <= input(16);
output(2, 135) <= input(17);
output(2, 136) <= input(18);
output(2, 137) <= input(19);
output(2, 138) <= input(20);
output(2, 139) <= input(21);
output(2, 140) <= input(22);
output(2, 141) <= input(23);
output(2, 142) <= input(24);
output(2, 143) <= input(25);
output(2, 144) <= input(44);
output(2, 145) <= input(43);
output(2, 146) <= input(40);
output(2, 147) <= input(41);
output(2, 148) <= input(37);
output(2, 149) <= input(34);
output(2, 150) <= input(33);
output(2, 151) <= input(16);
output(2, 152) <= input(17);
output(2, 153) <= input(18);
output(2, 154) <= input(19);
output(2, 155) <= input(20);
output(2, 156) <= input(21);
output(2, 157) <= input(22);
output(2, 158) <= input(23);
output(2, 159) <= input(24);
output(2, 160) <= input(45);
output(2, 161) <= input(46);
output(2, 162) <= input(42);
output(2, 163) <= input(39);
output(2, 164) <= input(38);
output(2, 165) <= input(35);
output(2, 166) <= input(36);
output(2, 167) <= input(32);
output(2, 168) <= input(0);
output(2, 169) <= input(1);
output(2, 170) <= input(2);
output(2, 171) <= input(3);
output(2, 172) <= input(4);
output(2, 173) <= input(5);
output(2, 174) <= input(6);
output(2, 175) <= input(7);
output(2, 176) <= input(48);
output(2, 177) <= input(45);
output(2, 178) <= input(46);
output(2, 179) <= input(42);
output(2, 180) <= input(39);
output(2, 181) <= input(38);
output(2, 182) <= input(35);
output(2, 183) <= input(36);
output(2, 184) <= input(32);
output(2, 185) <= input(0);
output(2, 186) <= input(1);
output(2, 187) <= input(2);
output(2, 188) <= input(3);
output(2, 189) <= input(4);
output(2, 190) <= input(5);
output(2, 191) <= input(6);
output(2, 192) <= input(50);
output(2, 193) <= input(48);
output(2, 194) <= input(45);
output(2, 195) <= input(46);
output(2, 196) <= input(42);
output(2, 197) <= input(39);
output(2, 198) <= input(38);
output(2, 199) <= input(35);
output(2, 200) <= input(36);
output(2, 201) <= input(32);
output(2, 202) <= input(0);
output(2, 203) <= input(1);
output(2, 204) <= input(2);
output(2, 205) <= input(3);
output(2, 206) <= input(4);
output(2, 207) <= input(5);
output(2, 208) <= input(51);
output(2, 209) <= input(49);
output(2, 210) <= input(47);
output(2, 211) <= input(44);
output(2, 212) <= input(43);
output(2, 213) <= input(40);
output(2, 214) <= input(41);
output(2, 215) <= input(37);
output(2, 216) <= input(34);
output(2, 217) <= input(33);
output(2, 218) <= input(16);
output(2, 219) <= input(17);
output(2, 220) <= input(18);
output(2, 221) <= input(19);
output(2, 222) <= input(20);
output(2, 223) <= input(21);
output(2, 224) <= input(52);
output(2, 225) <= input(51);
output(2, 226) <= input(49);
output(2, 227) <= input(47);
output(2, 228) <= input(44);
output(2, 229) <= input(43);
output(2, 230) <= input(40);
output(2, 231) <= input(41);
output(2, 232) <= input(37);
output(2, 233) <= input(34);
output(2, 234) <= input(33);
output(2, 235) <= input(16);
output(2, 236) <= input(17);
output(2, 237) <= input(18);
output(2, 238) <= input(19);
output(2, 239) <= input(20);
output(2, 240) <= input(53);
output(2, 241) <= input(54);
output(2, 242) <= input(50);
output(2, 243) <= input(48);
output(2, 244) <= input(45);
output(2, 245) <= input(46);
output(2, 246) <= input(42);
output(2, 247) <= input(39);
output(2, 248) <= input(38);
output(2, 249) <= input(35);
output(2, 250) <= input(36);
output(2, 251) <= input(32);
output(2, 252) <= input(0);
output(2, 253) <= input(1);
output(2, 254) <= input(2);
output(2, 255) <= input(3);
when "0111" =>
output(0, 0) <= input(0);
output(0, 1) <= input(1);
output(0, 2) <= input(2);
output(0, 3) <= input(3);
output(0, 4) <= input(4);
output(0, 5) <= input(5);
output(0, 6) <= input(6);
output(0, 7) <= input(7);
output(0, 8) <= input(8);
output(0, 9) <= input(9);
output(0, 10) <= input(10);
output(0, 11) <= input(11);
output(0, 12) <= input(12);
output(0, 13) <= input(13);
output(0, 14) <= input(14);
output(0, 15) <= input(15);
output(0, 16) <= input(16);
output(0, 17) <= input(0);
output(0, 18) <= input(1);
output(0, 19) <= input(2);
output(0, 20) <= input(3);
output(0, 21) <= input(4);
output(0, 22) <= input(5);
output(0, 23) <= input(6);
output(0, 24) <= input(7);
output(0, 25) <= input(8);
output(0, 26) <= input(9);
output(0, 27) <= input(10);
output(0, 28) <= input(11);
output(0, 29) <= input(12);
output(0, 30) <= input(13);
output(0, 31) <= input(14);
output(0, 32) <= input(17);
output(0, 33) <= input(16);
output(0, 34) <= input(0);
output(0, 35) <= input(1);
output(0, 36) <= input(2);
output(0, 37) <= input(3);
output(0, 38) <= input(4);
output(0, 39) <= input(5);
output(0, 40) <= input(6);
output(0, 41) <= input(7);
output(0, 42) <= input(8);
output(0, 43) <= input(9);
output(0, 44) <= input(10);
output(0, 45) <= input(11);
output(0, 46) <= input(12);
output(0, 47) <= input(13);
output(0, 48) <= input(18);
output(0, 49) <= input(17);
output(0, 50) <= input(16);
output(0, 51) <= input(0);
output(0, 52) <= input(1);
output(0, 53) <= input(2);
output(0, 54) <= input(3);
output(0, 55) <= input(4);
output(0, 56) <= input(5);
output(0, 57) <= input(6);
output(0, 58) <= input(7);
output(0, 59) <= input(8);
output(0, 60) <= input(9);
output(0, 61) <= input(10);
output(0, 62) <= input(11);
output(0, 63) <= input(12);
output(0, 64) <= input(19);
output(0, 65) <= input(18);
output(0, 66) <= input(17);
output(0, 67) <= input(16);
output(0, 68) <= input(0);
output(0, 69) <= input(1);
output(0, 70) <= input(2);
output(0, 71) <= input(3);
output(0, 72) <= input(4);
output(0, 73) <= input(5);
output(0, 74) <= input(6);
output(0, 75) <= input(7);
output(0, 76) <= input(8);
output(0, 77) <= input(9);
output(0, 78) <= input(10);
output(0, 79) <= input(11);
output(0, 80) <= input(20);
output(0, 81) <= input(21);
output(0, 82) <= input(22);
output(0, 83) <= input(23);
output(0, 84) <= input(24);
output(0, 85) <= input(25);
output(0, 86) <= input(26);
output(0, 87) <= input(27);
output(0, 88) <= input(28);
output(0, 89) <= input(29);
output(0, 90) <= input(30);
output(0, 91) <= input(31);
output(0, 92) <= input(32);
output(0, 93) <= input(33);
output(0, 94) <= input(34);
output(0, 95) <= input(35);
output(0, 96) <= input(36);
output(0, 97) <= input(20);
output(0, 98) <= input(21);
output(0, 99) <= input(22);
output(0, 100) <= input(23);
output(0, 101) <= input(24);
output(0, 102) <= input(25);
output(0, 103) <= input(26);
output(0, 104) <= input(27);
output(0, 105) <= input(28);
output(0, 106) <= input(29);
output(0, 107) <= input(30);
output(0, 108) <= input(31);
output(0, 109) <= input(32);
output(0, 110) <= input(33);
output(0, 111) <= input(34);
output(0, 112) <= input(37);
output(0, 113) <= input(36);
output(0, 114) <= input(20);
output(0, 115) <= input(21);
output(0, 116) <= input(22);
output(0, 117) <= input(23);
output(0, 118) <= input(24);
output(0, 119) <= input(25);
output(0, 120) <= input(26);
output(0, 121) <= input(27);
output(0, 122) <= input(28);
output(0, 123) <= input(29);
output(0, 124) <= input(30);
output(0, 125) <= input(31);
output(0, 126) <= input(32);
output(0, 127) <= input(33);
output(0, 128) <= input(38);
output(0, 129) <= input(37);
output(0, 130) <= input(36);
output(0, 131) <= input(20);
output(0, 132) <= input(21);
output(0, 133) <= input(22);
output(0, 134) <= input(23);
output(0, 135) <= input(24);
output(0, 136) <= input(25);
output(0, 137) <= input(26);
output(0, 138) <= input(27);
output(0, 139) <= input(28);
output(0, 140) <= input(29);
output(0, 141) <= input(30);
output(0, 142) <= input(31);
output(0, 143) <= input(32);
output(0, 144) <= input(39);
output(0, 145) <= input(38);
output(0, 146) <= input(37);
output(0, 147) <= input(36);
output(0, 148) <= input(20);
output(0, 149) <= input(21);
output(0, 150) <= input(22);
output(0, 151) <= input(23);
output(0, 152) <= input(24);
output(0, 153) <= input(25);
output(0, 154) <= input(26);
output(0, 155) <= input(27);
output(0, 156) <= input(28);
output(0, 157) <= input(29);
output(0, 158) <= input(30);
output(0, 159) <= input(31);
output(0, 160) <= input(40);
output(0, 161) <= input(41);
output(0, 162) <= input(42);
output(0, 163) <= input(43);
output(0, 164) <= input(44);
output(0, 165) <= input(19);
output(0, 166) <= input(18);
output(0, 167) <= input(17);
output(0, 168) <= input(16);
output(0, 169) <= input(0);
output(0, 170) <= input(1);
output(0, 171) <= input(2);
output(0, 172) <= input(3);
output(0, 173) <= input(4);
output(0, 174) <= input(5);
output(0, 175) <= input(6);
output(0, 176) <= input(45);
output(0, 177) <= input(40);
output(0, 178) <= input(41);
output(0, 179) <= input(42);
output(0, 180) <= input(43);
output(0, 181) <= input(44);
output(0, 182) <= input(19);
output(0, 183) <= input(18);
output(0, 184) <= input(17);
output(0, 185) <= input(16);
output(0, 186) <= input(0);
output(0, 187) <= input(1);
output(0, 188) <= input(2);
output(0, 189) <= input(3);
output(0, 190) <= input(4);
output(0, 191) <= input(5);
output(0, 192) <= input(46);
output(0, 193) <= input(45);
output(0, 194) <= input(40);
output(0, 195) <= input(41);
output(0, 196) <= input(42);
output(0, 197) <= input(43);
output(0, 198) <= input(44);
output(0, 199) <= input(19);
output(0, 200) <= input(18);
output(0, 201) <= input(17);
output(0, 202) <= input(16);
output(0, 203) <= input(0);
output(0, 204) <= input(1);
output(0, 205) <= input(2);
output(0, 206) <= input(3);
output(0, 207) <= input(4);
output(0, 208) <= input(47);
output(0, 209) <= input(46);
output(0, 210) <= input(45);
output(0, 211) <= input(40);
output(0, 212) <= input(41);
output(0, 213) <= input(42);
output(0, 214) <= input(43);
output(0, 215) <= input(44);
output(0, 216) <= input(19);
output(0, 217) <= input(18);
output(0, 218) <= input(17);
output(0, 219) <= input(16);
output(0, 220) <= input(0);
output(0, 221) <= input(1);
output(0, 222) <= input(2);
output(0, 223) <= input(3);
output(0, 224) <= input(48);
output(0, 225) <= input(47);
output(0, 226) <= input(46);
output(0, 227) <= input(45);
output(0, 228) <= input(40);
output(0, 229) <= input(41);
output(0, 230) <= input(42);
output(0, 231) <= input(43);
output(0, 232) <= input(44);
output(0, 233) <= input(19);
output(0, 234) <= input(18);
output(0, 235) <= input(17);
output(0, 236) <= input(16);
output(0, 237) <= input(0);
output(0, 238) <= input(1);
output(0, 239) <= input(2);
output(0, 240) <= input(49);
output(0, 241) <= input(50);
output(0, 242) <= input(51);
output(0, 243) <= input(52);
output(0, 244) <= input(53);
output(0, 245) <= input(39);
output(0, 246) <= input(38);
output(0, 247) <= input(37);
output(0, 248) <= input(36);
output(0, 249) <= input(20);
output(0, 250) <= input(21);
output(0, 251) <= input(22);
output(0, 252) <= input(23);
output(0, 253) <= input(24);
output(0, 254) <= input(25);
output(0, 255) <= input(26);
output(1, 0) <= input(54);
output(1, 1) <= input(55);
output(1, 2) <= input(56);
output(1, 3) <= input(57);
output(1, 4) <= input(58);
output(1, 5) <= input(59);
output(1, 6) <= input(60);
output(1, 7) <= input(61);
output(1, 8) <= input(62);
output(1, 9) <= input(63);
output(1, 10) <= input(64);
output(1, 11) <= input(65);
output(1, 12) <= input(66);
output(1, 13) <= input(67);
output(1, 14) <= input(68);
output(1, 15) <= input(69);
output(1, 16) <= input(70);
output(1, 17) <= input(54);
output(1, 18) <= input(55);
output(1, 19) <= input(56);
output(1, 20) <= input(57);
output(1, 21) <= input(58);
output(1, 22) <= input(59);
output(1, 23) <= input(60);
output(1, 24) <= input(61);
output(1, 25) <= input(62);
output(1, 26) <= input(63);
output(1, 27) <= input(64);
output(1, 28) <= input(65);
output(1, 29) <= input(66);
output(1, 30) <= input(67);
output(1, 31) <= input(68);
output(1, 32) <= input(71);
output(1, 33) <= input(70);
output(1, 34) <= input(54);
output(1, 35) <= input(55);
output(1, 36) <= input(56);
output(1, 37) <= input(57);
output(1, 38) <= input(58);
output(1, 39) <= input(59);
output(1, 40) <= input(60);
output(1, 41) <= input(61);
output(1, 42) <= input(62);
output(1, 43) <= input(63);
output(1, 44) <= input(64);
output(1, 45) <= input(65);
output(1, 46) <= input(66);
output(1, 47) <= input(67);
output(1, 48) <= input(72);
output(1, 49) <= input(71);
output(1, 50) <= input(70);
output(1, 51) <= input(54);
output(1, 52) <= input(55);
output(1, 53) <= input(56);
output(1, 54) <= input(57);
output(1, 55) <= input(58);
output(1, 56) <= input(59);
output(1, 57) <= input(60);
output(1, 58) <= input(61);
output(1, 59) <= input(62);
output(1, 60) <= input(63);
output(1, 61) <= input(64);
output(1, 62) <= input(65);
output(1, 63) <= input(66);
output(1, 64) <= input(73);
output(1, 65) <= input(72);
output(1, 66) <= input(71);
output(1, 67) <= input(70);
output(1, 68) <= input(54);
output(1, 69) <= input(55);
output(1, 70) <= input(56);
output(1, 71) <= input(57);
output(1, 72) <= input(58);
output(1, 73) <= input(59);
output(1, 74) <= input(60);
output(1, 75) <= input(61);
output(1, 76) <= input(62);
output(1, 77) <= input(63);
output(1, 78) <= input(64);
output(1, 79) <= input(65);
output(1, 80) <= input(74);
output(1, 81) <= input(73);
output(1, 82) <= input(72);
output(1, 83) <= input(71);
output(1, 84) <= input(70);
output(1, 85) <= input(54);
output(1, 86) <= input(55);
output(1, 87) <= input(56);
output(1, 88) <= input(57);
output(1, 89) <= input(58);
output(1, 90) <= input(59);
output(1, 91) <= input(60);
output(1, 92) <= input(61);
output(1, 93) <= input(62);
output(1, 94) <= input(63);
output(1, 95) <= input(64);
output(1, 96) <= input(75);
output(1, 97) <= input(74);
output(1, 98) <= input(73);
output(1, 99) <= input(72);
output(1, 100) <= input(71);
output(1, 101) <= input(70);
output(1, 102) <= input(54);
output(1, 103) <= input(55);
output(1, 104) <= input(56);
output(1, 105) <= input(57);
output(1, 106) <= input(58);
output(1, 107) <= input(59);
output(1, 108) <= input(60);
output(1, 109) <= input(61);
output(1, 110) <= input(62);
output(1, 111) <= input(63);
output(1, 112) <= input(76);
output(1, 113) <= input(75);
output(1, 114) <= input(74);
output(1, 115) <= input(73);
output(1, 116) <= input(72);
output(1, 117) <= input(71);
output(1, 118) <= input(70);
output(1, 119) <= input(54);
output(1, 120) <= input(55);
output(1, 121) <= input(56);
output(1, 122) <= input(57);
output(1, 123) <= input(58);
output(1, 124) <= input(59);
output(1, 125) <= input(60);
output(1, 126) <= input(61);
output(1, 127) <= input(62);
output(1, 128) <= input(77);
output(1, 129) <= input(76);
output(1, 130) <= input(75);
output(1, 131) <= input(74);
output(1, 132) <= input(73);
output(1, 133) <= input(72);
output(1, 134) <= input(71);
output(1, 135) <= input(70);
output(1, 136) <= input(54);
output(1, 137) <= input(55);
output(1, 138) <= input(56);
output(1, 139) <= input(57);
output(1, 140) <= input(58);
output(1, 141) <= input(59);
output(1, 142) <= input(60);
output(1, 143) <= input(61);
output(1, 144) <= input(78);
output(1, 145) <= input(77);
output(1, 146) <= input(76);
output(1, 147) <= input(75);
output(1, 148) <= input(74);
output(1, 149) <= input(73);
output(1, 150) <= input(72);
output(1, 151) <= input(71);
output(1, 152) <= input(70);
output(1, 153) <= input(54);
output(1, 154) <= input(55);
output(1, 155) <= input(56);
output(1, 156) <= input(57);
output(1, 157) <= input(58);
output(1, 158) <= input(59);
output(1, 159) <= input(60);
output(1, 160) <= input(79);
output(1, 161) <= input(78);
output(1, 162) <= input(77);
output(1, 163) <= input(76);
output(1, 164) <= input(75);
output(1, 165) <= input(74);
output(1, 166) <= input(73);
output(1, 167) <= input(72);
output(1, 168) <= input(71);
output(1, 169) <= input(70);
output(1, 170) <= input(54);
output(1, 171) <= input(55);
output(1, 172) <= input(56);
output(1, 173) <= input(57);
output(1, 174) <= input(58);
output(1, 175) <= input(59);
output(1, 176) <= input(80);
output(1, 177) <= input(79);
output(1, 178) <= input(78);
output(1, 179) <= input(77);
output(1, 180) <= input(76);
output(1, 181) <= input(75);
output(1, 182) <= input(74);
output(1, 183) <= input(73);
output(1, 184) <= input(72);
output(1, 185) <= input(71);
output(1, 186) <= input(70);
output(1, 187) <= input(54);
output(1, 188) <= input(55);
output(1, 189) <= input(56);
output(1, 190) <= input(57);
output(1, 191) <= input(58);
output(1, 192) <= input(81);
output(1, 193) <= input(80);
output(1, 194) <= input(79);
output(1, 195) <= input(78);
output(1, 196) <= input(77);
output(1, 197) <= input(76);
output(1, 198) <= input(75);
output(1, 199) <= input(74);
output(1, 200) <= input(73);
output(1, 201) <= input(72);
output(1, 202) <= input(71);
output(1, 203) <= input(70);
output(1, 204) <= input(54);
output(1, 205) <= input(55);
output(1, 206) <= input(56);
output(1, 207) <= input(57);
output(1, 208) <= input(82);
output(1, 209) <= input(81);
output(1, 210) <= input(80);
output(1, 211) <= input(79);
output(1, 212) <= input(78);
output(1, 213) <= input(77);
output(1, 214) <= input(76);
output(1, 215) <= input(75);
output(1, 216) <= input(74);
output(1, 217) <= input(73);
output(1, 218) <= input(72);
output(1, 219) <= input(71);
output(1, 220) <= input(70);
output(1, 221) <= input(54);
output(1, 222) <= input(55);
output(1, 223) <= input(56);
output(1, 224) <= input(83);
output(1, 225) <= input(82);
output(1, 226) <= input(81);
output(1, 227) <= input(80);
output(1, 228) <= input(79);
output(1, 229) <= input(78);
output(1, 230) <= input(77);
output(1, 231) <= input(76);
output(1, 232) <= input(75);
output(1, 233) <= input(74);
output(1, 234) <= input(73);
output(1, 235) <= input(72);
output(1, 236) <= input(71);
output(1, 237) <= input(70);
output(1, 238) <= input(54);
output(1, 239) <= input(55);
output(1, 240) <= input(84);
output(1, 241) <= input(83);
output(1, 242) <= input(82);
output(1, 243) <= input(81);
output(1, 244) <= input(80);
output(1, 245) <= input(79);
output(1, 246) <= input(78);
output(1, 247) <= input(77);
output(1, 248) <= input(76);
output(1, 249) <= input(75);
output(1, 250) <= input(74);
output(1, 251) <= input(73);
output(1, 252) <= input(72);
output(1, 253) <= input(71);
output(1, 254) <= input(70);
output(1, 255) <= input(54);
when "1000" =>
output(0, 0) <= input(0);
output(0, 1) <= input(1);
output(0, 2) <= input(2);
output(0, 3) <= input(3);
output(0, 4) <= input(4);
output(0, 5) <= input(5);
output(0, 6) <= input(6);
output(0, 7) <= input(7);
output(0, 8) <= input(8);
output(0, 9) <= input(9);
output(0, 10) <= input(10);
output(0, 11) <= input(11);
output(0, 12) <= input(12);
output(0, 13) <= input(13);
output(0, 14) <= input(14);
output(0, 15) <= input(15);
output(0, 16) <= input(16);
output(0, 17) <= input(0);
output(0, 18) <= input(1);
output(0, 19) <= input(2);
output(0, 20) <= input(3);
output(0, 21) <= input(4);
output(0, 22) <= input(5);
output(0, 23) <= input(6);
output(0, 24) <= input(7);
output(0, 25) <= input(8);
output(0, 26) <= input(9);
output(0, 27) <= input(10);
output(0, 28) <= input(11);
output(0, 29) <= input(12);
output(0, 30) <= input(13);
output(0, 31) <= input(14);
output(0, 32) <= input(17);
output(0, 33) <= input(16);
output(0, 34) <= input(0);
output(0, 35) <= input(1);
output(0, 36) <= input(2);
output(0, 37) <= input(3);
output(0, 38) <= input(4);
output(0, 39) <= input(5);
output(0, 40) <= input(6);
output(0, 41) <= input(7);
output(0, 42) <= input(8);
output(0, 43) <= input(9);
output(0, 44) <= input(10);
output(0, 45) <= input(11);
output(0, 46) <= input(12);
output(0, 47) <= input(13);
output(0, 48) <= input(18);
output(0, 49) <= input(17);
output(0, 50) <= input(16);
output(0, 51) <= input(0);
output(0, 52) <= input(1);
output(0, 53) <= input(2);
output(0, 54) <= input(3);
output(0, 55) <= input(4);
output(0, 56) <= input(5);
output(0, 57) <= input(6);
output(0, 58) <= input(7);
output(0, 59) <= input(8);
output(0, 60) <= input(9);
output(0, 61) <= input(10);
output(0, 62) <= input(11);
output(0, 63) <= input(12);
output(0, 64) <= input(19);
output(0, 65) <= input(18);
output(0, 66) <= input(17);
output(0, 67) <= input(16);
output(0, 68) <= input(0);
output(0, 69) <= input(1);
output(0, 70) <= input(2);
output(0, 71) <= input(3);
output(0, 72) <= input(4);
output(0, 73) <= input(5);
output(0, 74) <= input(6);
output(0, 75) <= input(7);
output(0, 76) <= input(8);
output(0, 77) <= input(9);
output(0, 78) <= input(10);
output(0, 79) <= input(11);
output(0, 80) <= input(20);
output(0, 81) <= input(21);
output(0, 82) <= input(22);
output(0, 83) <= input(23);
output(0, 84) <= input(24);
output(0, 85) <= input(25);
output(0, 86) <= input(26);
output(0, 87) <= input(27);
output(0, 88) <= input(28);
output(0, 89) <= input(29);
output(0, 90) <= input(30);
output(0, 91) <= input(31);
output(0, 92) <= input(32);
output(0, 93) <= input(33);
output(0, 94) <= input(34);
output(0, 95) <= input(35);
output(0, 96) <= input(36);
output(0, 97) <= input(20);
output(0, 98) <= input(21);
output(0, 99) <= input(22);
output(0, 100) <= input(23);
output(0, 101) <= input(24);
output(0, 102) <= input(25);
output(0, 103) <= input(26);
output(0, 104) <= input(27);
output(0, 105) <= input(28);
output(0, 106) <= input(29);
output(0, 107) <= input(30);
output(0, 108) <= input(31);
output(0, 109) <= input(32);
output(0, 110) <= input(33);
output(0, 111) <= input(34);
output(0, 112) <= input(37);
output(0, 113) <= input(36);
output(0, 114) <= input(20);
output(0, 115) <= input(21);
output(0, 116) <= input(22);
output(0, 117) <= input(23);
output(0, 118) <= input(24);
output(0, 119) <= input(25);
output(0, 120) <= input(26);
output(0, 121) <= input(27);
output(0, 122) <= input(28);
output(0, 123) <= input(29);
output(0, 124) <= input(30);
output(0, 125) <= input(31);
output(0, 126) <= input(32);
output(0, 127) <= input(33);
output(0, 128) <= input(38);
output(0, 129) <= input(37);
output(0, 130) <= input(36);
output(0, 131) <= input(20);
output(0, 132) <= input(21);
output(0, 133) <= input(22);
output(0, 134) <= input(23);
output(0, 135) <= input(24);
output(0, 136) <= input(25);
output(0, 137) <= input(26);
output(0, 138) <= input(27);
output(0, 139) <= input(28);
output(0, 140) <= input(29);
output(0, 141) <= input(30);
output(0, 142) <= input(31);
output(0, 143) <= input(32);
output(0, 144) <= input(39);
output(0, 145) <= input(38);
output(0, 146) <= input(37);
output(0, 147) <= input(36);
output(0, 148) <= input(20);
output(0, 149) <= input(21);
output(0, 150) <= input(22);
output(0, 151) <= input(23);
output(0, 152) <= input(24);
output(0, 153) <= input(25);
output(0, 154) <= input(26);
output(0, 155) <= input(27);
output(0, 156) <= input(28);
output(0, 157) <= input(29);
output(0, 158) <= input(30);
output(0, 159) <= input(31);
output(0, 160) <= input(40);
output(0, 161) <= input(41);
output(0, 162) <= input(42);
output(0, 163) <= input(43);
output(0, 164) <= input(44);
output(0, 165) <= input(19);
output(0, 166) <= input(18);
output(0, 167) <= input(17);
output(0, 168) <= input(16);
output(0, 169) <= input(0);
output(0, 170) <= input(1);
output(0, 171) <= input(2);
output(0, 172) <= input(3);
output(0, 173) <= input(4);
output(0, 174) <= input(5);
output(0, 175) <= input(6);
output(0, 176) <= input(45);
output(0, 177) <= input(40);
output(0, 178) <= input(41);
output(0, 179) <= input(42);
output(0, 180) <= input(43);
output(0, 181) <= input(44);
output(0, 182) <= input(19);
output(0, 183) <= input(18);
output(0, 184) <= input(17);
output(0, 185) <= input(16);
output(0, 186) <= input(0);
output(0, 187) <= input(1);
output(0, 188) <= input(2);
output(0, 189) <= input(3);
output(0, 190) <= input(4);
output(0, 191) <= input(5);
output(0, 192) <= input(46);
output(0, 193) <= input(45);
output(0, 194) <= input(40);
output(0, 195) <= input(41);
output(0, 196) <= input(42);
output(0, 197) <= input(43);
output(0, 198) <= input(44);
output(0, 199) <= input(19);
output(0, 200) <= input(18);
output(0, 201) <= input(17);
output(0, 202) <= input(16);
output(0, 203) <= input(0);
output(0, 204) <= input(1);
output(0, 205) <= input(2);
output(0, 206) <= input(3);
output(0, 207) <= input(4);
output(0, 208) <= input(47);
output(0, 209) <= input(46);
output(0, 210) <= input(45);
output(0, 211) <= input(40);
output(0, 212) <= input(41);
output(0, 213) <= input(42);
output(0, 214) <= input(43);
output(0, 215) <= input(44);
output(0, 216) <= input(19);
output(0, 217) <= input(18);
output(0, 218) <= input(17);
output(0, 219) <= input(16);
output(0, 220) <= input(0);
output(0, 221) <= input(1);
output(0, 222) <= input(2);
output(0, 223) <= input(3);
output(0, 224) <= input(48);
output(0, 225) <= input(47);
output(0, 226) <= input(46);
output(0, 227) <= input(45);
output(0, 228) <= input(40);
output(0, 229) <= input(41);
output(0, 230) <= input(42);
output(0, 231) <= input(43);
output(0, 232) <= input(44);
output(0, 233) <= input(19);
output(0, 234) <= input(18);
output(0, 235) <= input(17);
output(0, 236) <= input(16);
output(0, 237) <= input(0);
output(0, 238) <= input(1);
output(0, 239) <= input(2);
output(0, 240) <= input(49);
output(0, 241) <= input(50);
output(0, 242) <= input(51);
output(0, 243) <= input(52);
output(0, 244) <= input(53);
output(0, 245) <= input(39);
output(0, 246) <= input(38);
output(0, 247) <= input(37);
output(0, 248) <= input(36);
output(0, 249) <= input(20);
output(0, 250) <= input(21);
output(0, 251) <= input(22);
output(0, 252) <= input(23);
output(0, 253) <= input(24);
output(0, 254) <= input(25);
output(0, 255) <= input(26);
when "1001" =>
output(0, 0) <= input(0);
output(0, 1) <= input(1);
output(0, 2) <= input(2);
output(0, 3) <= input(3);
output(0, 4) <= input(4);
output(0, 5) <= input(5);
output(0, 6) <= input(6);
output(0, 7) <= input(7);
output(0, 8) <= input(8);
output(0, 9) <= input(9);
output(0, 10) <= input(10);
output(0, 11) <= input(11);
output(0, 12) <= input(12);
output(0, 13) <= input(13);
output(0, 14) <= input(14);
output(0, 15) <= input(15);
output(0, 16) <= input(16);
output(0, 17) <= input(0);
output(0, 18) <= input(1);
output(0, 19) <= input(2);
output(0, 20) <= input(3);
output(0, 21) <= input(4);
output(0, 22) <= input(5);
output(0, 23) <= input(6);
output(0, 24) <= input(7);
output(0, 25) <= input(8);
output(0, 26) <= input(9);
output(0, 27) <= input(10);
output(0, 28) <= input(11);
output(0, 29) <= input(12);
output(0, 30) <= input(13);
output(0, 31) <= input(14);
output(0, 32) <= input(17);
output(0, 33) <= input(18);
output(0, 34) <= input(19);
output(0, 35) <= input(20);
output(0, 36) <= input(21);
output(0, 37) <= input(22);
output(0, 38) <= input(23);
output(0, 39) <= input(24);
output(0, 40) <= input(25);
output(0, 41) <= input(26);
output(0, 42) <= input(27);
output(0, 43) <= input(28);
output(0, 44) <= input(29);
output(0, 45) <= input(30);
output(0, 46) <= input(31);
output(0, 47) <= input(32);
output(0, 48) <= input(33);
output(0, 49) <= input(17);
output(0, 50) <= input(18);
output(0, 51) <= input(19);
output(0, 52) <= input(20);
output(0, 53) <= input(21);
output(0, 54) <= input(22);
output(0, 55) <= input(23);
output(0, 56) <= input(24);
output(0, 57) <= input(25);
output(0, 58) <= input(26);
output(0, 59) <= input(27);
output(0, 60) <= input(28);
output(0, 61) <= input(29);
output(0, 62) <= input(30);
output(0, 63) <= input(31);
output(0, 64) <= input(34);
output(0, 65) <= input(33);
output(0, 66) <= input(17);
output(0, 67) <= input(18);
output(0, 68) <= input(19);
output(0, 69) <= input(20);
output(0, 70) <= input(21);
output(0, 71) <= input(22);
output(0, 72) <= input(23);
output(0, 73) <= input(24);
output(0, 74) <= input(25);
output(0, 75) <= input(26);
output(0, 76) <= input(27);
output(0, 77) <= input(28);
output(0, 78) <= input(29);
output(0, 79) <= input(30);
output(0, 80) <= input(35);
output(0, 81) <= input(36);
output(0, 82) <= input(37);
output(0, 83) <= input(16);
output(0, 84) <= input(0);
output(0, 85) <= input(1);
output(0, 86) <= input(2);
output(0, 87) <= input(3);
output(0, 88) <= input(4);
output(0, 89) <= input(5);
output(0, 90) <= input(6);
output(0, 91) <= input(7);
output(0, 92) <= input(8);
output(0, 93) <= input(9);
output(0, 94) <= input(10);
output(0, 95) <= input(11);
output(0, 96) <= input(38);
output(0, 97) <= input(35);
output(0, 98) <= input(36);
output(0, 99) <= input(37);
output(0, 100) <= input(16);
output(0, 101) <= input(0);
output(0, 102) <= input(1);
output(0, 103) <= input(2);
output(0, 104) <= input(3);
output(0, 105) <= input(4);
output(0, 106) <= input(5);
output(0, 107) <= input(6);
output(0, 108) <= input(7);
output(0, 109) <= input(8);
output(0, 110) <= input(9);
output(0, 111) <= input(10);
output(0, 112) <= input(39);
output(0, 113) <= input(40);
output(0, 114) <= input(34);
output(0, 115) <= input(33);
output(0, 116) <= input(17);
output(0, 117) <= input(18);
output(0, 118) <= input(19);
output(0, 119) <= input(20);
output(0, 120) <= input(21);
output(0, 121) <= input(22);
output(0, 122) <= input(23);
output(0, 123) <= input(24);
output(0, 124) <= input(25);
output(0, 125) <= input(26);
output(0, 126) <= input(27);
output(0, 127) <= input(28);
output(0, 128) <= input(41);
output(0, 129) <= input(39);
output(0, 130) <= input(40);
output(0, 131) <= input(34);
output(0, 132) <= input(33);
output(0, 133) <= input(17);
output(0, 134) <= input(18);
output(0, 135) <= input(19);
output(0, 136) <= input(20);
output(0, 137) <= input(21);
output(0, 138) <= input(22);
output(0, 139) <= input(23);
output(0, 140) <= input(24);
output(0, 141) <= input(25);
output(0, 142) <= input(26);
output(0, 143) <= input(27);
output(0, 144) <= input(42);
output(0, 145) <= input(41);
output(0, 146) <= input(39);
output(0, 147) <= input(40);
output(0, 148) <= input(34);
output(0, 149) <= input(33);
output(0, 150) <= input(17);
output(0, 151) <= input(18);
output(0, 152) <= input(19);
output(0, 153) <= input(20);
output(0, 154) <= input(21);
output(0, 155) <= input(22);
output(0, 156) <= input(23);
output(0, 157) <= input(24);
output(0, 158) <= input(25);
output(0, 159) <= input(26);
output(0, 160) <= input(43);
output(0, 161) <= input(44);
output(0, 162) <= input(45);
output(0, 163) <= input(38);
output(0, 164) <= input(35);
output(0, 165) <= input(36);
output(0, 166) <= input(37);
output(0, 167) <= input(16);
output(0, 168) <= input(0);
output(0, 169) <= input(1);
output(0, 170) <= input(2);
output(0, 171) <= input(3);
output(0, 172) <= input(4);
output(0, 173) <= input(5);
output(0, 174) <= input(6);
output(0, 175) <= input(7);
output(0, 176) <= input(46);
output(0, 177) <= input(43);
output(0, 178) <= input(44);
output(0, 179) <= input(45);
output(0, 180) <= input(38);
output(0, 181) <= input(35);
output(0, 182) <= input(36);
output(0, 183) <= input(37);
output(0, 184) <= input(16);
output(0, 185) <= input(0);
output(0, 186) <= input(1);
output(0, 187) <= input(2);
output(0, 188) <= input(3);
output(0, 189) <= input(4);
output(0, 190) <= input(5);
output(0, 191) <= input(6);
output(0, 192) <= input(47);
output(0, 193) <= input(46);
output(0, 194) <= input(43);
output(0, 195) <= input(44);
output(0, 196) <= input(45);
output(0, 197) <= input(38);
output(0, 198) <= input(35);
output(0, 199) <= input(36);
output(0, 200) <= input(37);
output(0, 201) <= input(16);
output(0, 202) <= input(0);
output(0, 203) <= input(1);
output(0, 204) <= input(2);
output(0, 205) <= input(3);
output(0, 206) <= input(4);
output(0, 207) <= input(5);
output(0, 208) <= input(48);
output(0, 209) <= input(49);
output(0, 210) <= input(50);
output(0, 211) <= input(42);
output(0, 212) <= input(41);
output(0, 213) <= input(39);
output(0, 214) <= input(40);
output(0, 215) <= input(34);
output(0, 216) <= input(33);
output(0, 217) <= input(17);
output(0, 218) <= input(18);
output(0, 219) <= input(19);
output(0, 220) <= input(20);
output(0, 221) <= input(21);
output(0, 222) <= input(22);
output(0, 223) <= input(23);
output(0, 224) <= input(51);
output(0, 225) <= input(48);
output(0, 226) <= input(49);
output(0, 227) <= input(50);
output(0, 228) <= input(42);
output(0, 229) <= input(41);
output(0, 230) <= input(39);
output(0, 231) <= input(40);
output(0, 232) <= input(34);
output(0, 233) <= input(33);
output(0, 234) <= input(17);
output(0, 235) <= input(18);
output(0, 236) <= input(19);
output(0, 237) <= input(20);
output(0, 238) <= input(21);
output(0, 239) <= input(22);
output(0, 240) <= input(52);
output(0, 241) <= input(53);
output(0, 242) <= input(47);
output(0, 243) <= input(46);
output(0, 244) <= input(43);
output(0, 245) <= input(44);
output(0, 246) <= input(45);
output(0, 247) <= input(38);
output(0, 248) <= input(35);
output(0, 249) <= input(36);
output(0, 250) <= input(37);
output(0, 251) <= input(16);
output(0, 252) <= input(0);
output(0, 253) <= input(1);
output(0, 254) <= input(2);
output(0, 255) <= input(3);
output(1, 0) <= input(0);
output(1, 1) <= input(1);
output(1, 2) <= input(2);
output(1, 3) <= input(3);
output(1, 4) <= input(4);
output(1, 5) <= input(5);
output(1, 6) <= input(6);
output(1, 7) <= input(7);
output(1, 8) <= input(8);
output(1, 9) <= input(9);
output(1, 10) <= input(10);
output(1, 11) <= input(11);
output(1, 12) <= input(12);
output(1, 13) <= input(13);
output(1, 14) <= input(14);
output(1, 15) <= input(15);
output(1, 16) <= input(18);
output(1, 17) <= input(19);
output(1, 18) <= input(20);
output(1, 19) <= input(21);
output(1, 20) <= input(22);
output(1, 21) <= input(23);
output(1, 22) <= input(24);
output(1, 23) <= input(25);
output(1, 24) <= input(26);
output(1, 25) <= input(27);
output(1, 26) <= input(28);
output(1, 27) <= input(29);
output(1, 28) <= input(30);
output(1, 29) <= input(31);
output(1, 30) <= input(32);
output(1, 31) <= input(54);
output(1, 32) <= input(17);
output(1, 33) <= input(18);
output(1, 34) <= input(19);
output(1, 35) <= input(20);
output(1, 36) <= input(21);
output(1, 37) <= input(22);
output(1, 38) <= input(23);
output(1, 39) <= input(24);
output(1, 40) <= input(25);
output(1, 41) <= input(26);
output(1, 42) <= input(27);
output(1, 43) <= input(28);
output(1, 44) <= input(29);
output(1, 45) <= input(30);
output(1, 46) <= input(31);
output(1, 47) <= input(32);
output(1, 48) <= input(37);
output(1, 49) <= input(16);
output(1, 50) <= input(0);
output(1, 51) <= input(1);
output(1, 52) <= input(2);
output(1, 53) <= input(3);
output(1, 54) <= input(4);
output(1, 55) <= input(5);
output(1, 56) <= input(6);
output(1, 57) <= input(7);
output(1, 58) <= input(8);
output(1, 59) <= input(9);
output(1, 60) <= input(10);
output(1, 61) <= input(11);
output(1, 62) <= input(12);
output(1, 63) <= input(13);
output(1, 64) <= input(36);
output(1, 65) <= input(37);
output(1, 66) <= input(16);
output(1, 67) <= input(0);
output(1, 68) <= input(1);
output(1, 69) <= input(2);
output(1, 70) <= input(3);
output(1, 71) <= input(4);
output(1, 72) <= input(5);
output(1, 73) <= input(6);
output(1, 74) <= input(7);
output(1, 75) <= input(8);
output(1, 76) <= input(9);
output(1, 77) <= input(10);
output(1, 78) <= input(11);
output(1, 79) <= input(12);
output(1, 80) <= input(34);
output(1, 81) <= input(33);
output(1, 82) <= input(17);
output(1, 83) <= input(18);
output(1, 84) <= input(19);
output(1, 85) <= input(20);
output(1, 86) <= input(21);
output(1, 87) <= input(22);
output(1, 88) <= input(23);
output(1, 89) <= input(24);
output(1, 90) <= input(25);
output(1, 91) <= input(26);
output(1, 92) <= input(27);
output(1, 93) <= input(28);
output(1, 94) <= input(29);
output(1, 95) <= input(30);
output(1, 96) <= input(40);
output(1, 97) <= input(34);
output(1, 98) <= input(33);
output(1, 99) <= input(17);
output(1, 100) <= input(18);
output(1, 101) <= input(19);
output(1, 102) <= input(20);
output(1, 103) <= input(21);
output(1, 104) <= input(22);
output(1, 105) <= input(23);
output(1, 106) <= input(24);
output(1, 107) <= input(25);
output(1, 108) <= input(26);
output(1, 109) <= input(27);
output(1, 110) <= input(28);
output(1, 111) <= input(29);
output(1, 112) <= input(38);
output(1, 113) <= input(35);
output(1, 114) <= input(36);
output(1, 115) <= input(37);
output(1, 116) <= input(16);
output(1, 117) <= input(0);
output(1, 118) <= input(1);
output(1, 119) <= input(2);
output(1, 120) <= input(3);
output(1, 121) <= input(4);
output(1, 122) <= input(5);
output(1, 123) <= input(6);
output(1, 124) <= input(7);
output(1, 125) <= input(8);
output(1, 126) <= input(9);
output(1, 127) <= input(10);
output(1, 128) <= input(39);
output(1, 129) <= input(40);
output(1, 130) <= input(34);
output(1, 131) <= input(33);
output(1, 132) <= input(17);
output(1, 133) <= input(18);
output(1, 134) <= input(19);
output(1, 135) <= input(20);
output(1, 136) <= input(21);
output(1, 137) <= input(22);
output(1, 138) <= input(23);
output(1, 139) <= input(24);
output(1, 140) <= input(25);
output(1, 141) <= input(26);
output(1, 142) <= input(27);
output(1, 143) <= input(28);
output(1, 144) <= input(41);
output(1, 145) <= input(39);
output(1, 146) <= input(40);
output(1, 147) <= input(34);
output(1, 148) <= input(33);
output(1, 149) <= input(17);
output(1, 150) <= input(18);
output(1, 151) <= input(19);
output(1, 152) <= input(20);
output(1, 153) <= input(21);
output(1, 154) <= input(22);
output(1, 155) <= input(23);
output(1, 156) <= input(24);
output(1, 157) <= input(25);
output(1, 158) <= input(26);
output(1, 159) <= input(27);
output(1, 160) <= input(44);
output(1, 161) <= input(45);
output(1, 162) <= input(38);
output(1, 163) <= input(35);
output(1, 164) <= input(36);
output(1, 165) <= input(37);
output(1, 166) <= input(16);
output(1, 167) <= input(0);
output(1, 168) <= input(1);
output(1, 169) <= input(2);
output(1, 170) <= input(3);
output(1, 171) <= input(4);
output(1, 172) <= input(5);
output(1, 173) <= input(6);
output(1, 174) <= input(7);
output(1, 175) <= input(8);
output(1, 176) <= input(43);
output(1, 177) <= input(44);
output(1, 178) <= input(45);
output(1, 179) <= input(38);
output(1, 180) <= input(35);
output(1, 181) <= input(36);
output(1, 182) <= input(37);
output(1, 183) <= input(16);
output(1, 184) <= input(0);
output(1, 185) <= input(1);
output(1, 186) <= input(2);
output(1, 187) <= input(3);
output(1, 188) <= input(4);
output(1, 189) <= input(5);
output(1, 190) <= input(6);
output(1, 191) <= input(7);
output(1, 192) <= input(50);
output(1, 193) <= input(42);
output(1, 194) <= input(41);
output(1, 195) <= input(39);
output(1, 196) <= input(40);
output(1, 197) <= input(34);
output(1, 198) <= input(33);
output(1, 199) <= input(17);
output(1, 200) <= input(18);
output(1, 201) <= input(19);
output(1, 202) <= input(20);
output(1, 203) <= input(21);
output(1, 204) <= input(22);
output(1, 205) <= input(23);
output(1, 206) <= input(24);
output(1, 207) <= input(25);
output(1, 208) <= input(49);
output(1, 209) <= input(50);
output(1, 210) <= input(42);
output(1, 211) <= input(41);
output(1, 212) <= input(39);
output(1, 213) <= input(40);
output(1, 214) <= input(34);
output(1, 215) <= input(33);
output(1, 216) <= input(17);
output(1, 217) <= input(18);
output(1, 218) <= input(19);
output(1, 219) <= input(20);
output(1, 220) <= input(21);
output(1, 221) <= input(22);
output(1, 222) <= input(23);
output(1, 223) <= input(24);
output(1, 224) <= input(47);
output(1, 225) <= input(46);
output(1, 226) <= input(43);
output(1, 227) <= input(44);
output(1, 228) <= input(45);
output(1, 229) <= input(38);
output(1, 230) <= input(35);
output(1, 231) <= input(36);
output(1, 232) <= input(37);
output(1, 233) <= input(16);
output(1, 234) <= input(0);
output(1, 235) <= input(1);
output(1, 236) <= input(2);
output(1, 237) <= input(3);
output(1, 238) <= input(4);
output(1, 239) <= input(5);
output(1, 240) <= input(48);
output(1, 241) <= input(49);
output(1, 242) <= input(50);
output(1, 243) <= input(42);
output(1, 244) <= input(41);
output(1, 245) <= input(39);
output(1, 246) <= input(40);
output(1, 247) <= input(34);
output(1, 248) <= input(33);
output(1, 249) <= input(17);
output(1, 250) <= input(18);
output(1, 251) <= input(19);
output(1, 252) <= input(20);
output(1, 253) <= input(21);
output(1, 254) <= input(22);
output(1, 255) <= input(23);
output(2, 0) <= input(0);
output(2, 1) <= input(1);
output(2, 2) <= input(2);
output(2, 3) <= input(3);
output(2, 4) <= input(4);
output(2, 5) <= input(5);
output(2, 6) <= input(6);
output(2, 7) <= input(7);
output(2, 8) <= input(8);
output(2, 9) <= input(9);
output(2, 10) <= input(10);
output(2, 11) <= input(11);
output(2, 12) <= input(12);
output(2, 13) <= input(13);
output(2, 14) <= input(14);
output(2, 15) <= input(15);
output(2, 16) <= input(18);
output(2, 17) <= input(19);
output(2, 18) <= input(20);
output(2, 19) <= input(21);
output(2, 20) <= input(22);
output(2, 21) <= input(23);
output(2, 22) <= input(24);
output(2, 23) <= input(25);
output(2, 24) <= input(26);
output(2, 25) <= input(27);
output(2, 26) <= input(28);
output(2, 27) <= input(29);
output(2, 28) <= input(30);
output(2, 29) <= input(31);
output(2, 30) <= input(32);
output(2, 31) <= input(54);
output(2, 32) <= input(16);
output(2, 33) <= input(0);
output(2, 34) <= input(1);
output(2, 35) <= input(2);
output(2, 36) <= input(3);
output(2, 37) <= input(4);
output(2, 38) <= input(5);
output(2, 39) <= input(6);
output(2, 40) <= input(7);
output(2, 41) <= input(8);
output(2, 42) <= input(9);
output(2, 43) <= input(10);
output(2, 44) <= input(11);
output(2, 45) <= input(12);
output(2, 46) <= input(13);
output(2, 47) <= input(14);
output(2, 48) <= input(17);
output(2, 49) <= input(18);
output(2, 50) <= input(19);
output(2, 51) <= input(20);
output(2, 52) <= input(21);
output(2, 53) <= input(22);
output(2, 54) <= input(23);
output(2, 55) <= input(24);
output(2, 56) <= input(25);
output(2, 57) <= input(26);
output(2, 58) <= input(27);
output(2, 59) <= input(28);
output(2, 60) <= input(29);
output(2, 61) <= input(30);
output(2, 62) <= input(31);
output(2, 63) <= input(32);
output(2, 64) <= input(33);
output(2, 65) <= input(17);
output(2, 66) <= input(18);
output(2, 67) <= input(19);
output(2, 68) <= input(20);
output(2, 69) <= input(21);
output(2, 70) <= input(22);
output(2, 71) <= input(23);
output(2, 72) <= input(24);
output(2, 73) <= input(25);
output(2, 74) <= input(26);
output(2, 75) <= input(27);
output(2, 76) <= input(28);
output(2, 77) <= input(29);
output(2, 78) <= input(30);
output(2, 79) <= input(31);
output(2, 80) <= input(36);
output(2, 81) <= input(37);
output(2, 82) <= input(16);
output(2, 83) <= input(0);
output(2, 84) <= input(1);
output(2, 85) <= input(2);
output(2, 86) <= input(3);
output(2, 87) <= input(4);
output(2, 88) <= input(5);
output(2, 89) <= input(6);
output(2, 90) <= input(7);
output(2, 91) <= input(8);
output(2, 92) <= input(9);
output(2, 93) <= input(10);
output(2, 94) <= input(11);
output(2, 95) <= input(12);
output(2, 96) <= input(34);
output(2, 97) <= input(33);
output(2, 98) <= input(17);
output(2, 99) <= input(18);
output(2, 100) <= input(19);
output(2, 101) <= input(20);
output(2, 102) <= input(21);
output(2, 103) <= input(22);
output(2, 104) <= input(23);
output(2, 105) <= input(24);
output(2, 106) <= input(25);
output(2, 107) <= input(26);
output(2, 108) <= input(27);
output(2, 109) <= input(28);
output(2, 110) <= input(29);
output(2, 111) <= input(30);
output(2, 112) <= input(35);
output(2, 113) <= input(36);
output(2, 114) <= input(37);
output(2, 115) <= input(16);
output(2, 116) <= input(0);
output(2, 117) <= input(1);
output(2, 118) <= input(2);
output(2, 119) <= input(3);
output(2, 120) <= input(4);
output(2, 121) <= input(5);
output(2, 122) <= input(6);
output(2, 123) <= input(7);
output(2, 124) <= input(8);
output(2, 125) <= input(9);
output(2, 126) <= input(10);
output(2, 127) <= input(11);
output(2, 128) <= input(38);
output(2, 129) <= input(35);
output(2, 130) <= input(36);
output(2, 131) <= input(37);
output(2, 132) <= input(16);
output(2, 133) <= input(0);
output(2, 134) <= input(1);
output(2, 135) <= input(2);
output(2, 136) <= input(3);
output(2, 137) <= input(4);
output(2, 138) <= input(5);
output(2, 139) <= input(6);
output(2, 140) <= input(7);
output(2, 141) <= input(8);
output(2, 142) <= input(9);
output(2, 143) <= input(10);
output(2, 144) <= input(39);
output(2, 145) <= input(40);
output(2, 146) <= input(34);
output(2, 147) <= input(33);
output(2, 148) <= input(17);
output(2, 149) <= input(18);
output(2, 150) <= input(19);
output(2, 151) <= input(20);
output(2, 152) <= input(21);
output(2, 153) <= input(22);
output(2, 154) <= input(23);
output(2, 155) <= input(24);
output(2, 156) <= input(25);
output(2, 157) <= input(26);
output(2, 158) <= input(27);
output(2, 159) <= input(28);
output(2, 160) <= input(45);
output(2, 161) <= input(38);
output(2, 162) <= input(35);
output(2, 163) <= input(36);
output(2, 164) <= input(37);
output(2, 165) <= input(16);
output(2, 166) <= input(0);
output(2, 167) <= input(1);
output(2, 168) <= input(2);
output(2, 169) <= input(3);
output(2, 170) <= input(4);
output(2, 171) <= input(5);
output(2, 172) <= input(6);
output(2, 173) <= input(7);
output(2, 174) <= input(8);
output(2, 175) <= input(9);
output(2, 176) <= input(41);
output(2, 177) <= input(39);
output(2, 178) <= input(40);
output(2, 179) <= input(34);
output(2, 180) <= input(33);
output(2, 181) <= input(17);
output(2, 182) <= input(18);
output(2, 183) <= input(19);
output(2, 184) <= input(20);
output(2, 185) <= input(21);
output(2, 186) <= input(22);
output(2, 187) <= input(23);
output(2, 188) <= input(24);
output(2, 189) <= input(25);
output(2, 190) <= input(26);
output(2, 191) <= input(27);
output(2, 192) <= input(42);
output(2, 193) <= input(41);
output(2, 194) <= input(39);
output(2, 195) <= input(40);
output(2, 196) <= input(34);
output(2, 197) <= input(33);
output(2, 198) <= input(17);
output(2, 199) <= input(18);
output(2, 200) <= input(19);
output(2, 201) <= input(20);
output(2, 202) <= input(21);
output(2, 203) <= input(22);
output(2, 204) <= input(23);
output(2, 205) <= input(24);
output(2, 206) <= input(25);
output(2, 207) <= input(26);
output(2, 208) <= input(43);
output(2, 209) <= input(44);
output(2, 210) <= input(45);
output(2, 211) <= input(38);
output(2, 212) <= input(35);
output(2, 213) <= input(36);
output(2, 214) <= input(37);
output(2, 215) <= input(16);
output(2, 216) <= input(0);
output(2, 217) <= input(1);
output(2, 218) <= input(2);
output(2, 219) <= input(3);
output(2, 220) <= input(4);
output(2, 221) <= input(5);
output(2, 222) <= input(6);
output(2, 223) <= input(7);
output(2, 224) <= input(50);
output(2, 225) <= input(42);
output(2, 226) <= input(41);
output(2, 227) <= input(39);
output(2, 228) <= input(40);
output(2, 229) <= input(34);
output(2, 230) <= input(33);
output(2, 231) <= input(17);
output(2, 232) <= input(18);
output(2, 233) <= input(19);
output(2, 234) <= input(20);
output(2, 235) <= input(21);
output(2, 236) <= input(22);
output(2, 237) <= input(23);
output(2, 238) <= input(24);
output(2, 239) <= input(25);
output(2, 240) <= input(46);
output(2, 241) <= input(43);
output(2, 242) <= input(44);
output(2, 243) <= input(45);
output(2, 244) <= input(38);
output(2, 245) <= input(35);
output(2, 246) <= input(36);
output(2, 247) <= input(37);
output(2, 248) <= input(16);
output(2, 249) <= input(0);
output(2, 250) <= input(1);
output(2, 251) <= input(2);
output(2, 252) <= input(3);
output(2, 253) <= input(4);
output(2, 254) <= input(5);
output(2, 255) <= input(6);
when "1010" =>
output(0, 0) <= input(0);
output(0, 1) <= input(1);
output(0, 2) <= input(2);
output(0, 3) <= input(3);
output(0, 4) <= input(4);
output(0, 5) <= input(5);
output(0, 6) <= input(6);
output(0, 7) <= input(7);
output(0, 8) <= input(8);
output(0, 9) <= input(9);
output(0, 10) <= input(10);
output(0, 11) <= input(11);
output(0, 12) <= input(12);
output(0, 13) <= input(13);
output(0, 14) <= input(14);
output(0, 15) <= input(15);
output(0, 16) <= input(16);
output(0, 17) <= input(17);
output(0, 18) <= input(18);
output(0, 19) <= input(19);
output(0, 20) <= input(20);
output(0, 21) <= input(21);
output(0, 22) <= input(22);
output(0, 23) <= input(23);
output(0, 24) <= input(24);
output(0, 25) <= input(25);
output(0, 26) <= input(26);
output(0, 27) <= input(27);
output(0, 28) <= input(28);
output(0, 29) <= input(29);
output(0, 30) <= input(30);
output(0, 31) <= input(31);
output(0, 32) <= input(32);
output(0, 33) <= input(0);
output(0, 34) <= input(1);
output(0, 35) <= input(2);
output(0, 36) <= input(3);
output(0, 37) <= input(4);
output(0, 38) <= input(5);
output(0, 39) <= input(6);
output(0, 40) <= input(7);
output(0, 41) <= input(8);
output(0, 42) <= input(9);
output(0, 43) <= input(10);
output(0, 44) <= input(11);
output(0, 45) <= input(12);
output(0, 46) <= input(13);
output(0, 47) <= input(14);
output(0, 48) <= input(33);
output(0, 49) <= input(16);
output(0, 50) <= input(17);
output(0, 51) <= input(18);
output(0, 52) <= input(19);
output(0, 53) <= input(20);
output(0, 54) <= input(21);
output(0, 55) <= input(22);
output(0, 56) <= input(23);
output(0, 57) <= input(24);
output(0, 58) <= input(25);
output(0, 59) <= input(26);
output(0, 60) <= input(27);
output(0, 61) <= input(28);
output(0, 62) <= input(29);
output(0, 63) <= input(30);
output(0, 64) <= input(34);
output(0, 65) <= input(32);
output(0, 66) <= input(0);
output(0, 67) <= input(1);
output(0, 68) <= input(2);
output(0, 69) <= input(3);
output(0, 70) <= input(4);
output(0, 71) <= input(5);
output(0, 72) <= input(6);
output(0, 73) <= input(7);
output(0, 74) <= input(8);
output(0, 75) <= input(9);
output(0, 76) <= input(10);
output(0, 77) <= input(11);
output(0, 78) <= input(12);
output(0, 79) <= input(13);
output(0, 80) <= input(35);
output(0, 81) <= input(33);
output(0, 82) <= input(16);
output(0, 83) <= input(17);
output(0, 84) <= input(18);
output(0, 85) <= input(19);
output(0, 86) <= input(20);
output(0, 87) <= input(21);
output(0, 88) <= input(22);
output(0, 89) <= input(23);
output(0, 90) <= input(24);
output(0, 91) <= input(25);
output(0, 92) <= input(26);
output(0, 93) <= input(27);
output(0, 94) <= input(28);
output(0, 95) <= input(29);
output(0, 96) <= input(36);
output(0, 97) <= input(34);
output(0, 98) <= input(32);
output(0, 99) <= input(0);
output(0, 100) <= input(1);
output(0, 101) <= input(2);
output(0, 102) <= input(3);
output(0, 103) <= input(4);
output(0, 104) <= input(5);
output(0, 105) <= input(6);
output(0, 106) <= input(7);
output(0, 107) <= input(8);
output(0, 108) <= input(9);
output(0, 109) <= input(10);
output(0, 110) <= input(11);
output(0, 111) <= input(12);
output(0, 112) <= input(37);
output(0, 113) <= input(35);
output(0, 114) <= input(33);
output(0, 115) <= input(16);
output(0, 116) <= input(17);
output(0, 117) <= input(18);
output(0, 118) <= input(19);
output(0, 119) <= input(20);
output(0, 120) <= input(21);
output(0, 121) <= input(22);
output(0, 122) <= input(23);
output(0, 123) <= input(24);
output(0, 124) <= input(25);
output(0, 125) <= input(26);
output(0, 126) <= input(27);
output(0, 127) <= input(28);
output(0, 128) <= input(38);
output(0, 129) <= input(37);
output(0, 130) <= input(35);
output(0, 131) <= input(33);
output(0, 132) <= input(16);
output(0, 133) <= input(17);
output(0, 134) <= input(18);
output(0, 135) <= input(19);
output(0, 136) <= input(20);
output(0, 137) <= input(21);
output(0, 138) <= input(22);
output(0, 139) <= input(23);
output(0, 140) <= input(24);
output(0, 141) <= input(25);
output(0, 142) <= input(26);
output(0, 143) <= input(27);
output(0, 144) <= input(39);
output(0, 145) <= input(40);
output(0, 146) <= input(36);
output(0, 147) <= input(34);
output(0, 148) <= input(32);
output(0, 149) <= input(0);
output(0, 150) <= input(1);
output(0, 151) <= input(2);
output(0, 152) <= input(3);
output(0, 153) <= input(4);
output(0, 154) <= input(5);
output(0, 155) <= input(6);
output(0, 156) <= input(7);
output(0, 157) <= input(8);
output(0, 158) <= input(9);
output(0, 159) <= input(10);
output(0, 160) <= input(41);
output(0, 161) <= input(38);
output(0, 162) <= input(37);
output(0, 163) <= input(35);
output(0, 164) <= input(33);
output(0, 165) <= input(16);
output(0, 166) <= input(17);
output(0, 167) <= input(18);
output(0, 168) <= input(19);
output(0, 169) <= input(20);
output(0, 170) <= input(21);
output(0, 171) <= input(22);
output(0, 172) <= input(23);
output(0, 173) <= input(24);
output(0, 174) <= input(25);
output(0, 175) <= input(26);
output(0, 176) <= input(42);
output(0, 177) <= input(39);
output(0, 178) <= input(40);
output(0, 179) <= input(36);
output(0, 180) <= input(34);
output(0, 181) <= input(32);
output(0, 182) <= input(0);
output(0, 183) <= input(1);
output(0, 184) <= input(2);
output(0, 185) <= input(3);
output(0, 186) <= input(4);
output(0, 187) <= input(5);
output(0, 188) <= input(6);
output(0, 189) <= input(7);
output(0, 190) <= input(8);
output(0, 191) <= input(9);
output(0, 192) <= input(43);
output(0, 193) <= input(41);
output(0, 194) <= input(38);
output(0, 195) <= input(37);
output(0, 196) <= input(35);
output(0, 197) <= input(33);
output(0, 198) <= input(16);
output(0, 199) <= input(17);
output(0, 200) <= input(18);
output(0, 201) <= input(19);
output(0, 202) <= input(20);
output(0, 203) <= input(21);
output(0, 204) <= input(22);
output(0, 205) <= input(23);
output(0, 206) <= input(24);
output(0, 207) <= input(25);
output(0, 208) <= input(44);
output(0, 209) <= input(42);
output(0, 210) <= input(39);
output(0, 211) <= input(40);
output(0, 212) <= input(36);
output(0, 213) <= input(34);
output(0, 214) <= input(32);
output(0, 215) <= input(0);
output(0, 216) <= input(1);
output(0, 217) <= input(2);
output(0, 218) <= input(3);
output(0, 219) <= input(4);
output(0, 220) <= input(5);
output(0, 221) <= input(6);
output(0, 222) <= input(7);
output(0, 223) <= input(8);
output(0, 224) <= input(45);
output(0, 225) <= input(43);
output(0, 226) <= input(41);
output(0, 227) <= input(38);
output(0, 228) <= input(37);
output(0, 229) <= input(35);
output(0, 230) <= input(33);
output(0, 231) <= input(16);
output(0, 232) <= input(17);
output(0, 233) <= input(18);
output(0, 234) <= input(19);
output(0, 235) <= input(20);
output(0, 236) <= input(21);
output(0, 237) <= input(22);
output(0, 238) <= input(23);
output(0, 239) <= input(24);
output(0, 240) <= input(46);
output(0, 241) <= input(44);
output(0, 242) <= input(42);
output(0, 243) <= input(39);
output(0, 244) <= input(40);
output(0, 245) <= input(36);
output(0, 246) <= input(34);
output(0, 247) <= input(32);
output(0, 248) <= input(0);
output(0, 249) <= input(1);
output(0, 250) <= input(2);
output(0, 251) <= input(3);
output(0, 252) <= input(4);
output(0, 253) <= input(5);
output(0, 254) <= input(6);
output(0, 255) <= input(7);
output(1, 0) <= input(17);
output(1, 1) <= input(18);
output(1, 2) <= input(19);
output(1, 3) <= input(20);
output(1, 4) <= input(21);
output(1, 5) <= input(22);
output(1, 6) <= input(23);
output(1, 7) <= input(24);
output(1, 8) <= input(25);
output(1, 9) <= input(26);
output(1, 10) <= input(27);
output(1, 11) <= input(28);
output(1, 12) <= input(29);
output(1, 13) <= input(30);
output(1, 14) <= input(31);
output(1, 15) <= input(47);
output(1, 16) <= input(0);
output(1, 17) <= input(1);
output(1, 18) <= input(2);
output(1, 19) <= input(3);
output(1, 20) <= input(4);
output(1, 21) <= input(5);
output(1, 22) <= input(6);
output(1, 23) <= input(7);
output(1, 24) <= input(8);
output(1, 25) <= input(9);
output(1, 26) <= input(10);
output(1, 27) <= input(11);
output(1, 28) <= input(12);
output(1, 29) <= input(13);
output(1, 30) <= input(14);
output(1, 31) <= input(15);
output(1, 32) <= input(16);
output(1, 33) <= input(17);
output(1, 34) <= input(18);
output(1, 35) <= input(19);
output(1, 36) <= input(20);
output(1, 37) <= input(21);
output(1, 38) <= input(22);
output(1, 39) <= input(23);
output(1, 40) <= input(24);
output(1, 41) <= input(25);
output(1, 42) <= input(26);
output(1, 43) <= input(27);
output(1, 44) <= input(28);
output(1, 45) <= input(29);
output(1, 46) <= input(30);
output(1, 47) <= input(31);
output(1, 48) <= input(32);
output(1, 49) <= input(0);
output(1, 50) <= input(1);
output(1, 51) <= input(2);
output(1, 52) <= input(3);
output(1, 53) <= input(4);
output(1, 54) <= input(5);
output(1, 55) <= input(6);
output(1, 56) <= input(7);
output(1, 57) <= input(8);
output(1, 58) <= input(9);
output(1, 59) <= input(10);
output(1, 60) <= input(11);
output(1, 61) <= input(12);
output(1, 62) <= input(13);
output(1, 63) <= input(14);
output(1, 64) <= input(33);
output(1, 65) <= input(16);
output(1, 66) <= input(17);
output(1, 67) <= input(18);
output(1, 68) <= input(19);
output(1, 69) <= input(20);
output(1, 70) <= input(21);
output(1, 71) <= input(22);
output(1, 72) <= input(23);
output(1, 73) <= input(24);
output(1, 74) <= input(25);
output(1, 75) <= input(26);
output(1, 76) <= input(27);
output(1, 77) <= input(28);
output(1, 78) <= input(29);
output(1, 79) <= input(30);
output(1, 80) <= input(34);
output(1, 81) <= input(32);
output(1, 82) <= input(0);
output(1, 83) <= input(1);
output(1, 84) <= input(2);
output(1, 85) <= input(3);
output(1, 86) <= input(4);
output(1, 87) <= input(5);
output(1, 88) <= input(6);
output(1, 89) <= input(7);
output(1, 90) <= input(8);
output(1, 91) <= input(9);
output(1, 92) <= input(10);
output(1, 93) <= input(11);
output(1, 94) <= input(12);
output(1, 95) <= input(13);
output(1, 96) <= input(35);
output(1, 97) <= input(33);
output(1, 98) <= input(16);
output(1, 99) <= input(17);
output(1, 100) <= input(18);
output(1, 101) <= input(19);
output(1, 102) <= input(20);
output(1, 103) <= input(21);
output(1, 104) <= input(22);
output(1, 105) <= input(23);
output(1, 106) <= input(24);
output(1, 107) <= input(25);
output(1, 108) <= input(26);
output(1, 109) <= input(27);
output(1, 110) <= input(28);
output(1, 111) <= input(29);
output(1, 112) <= input(36);
output(1, 113) <= input(34);
output(1, 114) <= input(32);
output(1, 115) <= input(0);
output(1, 116) <= input(1);
output(1, 117) <= input(2);
output(1, 118) <= input(3);
output(1, 119) <= input(4);
output(1, 120) <= input(5);
output(1, 121) <= input(6);
output(1, 122) <= input(7);
output(1, 123) <= input(8);
output(1, 124) <= input(9);
output(1, 125) <= input(10);
output(1, 126) <= input(11);
output(1, 127) <= input(12);
output(1, 128) <= input(37);
output(1, 129) <= input(35);
output(1, 130) <= input(33);
output(1, 131) <= input(16);
output(1, 132) <= input(17);
output(1, 133) <= input(18);
output(1, 134) <= input(19);
output(1, 135) <= input(20);
output(1, 136) <= input(21);
output(1, 137) <= input(22);
output(1, 138) <= input(23);
output(1, 139) <= input(24);
output(1, 140) <= input(25);
output(1, 141) <= input(26);
output(1, 142) <= input(27);
output(1, 143) <= input(28);
output(1, 144) <= input(40);
output(1, 145) <= input(36);
output(1, 146) <= input(34);
output(1, 147) <= input(32);
output(1, 148) <= input(0);
output(1, 149) <= input(1);
output(1, 150) <= input(2);
output(1, 151) <= input(3);
output(1, 152) <= input(4);
output(1, 153) <= input(5);
output(1, 154) <= input(6);
output(1, 155) <= input(7);
output(1, 156) <= input(8);
output(1, 157) <= input(9);
output(1, 158) <= input(10);
output(1, 159) <= input(11);
output(1, 160) <= input(38);
output(1, 161) <= input(37);
output(1, 162) <= input(35);
output(1, 163) <= input(33);
output(1, 164) <= input(16);
output(1, 165) <= input(17);
output(1, 166) <= input(18);
output(1, 167) <= input(19);
output(1, 168) <= input(20);
output(1, 169) <= input(21);
output(1, 170) <= input(22);
output(1, 171) <= input(23);
output(1, 172) <= input(24);
output(1, 173) <= input(25);
output(1, 174) <= input(26);
output(1, 175) <= input(27);
output(1, 176) <= input(39);
output(1, 177) <= input(40);
output(1, 178) <= input(36);
output(1, 179) <= input(34);
output(1, 180) <= input(32);
output(1, 181) <= input(0);
output(1, 182) <= input(1);
output(1, 183) <= input(2);
output(1, 184) <= input(3);
output(1, 185) <= input(4);
output(1, 186) <= input(5);
output(1, 187) <= input(6);
output(1, 188) <= input(7);
output(1, 189) <= input(8);
output(1, 190) <= input(9);
output(1, 191) <= input(10);
output(1, 192) <= input(41);
output(1, 193) <= input(38);
output(1, 194) <= input(37);
output(1, 195) <= input(35);
output(1, 196) <= input(33);
output(1, 197) <= input(16);
output(1, 198) <= input(17);
output(1, 199) <= input(18);
output(1, 200) <= input(19);
output(1, 201) <= input(20);
output(1, 202) <= input(21);
output(1, 203) <= input(22);
output(1, 204) <= input(23);
output(1, 205) <= input(24);
output(1, 206) <= input(25);
output(1, 207) <= input(26);
output(1, 208) <= input(42);
output(1, 209) <= input(39);
output(1, 210) <= input(40);
output(1, 211) <= input(36);
output(1, 212) <= input(34);
output(1, 213) <= input(32);
output(1, 214) <= input(0);
output(1, 215) <= input(1);
output(1, 216) <= input(2);
output(1, 217) <= input(3);
output(1, 218) <= input(4);
output(1, 219) <= input(5);
output(1, 220) <= input(6);
output(1, 221) <= input(7);
output(1, 222) <= input(8);
output(1, 223) <= input(9);
output(1, 224) <= input(43);
output(1, 225) <= input(41);
output(1, 226) <= input(38);
output(1, 227) <= input(37);
output(1, 228) <= input(35);
output(1, 229) <= input(33);
output(1, 230) <= input(16);
output(1, 231) <= input(17);
output(1, 232) <= input(18);
output(1, 233) <= input(19);
output(1, 234) <= input(20);
output(1, 235) <= input(21);
output(1, 236) <= input(22);
output(1, 237) <= input(23);
output(1, 238) <= input(24);
output(1, 239) <= input(25);
output(1, 240) <= input(44);
output(1, 241) <= input(42);
output(1, 242) <= input(39);
output(1, 243) <= input(40);
output(1, 244) <= input(36);
output(1, 245) <= input(34);
output(1, 246) <= input(32);
output(1, 247) <= input(0);
output(1, 248) <= input(1);
output(1, 249) <= input(2);
output(1, 250) <= input(3);
output(1, 251) <= input(4);
output(1, 252) <= input(5);
output(1, 253) <= input(6);
output(1, 254) <= input(7);
output(1, 255) <= input(8);
when "1011" =>
output(0, 0) <= input(0);
output(0, 1) <= input(1);
output(0, 2) <= input(2);
output(0, 3) <= input(3);
output(0, 4) <= input(4);
output(0, 5) <= input(5);
output(0, 6) <= input(6);
output(0, 7) <= input(7);
output(0, 8) <= input(8);
output(0, 9) <= input(9);
output(0, 10) <= input(10);
output(0, 11) <= input(11);
output(0, 12) <= input(12);
output(0, 13) <= input(13);
output(0, 14) <= input(14);
output(0, 15) <= input(15);
output(0, 16) <= input(16);
output(0, 17) <= input(17);
output(0, 18) <= input(18);
output(0, 19) <= input(19);
output(0, 20) <= input(20);
output(0, 21) <= input(21);
output(0, 22) <= input(22);
output(0, 23) <= input(23);
output(0, 24) <= input(24);
output(0, 25) <= input(25);
output(0, 26) <= input(26);
output(0, 27) <= input(27);
output(0, 28) <= input(28);
output(0, 29) <= input(29);
output(0, 30) <= input(30);
output(0, 31) <= input(31);
output(0, 32) <= input(32);
output(0, 33) <= input(0);
output(0, 34) <= input(1);
output(0, 35) <= input(2);
output(0, 36) <= input(3);
output(0, 37) <= input(4);
output(0, 38) <= input(5);
output(0, 39) <= input(6);
output(0, 40) <= input(7);
output(0, 41) <= input(8);
output(0, 42) <= input(9);
output(0, 43) <= input(10);
output(0, 44) <= input(11);
output(0, 45) <= input(12);
output(0, 46) <= input(13);
output(0, 47) <= input(14);
output(0, 48) <= input(33);
output(0, 49) <= input(16);
output(0, 50) <= input(17);
output(0, 51) <= input(18);
output(0, 52) <= input(19);
output(0, 53) <= input(20);
output(0, 54) <= input(21);
output(0, 55) <= input(22);
output(0, 56) <= input(23);
output(0, 57) <= input(24);
output(0, 58) <= input(25);
output(0, 59) <= input(26);
output(0, 60) <= input(27);
output(0, 61) <= input(28);
output(0, 62) <= input(29);
output(0, 63) <= input(30);
output(0, 64) <= input(34);
output(0, 65) <= input(32);
output(0, 66) <= input(0);
output(0, 67) <= input(1);
output(0, 68) <= input(2);
output(0, 69) <= input(3);
output(0, 70) <= input(4);
output(0, 71) <= input(5);
output(0, 72) <= input(6);
output(0, 73) <= input(7);
output(0, 74) <= input(8);
output(0, 75) <= input(9);
output(0, 76) <= input(10);
output(0, 77) <= input(11);
output(0, 78) <= input(12);
output(0, 79) <= input(13);
output(0, 80) <= input(35);
output(0, 81) <= input(33);
output(0, 82) <= input(16);
output(0, 83) <= input(17);
output(0, 84) <= input(18);
output(0, 85) <= input(19);
output(0, 86) <= input(20);
output(0, 87) <= input(21);
output(0, 88) <= input(22);
output(0, 89) <= input(23);
output(0, 90) <= input(24);
output(0, 91) <= input(25);
output(0, 92) <= input(26);
output(0, 93) <= input(27);
output(0, 94) <= input(28);
output(0, 95) <= input(29);
output(0, 96) <= input(36);
output(0, 97) <= input(34);
output(0, 98) <= input(32);
output(0, 99) <= input(0);
output(0, 100) <= input(1);
output(0, 101) <= input(2);
output(0, 102) <= input(3);
output(0, 103) <= input(4);
output(0, 104) <= input(5);
output(0, 105) <= input(6);
output(0, 106) <= input(7);
output(0, 107) <= input(8);
output(0, 108) <= input(9);
output(0, 109) <= input(10);
output(0, 110) <= input(11);
output(0, 111) <= input(12);
output(0, 112) <= input(36);
output(0, 113) <= input(34);
output(0, 114) <= input(32);
output(0, 115) <= input(0);
output(0, 116) <= input(1);
output(0, 117) <= input(2);
output(0, 118) <= input(3);
output(0, 119) <= input(4);
output(0, 120) <= input(5);
output(0, 121) <= input(6);
output(0, 122) <= input(7);
output(0, 123) <= input(8);
output(0, 124) <= input(9);
output(0, 125) <= input(10);
output(0, 126) <= input(11);
output(0, 127) <= input(12);
output(0, 128) <= input(37);
output(0, 129) <= input(35);
output(0, 130) <= input(33);
output(0, 131) <= input(16);
output(0, 132) <= input(17);
output(0, 133) <= input(18);
output(0, 134) <= input(19);
output(0, 135) <= input(20);
output(0, 136) <= input(21);
output(0, 137) <= input(22);
output(0, 138) <= input(23);
output(0, 139) <= input(24);
output(0, 140) <= input(25);
output(0, 141) <= input(26);
output(0, 142) <= input(27);
output(0, 143) <= input(28);
output(0, 144) <= input(38);
output(0, 145) <= input(36);
output(0, 146) <= input(34);
output(0, 147) <= input(32);
output(0, 148) <= input(0);
output(0, 149) <= input(1);
output(0, 150) <= input(2);
output(0, 151) <= input(3);
output(0, 152) <= input(4);
output(0, 153) <= input(5);
output(0, 154) <= input(6);
output(0, 155) <= input(7);
output(0, 156) <= input(8);
output(0, 157) <= input(9);
output(0, 158) <= input(10);
output(0, 159) <= input(11);
output(0, 160) <= input(39);
output(0, 161) <= input(37);
output(0, 162) <= input(35);
output(0, 163) <= input(33);
output(0, 164) <= input(16);
output(0, 165) <= input(17);
output(0, 166) <= input(18);
output(0, 167) <= input(19);
output(0, 168) <= input(20);
output(0, 169) <= input(21);
output(0, 170) <= input(22);
output(0, 171) <= input(23);
output(0, 172) <= input(24);
output(0, 173) <= input(25);
output(0, 174) <= input(26);
output(0, 175) <= input(27);
output(0, 176) <= input(40);
output(0, 177) <= input(38);
output(0, 178) <= input(36);
output(0, 179) <= input(34);
output(0, 180) <= input(32);
output(0, 181) <= input(0);
output(0, 182) <= input(1);
output(0, 183) <= input(2);
output(0, 184) <= input(3);
output(0, 185) <= input(4);
output(0, 186) <= input(5);
output(0, 187) <= input(6);
output(0, 188) <= input(7);
output(0, 189) <= input(8);
output(0, 190) <= input(9);
output(0, 191) <= input(10);
output(0, 192) <= input(41);
output(0, 193) <= input(39);
output(0, 194) <= input(37);
output(0, 195) <= input(35);
output(0, 196) <= input(33);
output(0, 197) <= input(16);
output(0, 198) <= input(17);
output(0, 199) <= input(18);
output(0, 200) <= input(19);
output(0, 201) <= input(20);
output(0, 202) <= input(21);
output(0, 203) <= input(22);
output(0, 204) <= input(23);
output(0, 205) <= input(24);
output(0, 206) <= input(25);
output(0, 207) <= input(26);
output(0, 208) <= input(42);
output(0, 209) <= input(40);
output(0, 210) <= input(38);
output(0, 211) <= input(36);
output(0, 212) <= input(34);
output(0, 213) <= input(32);
output(0, 214) <= input(0);
output(0, 215) <= input(1);
output(0, 216) <= input(2);
output(0, 217) <= input(3);
output(0, 218) <= input(4);
output(0, 219) <= input(5);
output(0, 220) <= input(6);
output(0, 221) <= input(7);
output(0, 222) <= input(8);
output(0, 223) <= input(9);
output(0, 224) <= input(43);
output(0, 225) <= input(41);
output(0, 226) <= input(39);
output(0, 227) <= input(37);
output(0, 228) <= input(35);
output(0, 229) <= input(33);
output(0, 230) <= input(16);
output(0, 231) <= input(17);
output(0, 232) <= input(18);
output(0, 233) <= input(19);
output(0, 234) <= input(20);
output(0, 235) <= input(21);
output(0, 236) <= input(22);
output(0, 237) <= input(23);
output(0, 238) <= input(24);
output(0, 239) <= input(25);
output(0, 240) <= input(43);
output(0, 241) <= input(41);
output(0, 242) <= input(39);
output(0, 243) <= input(37);
output(0, 244) <= input(35);
output(0, 245) <= input(33);
output(0, 246) <= input(16);
output(0, 247) <= input(17);
output(0, 248) <= input(18);
output(0, 249) <= input(19);
output(0, 250) <= input(20);
output(0, 251) <= input(21);
output(0, 252) <= input(22);
output(0, 253) <= input(23);
output(0, 254) <= input(24);
output(0, 255) <= input(25);
output(1, 0) <= input(0);
output(1, 1) <= input(1);
output(1, 2) <= input(2);
output(1, 3) <= input(3);
output(1, 4) <= input(4);
output(1, 5) <= input(5);
output(1, 6) <= input(6);
output(1, 7) <= input(7);
output(1, 8) <= input(8);
output(1, 9) <= input(9);
output(1, 10) <= input(10);
output(1, 11) <= input(11);
output(1, 12) <= input(12);
output(1, 13) <= input(13);
output(1, 14) <= input(14);
output(1, 15) <= input(15);
output(1, 16) <= input(16);
output(1, 17) <= input(17);
output(1, 18) <= input(18);
output(1, 19) <= input(19);
output(1, 20) <= input(20);
output(1, 21) <= input(21);
output(1, 22) <= input(22);
output(1, 23) <= input(23);
output(1, 24) <= input(24);
output(1, 25) <= input(25);
output(1, 26) <= input(26);
output(1, 27) <= input(27);
output(1, 28) <= input(28);
output(1, 29) <= input(29);
output(1, 30) <= input(30);
output(1, 31) <= input(31);
output(1, 32) <= input(32);
output(1, 33) <= input(0);
output(1, 34) <= input(1);
output(1, 35) <= input(2);
output(1, 36) <= input(3);
output(1, 37) <= input(4);
output(1, 38) <= input(5);
output(1, 39) <= input(6);
output(1, 40) <= input(7);
output(1, 41) <= input(8);
output(1, 42) <= input(9);
output(1, 43) <= input(10);
output(1, 44) <= input(11);
output(1, 45) <= input(12);
output(1, 46) <= input(13);
output(1, 47) <= input(14);
output(1, 48) <= input(32);
output(1, 49) <= input(0);
output(1, 50) <= input(1);
output(1, 51) <= input(2);
output(1, 52) <= input(3);
output(1, 53) <= input(4);
output(1, 54) <= input(5);
output(1, 55) <= input(6);
output(1, 56) <= input(7);
output(1, 57) <= input(8);
output(1, 58) <= input(9);
output(1, 59) <= input(10);
output(1, 60) <= input(11);
output(1, 61) <= input(12);
output(1, 62) <= input(13);
output(1, 63) <= input(14);
output(1, 64) <= input(33);
output(1, 65) <= input(16);
output(1, 66) <= input(17);
output(1, 67) <= input(18);
output(1, 68) <= input(19);
output(1, 69) <= input(20);
output(1, 70) <= input(21);
output(1, 71) <= input(22);
output(1, 72) <= input(23);
output(1, 73) <= input(24);
output(1, 74) <= input(25);
output(1, 75) <= input(26);
output(1, 76) <= input(27);
output(1, 77) <= input(28);
output(1, 78) <= input(29);
output(1, 79) <= input(30);
output(1, 80) <= input(34);
output(1, 81) <= input(32);
output(1, 82) <= input(0);
output(1, 83) <= input(1);
output(1, 84) <= input(2);
output(1, 85) <= input(3);
output(1, 86) <= input(4);
output(1, 87) <= input(5);
output(1, 88) <= input(6);
output(1, 89) <= input(7);
output(1, 90) <= input(8);
output(1, 91) <= input(9);
output(1, 92) <= input(10);
output(1, 93) <= input(11);
output(1, 94) <= input(12);
output(1, 95) <= input(13);
output(1, 96) <= input(35);
output(1, 97) <= input(33);
output(1, 98) <= input(16);
output(1, 99) <= input(17);
output(1, 100) <= input(18);
output(1, 101) <= input(19);
output(1, 102) <= input(20);
output(1, 103) <= input(21);
output(1, 104) <= input(22);
output(1, 105) <= input(23);
output(1, 106) <= input(24);
output(1, 107) <= input(25);
output(1, 108) <= input(26);
output(1, 109) <= input(27);
output(1, 110) <= input(28);
output(1, 111) <= input(29);
output(1, 112) <= input(35);
output(1, 113) <= input(33);
output(1, 114) <= input(16);
output(1, 115) <= input(17);
output(1, 116) <= input(18);
output(1, 117) <= input(19);
output(1, 118) <= input(20);
output(1, 119) <= input(21);
output(1, 120) <= input(22);
output(1, 121) <= input(23);
output(1, 122) <= input(24);
output(1, 123) <= input(25);
output(1, 124) <= input(26);
output(1, 125) <= input(27);
output(1, 126) <= input(28);
output(1, 127) <= input(29);
output(1, 128) <= input(36);
output(1, 129) <= input(34);
output(1, 130) <= input(32);
output(1, 131) <= input(0);
output(1, 132) <= input(1);
output(1, 133) <= input(2);
output(1, 134) <= input(3);
output(1, 135) <= input(4);
output(1, 136) <= input(5);
output(1, 137) <= input(6);
output(1, 138) <= input(7);
output(1, 139) <= input(8);
output(1, 140) <= input(9);
output(1, 141) <= input(10);
output(1, 142) <= input(11);
output(1, 143) <= input(12);
output(1, 144) <= input(37);
output(1, 145) <= input(35);
output(1, 146) <= input(33);
output(1, 147) <= input(16);
output(1, 148) <= input(17);
output(1, 149) <= input(18);
output(1, 150) <= input(19);
output(1, 151) <= input(20);
output(1, 152) <= input(21);
output(1, 153) <= input(22);
output(1, 154) <= input(23);
output(1, 155) <= input(24);
output(1, 156) <= input(25);
output(1, 157) <= input(26);
output(1, 158) <= input(27);
output(1, 159) <= input(28);
output(1, 160) <= input(38);
output(1, 161) <= input(36);
output(1, 162) <= input(34);
output(1, 163) <= input(32);
output(1, 164) <= input(0);
output(1, 165) <= input(1);
output(1, 166) <= input(2);
output(1, 167) <= input(3);
output(1, 168) <= input(4);
output(1, 169) <= input(5);
output(1, 170) <= input(6);
output(1, 171) <= input(7);
output(1, 172) <= input(8);
output(1, 173) <= input(9);
output(1, 174) <= input(10);
output(1, 175) <= input(11);
output(1, 176) <= input(38);
output(1, 177) <= input(36);
output(1, 178) <= input(34);
output(1, 179) <= input(32);
output(1, 180) <= input(0);
output(1, 181) <= input(1);
output(1, 182) <= input(2);
output(1, 183) <= input(3);
output(1, 184) <= input(4);
output(1, 185) <= input(5);
output(1, 186) <= input(6);
output(1, 187) <= input(7);
output(1, 188) <= input(8);
output(1, 189) <= input(9);
output(1, 190) <= input(10);
output(1, 191) <= input(11);
output(1, 192) <= input(39);
output(1, 193) <= input(37);
output(1, 194) <= input(35);
output(1, 195) <= input(33);
output(1, 196) <= input(16);
output(1, 197) <= input(17);
output(1, 198) <= input(18);
output(1, 199) <= input(19);
output(1, 200) <= input(20);
output(1, 201) <= input(21);
output(1, 202) <= input(22);
output(1, 203) <= input(23);
output(1, 204) <= input(24);
output(1, 205) <= input(25);
output(1, 206) <= input(26);
output(1, 207) <= input(27);
output(1, 208) <= input(40);
output(1, 209) <= input(38);
output(1, 210) <= input(36);
output(1, 211) <= input(34);
output(1, 212) <= input(32);
output(1, 213) <= input(0);
output(1, 214) <= input(1);
output(1, 215) <= input(2);
output(1, 216) <= input(3);
output(1, 217) <= input(4);
output(1, 218) <= input(5);
output(1, 219) <= input(6);
output(1, 220) <= input(7);
output(1, 221) <= input(8);
output(1, 222) <= input(9);
output(1, 223) <= input(10);
output(1, 224) <= input(41);
output(1, 225) <= input(39);
output(1, 226) <= input(37);
output(1, 227) <= input(35);
output(1, 228) <= input(33);
output(1, 229) <= input(16);
output(1, 230) <= input(17);
output(1, 231) <= input(18);
output(1, 232) <= input(19);
output(1, 233) <= input(20);
output(1, 234) <= input(21);
output(1, 235) <= input(22);
output(1, 236) <= input(23);
output(1, 237) <= input(24);
output(1, 238) <= input(25);
output(1, 239) <= input(26);
output(1, 240) <= input(41);
output(1, 241) <= input(39);
output(1, 242) <= input(37);
output(1, 243) <= input(35);
output(1, 244) <= input(33);
output(1, 245) <= input(16);
output(1, 246) <= input(17);
output(1, 247) <= input(18);
output(1, 248) <= input(19);
output(1, 249) <= input(20);
output(1, 250) <= input(21);
output(1, 251) <= input(22);
output(1, 252) <= input(23);
output(1, 253) <= input(24);
output(1, 254) <= input(25);
output(1, 255) <= input(26);
output(2, 0) <= input(0);
output(2, 1) <= input(1);
output(2, 2) <= input(2);
output(2, 3) <= input(3);
output(2, 4) <= input(4);
output(2, 5) <= input(5);
output(2, 6) <= input(6);
output(2, 7) <= input(7);
output(2, 8) <= input(8);
output(2, 9) <= input(9);
output(2, 10) <= input(10);
output(2, 11) <= input(11);
output(2, 12) <= input(12);
output(2, 13) <= input(13);
output(2, 14) <= input(14);
output(2, 15) <= input(15);
output(2, 16) <= input(16);
output(2, 17) <= input(17);
output(2, 18) <= input(18);
output(2, 19) <= input(19);
output(2, 20) <= input(20);
output(2, 21) <= input(21);
output(2, 22) <= input(22);
output(2, 23) <= input(23);
output(2, 24) <= input(24);
output(2, 25) <= input(25);
output(2, 26) <= input(26);
output(2, 27) <= input(27);
output(2, 28) <= input(28);
output(2, 29) <= input(29);
output(2, 30) <= input(30);
output(2, 31) <= input(31);
output(2, 32) <= input(16);
output(2, 33) <= input(17);
output(2, 34) <= input(18);
output(2, 35) <= input(19);
output(2, 36) <= input(20);
output(2, 37) <= input(21);
output(2, 38) <= input(22);
output(2, 39) <= input(23);
output(2, 40) <= input(24);
output(2, 41) <= input(25);
output(2, 42) <= input(26);
output(2, 43) <= input(27);
output(2, 44) <= input(28);
output(2, 45) <= input(29);
output(2, 46) <= input(30);
output(2, 47) <= input(31);
output(2, 48) <= input(32);
output(2, 49) <= input(0);
output(2, 50) <= input(1);
output(2, 51) <= input(2);
output(2, 52) <= input(3);
output(2, 53) <= input(4);
output(2, 54) <= input(5);
output(2, 55) <= input(6);
output(2, 56) <= input(7);
output(2, 57) <= input(8);
output(2, 58) <= input(9);
output(2, 59) <= input(10);
output(2, 60) <= input(11);
output(2, 61) <= input(12);
output(2, 62) <= input(13);
output(2, 63) <= input(14);
output(2, 64) <= input(33);
output(2, 65) <= input(16);
output(2, 66) <= input(17);
output(2, 67) <= input(18);
output(2, 68) <= input(19);
output(2, 69) <= input(20);
output(2, 70) <= input(21);
output(2, 71) <= input(22);
output(2, 72) <= input(23);
output(2, 73) <= input(24);
output(2, 74) <= input(25);
output(2, 75) <= input(26);
output(2, 76) <= input(27);
output(2, 77) <= input(28);
output(2, 78) <= input(29);
output(2, 79) <= input(30);
output(2, 80) <= input(33);
output(2, 81) <= input(16);
output(2, 82) <= input(17);
output(2, 83) <= input(18);
output(2, 84) <= input(19);
output(2, 85) <= input(20);
output(2, 86) <= input(21);
output(2, 87) <= input(22);
output(2, 88) <= input(23);
output(2, 89) <= input(24);
output(2, 90) <= input(25);
output(2, 91) <= input(26);
output(2, 92) <= input(27);
output(2, 93) <= input(28);
output(2, 94) <= input(29);
output(2, 95) <= input(30);
output(2, 96) <= input(34);
output(2, 97) <= input(32);
output(2, 98) <= input(0);
output(2, 99) <= input(1);
output(2, 100) <= input(2);
output(2, 101) <= input(3);
output(2, 102) <= input(4);
output(2, 103) <= input(5);
output(2, 104) <= input(6);
output(2, 105) <= input(7);
output(2, 106) <= input(8);
output(2, 107) <= input(9);
output(2, 108) <= input(10);
output(2, 109) <= input(11);
output(2, 110) <= input(12);
output(2, 111) <= input(13);
output(2, 112) <= input(34);
output(2, 113) <= input(32);
output(2, 114) <= input(0);
output(2, 115) <= input(1);
output(2, 116) <= input(2);
output(2, 117) <= input(3);
output(2, 118) <= input(4);
output(2, 119) <= input(5);
output(2, 120) <= input(6);
output(2, 121) <= input(7);
output(2, 122) <= input(8);
output(2, 123) <= input(9);
output(2, 124) <= input(10);
output(2, 125) <= input(11);
output(2, 126) <= input(12);
output(2, 127) <= input(13);
output(2, 128) <= input(35);
output(2, 129) <= input(33);
output(2, 130) <= input(16);
output(2, 131) <= input(17);
output(2, 132) <= input(18);
output(2, 133) <= input(19);
output(2, 134) <= input(20);
output(2, 135) <= input(21);
output(2, 136) <= input(22);
output(2, 137) <= input(23);
output(2, 138) <= input(24);
output(2, 139) <= input(25);
output(2, 140) <= input(26);
output(2, 141) <= input(27);
output(2, 142) <= input(28);
output(2, 143) <= input(29);
output(2, 144) <= input(36);
output(2, 145) <= input(34);
output(2, 146) <= input(32);
output(2, 147) <= input(0);
output(2, 148) <= input(1);
output(2, 149) <= input(2);
output(2, 150) <= input(3);
output(2, 151) <= input(4);
output(2, 152) <= input(5);
output(2, 153) <= input(6);
output(2, 154) <= input(7);
output(2, 155) <= input(8);
output(2, 156) <= input(9);
output(2, 157) <= input(10);
output(2, 158) <= input(11);
output(2, 159) <= input(12);
output(2, 160) <= input(36);
output(2, 161) <= input(34);
output(2, 162) <= input(32);
output(2, 163) <= input(0);
output(2, 164) <= input(1);
output(2, 165) <= input(2);
output(2, 166) <= input(3);
output(2, 167) <= input(4);
output(2, 168) <= input(5);
output(2, 169) <= input(6);
output(2, 170) <= input(7);
output(2, 171) <= input(8);
output(2, 172) <= input(9);
output(2, 173) <= input(10);
output(2, 174) <= input(11);
output(2, 175) <= input(12);
output(2, 176) <= input(37);
output(2, 177) <= input(35);
output(2, 178) <= input(33);
output(2, 179) <= input(16);
output(2, 180) <= input(17);
output(2, 181) <= input(18);
output(2, 182) <= input(19);
output(2, 183) <= input(20);
output(2, 184) <= input(21);
output(2, 185) <= input(22);
output(2, 186) <= input(23);
output(2, 187) <= input(24);
output(2, 188) <= input(25);
output(2, 189) <= input(26);
output(2, 190) <= input(27);
output(2, 191) <= input(28);
output(2, 192) <= input(38);
output(2, 193) <= input(36);
output(2, 194) <= input(34);
output(2, 195) <= input(32);
output(2, 196) <= input(0);
output(2, 197) <= input(1);
output(2, 198) <= input(2);
output(2, 199) <= input(3);
output(2, 200) <= input(4);
output(2, 201) <= input(5);
output(2, 202) <= input(6);
output(2, 203) <= input(7);
output(2, 204) <= input(8);
output(2, 205) <= input(9);
output(2, 206) <= input(10);
output(2, 207) <= input(11);
output(2, 208) <= input(38);
output(2, 209) <= input(36);
output(2, 210) <= input(34);
output(2, 211) <= input(32);
output(2, 212) <= input(0);
output(2, 213) <= input(1);
output(2, 214) <= input(2);
output(2, 215) <= input(3);
output(2, 216) <= input(4);
output(2, 217) <= input(5);
output(2, 218) <= input(6);
output(2, 219) <= input(7);
output(2, 220) <= input(8);
output(2, 221) <= input(9);
output(2, 222) <= input(10);
output(2, 223) <= input(11);
output(2, 224) <= input(39);
output(2, 225) <= input(37);
output(2, 226) <= input(35);
output(2, 227) <= input(33);
output(2, 228) <= input(16);
output(2, 229) <= input(17);
output(2, 230) <= input(18);
output(2, 231) <= input(19);
output(2, 232) <= input(20);
output(2, 233) <= input(21);
output(2, 234) <= input(22);
output(2, 235) <= input(23);
output(2, 236) <= input(24);
output(2, 237) <= input(25);
output(2, 238) <= input(26);
output(2, 239) <= input(27);
output(2, 240) <= input(39);
output(2, 241) <= input(37);
output(2, 242) <= input(35);
output(2, 243) <= input(33);
output(2, 244) <= input(16);
output(2, 245) <= input(17);
output(2, 246) <= input(18);
output(2, 247) <= input(19);
output(2, 248) <= input(20);
output(2, 249) <= input(21);
output(2, 250) <= input(22);
output(2, 251) <= input(23);
output(2, 252) <= input(24);
output(2, 253) <= input(25);
output(2, 254) <= input(26);
output(2, 255) <= input(27);
when "1100" =>
output(0, 0) <= input(0);
output(0, 1) <= input(1);
output(0, 2) <= input(2);
output(0, 3) <= input(3);
output(0, 4) <= input(4);
output(0, 5) <= input(5);
output(0, 6) <= input(6);
output(0, 7) <= input(7);
output(0, 8) <= input(8);
output(0, 9) <= input(9);
output(0, 10) <= input(10);
output(0, 11) <= input(11);
output(0, 12) <= input(12);
output(0, 13) <= input(13);
output(0, 14) <= input(14);
output(0, 15) <= input(15);
output(0, 16) <= input(0);
output(0, 17) <= input(1);
output(0, 18) <= input(2);
output(0, 19) <= input(3);
output(0, 20) <= input(4);
output(0, 21) <= input(5);
output(0, 22) <= input(6);
output(0, 23) <= input(7);
output(0, 24) <= input(8);
output(0, 25) <= input(9);
output(0, 26) <= input(10);
output(0, 27) <= input(11);
output(0, 28) <= input(12);
output(0, 29) <= input(13);
output(0, 30) <= input(14);
output(0, 31) <= input(15);
output(0, 32) <= input(16);
output(0, 33) <= input(17);
output(0, 34) <= input(18);
output(0, 35) <= input(19);
output(0, 36) <= input(20);
output(0, 37) <= input(21);
output(0, 38) <= input(22);
output(0, 39) <= input(23);
output(0, 40) <= input(24);
output(0, 41) <= input(25);
output(0, 42) <= input(26);
output(0, 43) <= input(27);
output(0, 44) <= input(28);
output(0, 45) <= input(29);
output(0, 46) <= input(30);
output(0, 47) <= input(31);
output(0, 48) <= input(16);
output(0, 49) <= input(17);
output(0, 50) <= input(18);
output(0, 51) <= input(19);
output(0, 52) <= input(20);
output(0, 53) <= input(21);
output(0, 54) <= input(22);
output(0, 55) <= input(23);
output(0, 56) <= input(24);
output(0, 57) <= input(25);
output(0, 58) <= input(26);
output(0, 59) <= input(27);
output(0, 60) <= input(28);
output(0, 61) <= input(29);
output(0, 62) <= input(30);
output(0, 63) <= input(31);
output(0, 64) <= input(32);
output(0, 65) <= input(0);
output(0, 66) <= input(1);
output(0, 67) <= input(2);
output(0, 68) <= input(3);
output(0, 69) <= input(4);
output(0, 70) <= input(5);
output(0, 71) <= input(6);
output(0, 72) <= input(7);
output(0, 73) <= input(8);
output(0, 74) <= input(9);
output(0, 75) <= input(10);
output(0, 76) <= input(11);
output(0, 77) <= input(12);
output(0, 78) <= input(13);
output(0, 79) <= input(14);
output(0, 80) <= input(32);
output(0, 81) <= input(0);
output(0, 82) <= input(1);
output(0, 83) <= input(2);
output(0, 84) <= input(3);
output(0, 85) <= input(4);
output(0, 86) <= input(5);
output(0, 87) <= input(6);
output(0, 88) <= input(7);
output(0, 89) <= input(8);
output(0, 90) <= input(9);
output(0, 91) <= input(10);
output(0, 92) <= input(11);
output(0, 93) <= input(12);
output(0, 94) <= input(13);
output(0, 95) <= input(14);
output(0, 96) <= input(33);
output(0, 97) <= input(16);
output(0, 98) <= input(17);
output(0, 99) <= input(18);
output(0, 100) <= input(19);
output(0, 101) <= input(20);
output(0, 102) <= input(21);
output(0, 103) <= input(22);
output(0, 104) <= input(23);
output(0, 105) <= input(24);
output(0, 106) <= input(25);
output(0, 107) <= input(26);
output(0, 108) <= input(27);
output(0, 109) <= input(28);
output(0, 110) <= input(29);
output(0, 111) <= input(30);
output(0, 112) <= input(33);
output(0, 113) <= input(16);
output(0, 114) <= input(17);
output(0, 115) <= input(18);
output(0, 116) <= input(19);
output(0, 117) <= input(20);
output(0, 118) <= input(21);
output(0, 119) <= input(22);
output(0, 120) <= input(23);
output(0, 121) <= input(24);
output(0, 122) <= input(25);
output(0, 123) <= input(26);
output(0, 124) <= input(27);
output(0, 125) <= input(28);
output(0, 126) <= input(29);
output(0, 127) <= input(30);
output(0, 128) <= input(34);
output(0, 129) <= input(32);
output(0, 130) <= input(0);
output(0, 131) <= input(1);
output(0, 132) <= input(2);
output(0, 133) <= input(3);
output(0, 134) <= input(4);
output(0, 135) <= input(5);
output(0, 136) <= input(6);
output(0, 137) <= input(7);
output(0, 138) <= input(8);
output(0, 139) <= input(9);
output(0, 140) <= input(10);
output(0, 141) <= input(11);
output(0, 142) <= input(12);
output(0, 143) <= input(13);
output(0, 144) <= input(34);
output(0, 145) <= input(32);
output(0, 146) <= input(0);
output(0, 147) <= input(1);
output(0, 148) <= input(2);
output(0, 149) <= input(3);
output(0, 150) <= input(4);
output(0, 151) <= input(5);
output(0, 152) <= input(6);
output(0, 153) <= input(7);
output(0, 154) <= input(8);
output(0, 155) <= input(9);
output(0, 156) <= input(10);
output(0, 157) <= input(11);
output(0, 158) <= input(12);
output(0, 159) <= input(13);
output(0, 160) <= input(35);
output(0, 161) <= input(33);
output(0, 162) <= input(16);
output(0, 163) <= input(17);
output(0, 164) <= input(18);
output(0, 165) <= input(19);
output(0, 166) <= input(20);
output(0, 167) <= input(21);
output(0, 168) <= input(22);
output(0, 169) <= input(23);
output(0, 170) <= input(24);
output(0, 171) <= input(25);
output(0, 172) <= input(26);
output(0, 173) <= input(27);
output(0, 174) <= input(28);
output(0, 175) <= input(29);
output(0, 176) <= input(35);
output(0, 177) <= input(33);
output(0, 178) <= input(16);
output(0, 179) <= input(17);
output(0, 180) <= input(18);
output(0, 181) <= input(19);
output(0, 182) <= input(20);
output(0, 183) <= input(21);
output(0, 184) <= input(22);
output(0, 185) <= input(23);
output(0, 186) <= input(24);
output(0, 187) <= input(25);
output(0, 188) <= input(26);
output(0, 189) <= input(27);
output(0, 190) <= input(28);
output(0, 191) <= input(29);
output(0, 192) <= input(36);
output(0, 193) <= input(34);
output(0, 194) <= input(32);
output(0, 195) <= input(0);
output(0, 196) <= input(1);
output(0, 197) <= input(2);
output(0, 198) <= input(3);
output(0, 199) <= input(4);
output(0, 200) <= input(5);
output(0, 201) <= input(6);
output(0, 202) <= input(7);
output(0, 203) <= input(8);
output(0, 204) <= input(9);
output(0, 205) <= input(10);
output(0, 206) <= input(11);
output(0, 207) <= input(12);
output(0, 208) <= input(36);
output(0, 209) <= input(34);
output(0, 210) <= input(32);
output(0, 211) <= input(0);
output(0, 212) <= input(1);
output(0, 213) <= input(2);
output(0, 214) <= input(3);
output(0, 215) <= input(4);
output(0, 216) <= input(5);
output(0, 217) <= input(6);
output(0, 218) <= input(7);
output(0, 219) <= input(8);
output(0, 220) <= input(9);
output(0, 221) <= input(10);
output(0, 222) <= input(11);
output(0, 223) <= input(12);
output(0, 224) <= input(37);
output(0, 225) <= input(35);
output(0, 226) <= input(33);
output(0, 227) <= input(16);
output(0, 228) <= input(17);
output(0, 229) <= input(18);
output(0, 230) <= input(19);
output(0, 231) <= input(20);
output(0, 232) <= input(21);
output(0, 233) <= input(22);
output(0, 234) <= input(23);
output(0, 235) <= input(24);
output(0, 236) <= input(25);
output(0, 237) <= input(26);
output(0, 238) <= input(27);
output(0, 239) <= input(28);
output(0, 240) <= input(37);
output(0, 241) <= input(35);
output(0, 242) <= input(33);
output(0, 243) <= input(16);
output(0, 244) <= input(17);
output(0, 245) <= input(18);
output(0, 246) <= input(19);
output(0, 247) <= input(20);
output(0, 248) <= input(21);
output(0, 249) <= input(22);
output(0, 250) <= input(23);
output(0, 251) <= input(24);
output(0, 252) <= input(25);
output(0, 253) <= input(26);
output(0, 254) <= input(27);
output(0, 255) <= input(28);
output(1, 0) <= input(0);
output(1, 1) <= input(1);
output(1, 2) <= input(2);
output(1, 3) <= input(3);
output(1, 4) <= input(4);
output(1, 5) <= input(5);
output(1, 6) <= input(6);
output(1, 7) <= input(7);
output(1, 8) <= input(8);
output(1, 9) <= input(9);
output(1, 10) <= input(10);
output(1, 11) <= input(11);
output(1, 12) <= input(12);
output(1, 13) <= input(13);
output(1, 14) <= input(14);
output(1, 15) <= input(15);
output(1, 16) <= input(0);
output(1, 17) <= input(1);
output(1, 18) <= input(2);
output(1, 19) <= input(3);
output(1, 20) <= input(4);
output(1, 21) <= input(5);
output(1, 22) <= input(6);
output(1, 23) <= input(7);
output(1, 24) <= input(8);
output(1, 25) <= input(9);
output(1, 26) <= input(10);
output(1, 27) <= input(11);
output(1, 28) <= input(12);
output(1, 29) <= input(13);
output(1, 30) <= input(14);
output(1, 31) <= input(15);
output(1, 32) <= input(16);
output(1, 33) <= input(17);
output(1, 34) <= input(18);
output(1, 35) <= input(19);
output(1, 36) <= input(20);
output(1, 37) <= input(21);
output(1, 38) <= input(22);
output(1, 39) <= input(23);
output(1, 40) <= input(24);
output(1, 41) <= input(25);
output(1, 42) <= input(26);
output(1, 43) <= input(27);
output(1, 44) <= input(28);
output(1, 45) <= input(29);
output(1, 46) <= input(30);
output(1, 47) <= input(31);
output(1, 48) <= input(16);
output(1, 49) <= input(17);
output(1, 50) <= input(18);
output(1, 51) <= input(19);
output(1, 52) <= input(20);
output(1, 53) <= input(21);
output(1, 54) <= input(22);
output(1, 55) <= input(23);
output(1, 56) <= input(24);
output(1, 57) <= input(25);
output(1, 58) <= input(26);
output(1, 59) <= input(27);
output(1, 60) <= input(28);
output(1, 61) <= input(29);
output(1, 62) <= input(30);
output(1, 63) <= input(31);
output(1, 64) <= input(16);
output(1, 65) <= input(17);
output(1, 66) <= input(18);
output(1, 67) <= input(19);
output(1, 68) <= input(20);
output(1, 69) <= input(21);
output(1, 70) <= input(22);
output(1, 71) <= input(23);
output(1, 72) <= input(24);
output(1, 73) <= input(25);
output(1, 74) <= input(26);
output(1, 75) <= input(27);
output(1, 76) <= input(28);
output(1, 77) <= input(29);
output(1, 78) <= input(30);
output(1, 79) <= input(31);
output(1, 80) <= input(32);
output(1, 81) <= input(0);
output(1, 82) <= input(1);
output(1, 83) <= input(2);
output(1, 84) <= input(3);
output(1, 85) <= input(4);
output(1, 86) <= input(5);
output(1, 87) <= input(6);
output(1, 88) <= input(7);
output(1, 89) <= input(8);
output(1, 90) <= input(9);
output(1, 91) <= input(10);
output(1, 92) <= input(11);
output(1, 93) <= input(12);
output(1, 94) <= input(13);
output(1, 95) <= input(14);
output(1, 96) <= input(32);
output(1, 97) <= input(0);
output(1, 98) <= input(1);
output(1, 99) <= input(2);
output(1, 100) <= input(3);
output(1, 101) <= input(4);
output(1, 102) <= input(5);
output(1, 103) <= input(6);
output(1, 104) <= input(7);
output(1, 105) <= input(8);
output(1, 106) <= input(9);
output(1, 107) <= input(10);
output(1, 108) <= input(11);
output(1, 109) <= input(12);
output(1, 110) <= input(13);
output(1, 111) <= input(14);
output(1, 112) <= input(32);
output(1, 113) <= input(0);
output(1, 114) <= input(1);
output(1, 115) <= input(2);
output(1, 116) <= input(3);
output(1, 117) <= input(4);
output(1, 118) <= input(5);
output(1, 119) <= input(6);
output(1, 120) <= input(7);
output(1, 121) <= input(8);
output(1, 122) <= input(9);
output(1, 123) <= input(10);
output(1, 124) <= input(11);
output(1, 125) <= input(12);
output(1, 126) <= input(13);
output(1, 127) <= input(14);
output(1, 128) <= input(33);
output(1, 129) <= input(16);
output(1, 130) <= input(17);
output(1, 131) <= input(18);
output(1, 132) <= input(19);
output(1, 133) <= input(20);
output(1, 134) <= input(21);
output(1, 135) <= input(22);
output(1, 136) <= input(23);
output(1, 137) <= input(24);
output(1, 138) <= input(25);
output(1, 139) <= input(26);
output(1, 140) <= input(27);
output(1, 141) <= input(28);
output(1, 142) <= input(29);
output(1, 143) <= input(30);
output(1, 144) <= input(33);
output(1, 145) <= input(16);
output(1, 146) <= input(17);
output(1, 147) <= input(18);
output(1, 148) <= input(19);
output(1, 149) <= input(20);
output(1, 150) <= input(21);
output(1, 151) <= input(22);
output(1, 152) <= input(23);
output(1, 153) <= input(24);
output(1, 154) <= input(25);
output(1, 155) <= input(26);
output(1, 156) <= input(27);
output(1, 157) <= input(28);
output(1, 158) <= input(29);
output(1, 159) <= input(30);
output(1, 160) <= input(34);
output(1, 161) <= input(32);
output(1, 162) <= input(0);
output(1, 163) <= input(1);
output(1, 164) <= input(2);
output(1, 165) <= input(3);
output(1, 166) <= input(4);
output(1, 167) <= input(5);
output(1, 168) <= input(6);
output(1, 169) <= input(7);
output(1, 170) <= input(8);
output(1, 171) <= input(9);
output(1, 172) <= input(10);
output(1, 173) <= input(11);
output(1, 174) <= input(12);
output(1, 175) <= input(13);
output(1, 176) <= input(34);
output(1, 177) <= input(32);
output(1, 178) <= input(0);
output(1, 179) <= input(1);
output(1, 180) <= input(2);
output(1, 181) <= input(3);
output(1, 182) <= input(4);
output(1, 183) <= input(5);
output(1, 184) <= input(6);
output(1, 185) <= input(7);
output(1, 186) <= input(8);
output(1, 187) <= input(9);
output(1, 188) <= input(10);
output(1, 189) <= input(11);
output(1, 190) <= input(12);
output(1, 191) <= input(13);
output(1, 192) <= input(34);
output(1, 193) <= input(32);
output(1, 194) <= input(0);
output(1, 195) <= input(1);
output(1, 196) <= input(2);
output(1, 197) <= input(3);
output(1, 198) <= input(4);
output(1, 199) <= input(5);
output(1, 200) <= input(6);
output(1, 201) <= input(7);
output(1, 202) <= input(8);
output(1, 203) <= input(9);
output(1, 204) <= input(10);
output(1, 205) <= input(11);
output(1, 206) <= input(12);
output(1, 207) <= input(13);
output(1, 208) <= input(35);
output(1, 209) <= input(33);
output(1, 210) <= input(16);
output(1, 211) <= input(17);
output(1, 212) <= input(18);
output(1, 213) <= input(19);
output(1, 214) <= input(20);
output(1, 215) <= input(21);
output(1, 216) <= input(22);
output(1, 217) <= input(23);
output(1, 218) <= input(24);
output(1, 219) <= input(25);
output(1, 220) <= input(26);
output(1, 221) <= input(27);
output(1, 222) <= input(28);
output(1, 223) <= input(29);
output(1, 224) <= input(35);
output(1, 225) <= input(33);
output(1, 226) <= input(16);
output(1, 227) <= input(17);
output(1, 228) <= input(18);
output(1, 229) <= input(19);
output(1, 230) <= input(20);
output(1, 231) <= input(21);
output(1, 232) <= input(22);
output(1, 233) <= input(23);
output(1, 234) <= input(24);
output(1, 235) <= input(25);
output(1, 236) <= input(26);
output(1, 237) <= input(27);
output(1, 238) <= input(28);
output(1, 239) <= input(29);
output(1, 240) <= input(35);
output(1, 241) <= input(33);
output(1, 242) <= input(16);
output(1, 243) <= input(17);
output(1, 244) <= input(18);
output(1, 245) <= input(19);
output(1, 246) <= input(20);
output(1, 247) <= input(21);
output(1, 248) <= input(22);
output(1, 249) <= input(23);
output(1, 250) <= input(24);
output(1, 251) <= input(25);
output(1, 252) <= input(26);
output(1, 253) <= input(27);
output(1, 254) <= input(28);
output(1, 255) <= input(29);
output(2, 0) <= input(0);
output(2, 1) <= input(1);
output(2, 2) <= input(2);
output(2, 3) <= input(3);
output(2, 4) <= input(4);
output(2, 5) <= input(5);
output(2, 6) <= input(6);
output(2, 7) <= input(7);
output(2, 8) <= input(8);
output(2, 9) <= input(9);
output(2, 10) <= input(10);
output(2, 11) <= input(11);
output(2, 12) <= input(12);
output(2, 13) <= input(13);
output(2, 14) <= input(14);
output(2, 15) <= input(15);
output(2, 16) <= input(0);
output(2, 17) <= input(1);
output(2, 18) <= input(2);
output(2, 19) <= input(3);
output(2, 20) <= input(4);
output(2, 21) <= input(5);
output(2, 22) <= input(6);
output(2, 23) <= input(7);
output(2, 24) <= input(8);
output(2, 25) <= input(9);
output(2, 26) <= input(10);
output(2, 27) <= input(11);
output(2, 28) <= input(12);
output(2, 29) <= input(13);
output(2, 30) <= input(14);
output(2, 31) <= input(15);
output(2, 32) <= input(0);
output(2, 33) <= input(1);
output(2, 34) <= input(2);
output(2, 35) <= input(3);
output(2, 36) <= input(4);
output(2, 37) <= input(5);
output(2, 38) <= input(6);
output(2, 39) <= input(7);
output(2, 40) <= input(8);
output(2, 41) <= input(9);
output(2, 42) <= input(10);
output(2, 43) <= input(11);
output(2, 44) <= input(12);
output(2, 45) <= input(13);
output(2, 46) <= input(14);
output(2, 47) <= input(15);
output(2, 48) <= input(0);
output(2, 49) <= input(1);
output(2, 50) <= input(2);
output(2, 51) <= input(3);
output(2, 52) <= input(4);
output(2, 53) <= input(5);
output(2, 54) <= input(6);
output(2, 55) <= input(7);
output(2, 56) <= input(8);
output(2, 57) <= input(9);
output(2, 58) <= input(10);
output(2, 59) <= input(11);
output(2, 60) <= input(12);
output(2, 61) <= input(13);
output(2, 62) <= input(14);
output(2, 63) <= input(15);
output(2, 64) <= input(16);
output(2, 65) <= input(17);
output(2, 66) <= input(18);
output(2, 67) <= input(19);
output(2, 68) <= input(20);
output(2, 69) <= input(21);
output(2, 70) <= input(22);
output(2, 71) <= input(23);
output(2, 72) <= input(24);
output(2, 73) <= input(25);
output(2, 74) <= input(26);
output(2, 75) <= input(27);
output(2, 76) <= input(28);
output(2, 77) <= input(29);
output(2, 78) <= input(30);
output(2, 79) <= input(31);
output(2, 80) <= input(16);
output(2, 81) <= input(17);
output(2, 82) <= input(18);
output(2, 83) <= input(19);
output(2, 84) <= input(20);
output(2, 85) <= input(21);
output(2, 86) <= input(22);
output(2, 87) <= input(23);
output(2, 88) <= input(24);
output(2, 89) <= input(25);
output(2, 90) <= input(26);
output(2, 91) <= input(27);
output(2, 92) <= input(28);
output(2, 93) <= input(29);
output(2, 94) <= input(30);
output(2, 95) <= input(31);
output(2, 96) <= input(16);
output(2, 97) <= input(17);
output(2, 98) <= input(18);
output(2, 99) <= input(19);
output(2, 100) <= input(20);
output(2, 101) <= input(21);
output(2, 102) <= input(22);
output(2, 103) <= input(23);
output(2, 104) <= input(24);
output(2, 105) <= input(25);
output(2, 106) <= input(26);
output(2, 107) <= input(27);
output(2, 108) <= input(28);
output(2, 109) <= input(29);
output(2, 110) <= input(30);
output(2, 111) <= input(31);
output(2, 112) <= input(16);
output(2, 113) <= input(17);
output(2, 114) <= input(18);
output(2, 115) <= input(19);
output(2, 116) <= input(20);
output(2, 117) <= input(21);
output(2, 118) <= input(22);
output(2, 119) <= input(23);
output(2, 120) <= input(24);
output(2, 121) <= input(25);
output(2, 122) <= input(26);
output(2, 123) <= input(27);
output(2, 124) <= input(28);
output(2, 125) <= input(29);
output(2, 126) <= input(30);
output(2, 127) <= input(31);
output(2, 128) <= input(32);
output(2, 129) <= input(0);
output(2, 130) <= input(1);
output(2, 131) <= input(2);
output(2, 132) <= input(3);
output(2, 133) <= input(4);
output(2, 134) <= input(5);
output(2, 135) <= input(6);
output(2, 136) <= input(7);
output(2, 137) <= input(8);
output(2, 138) <= input(9);
output(2, 139) <= input(10);
output(2, 140) <= input(11);
output(2, 141) <= input(12);
output(2, 142) <= input(13);
output(2, 143) <= input(14);
output(2, 144) <= input(32);
output(2, 145) <= input(0);
output(2, 146) <= input(1);
output(2, 147) <= input(2);
output(2, 148) <= input(3);
output(2, 149) <= input(4);
output(2, 150) <= input(5);
output(2, 151) <= input(6);
output(2, 152) <= input(7);
output(2, 153) <= input(8);
output(2, 154) <= input(9);
output(2, 155) <= input(10);
output(2, 156) <= input(11);
output(2, 157) <= input(12);
output(2, 158) <= input(13);
output(2, 159) <= input(14);
output(2, 160) <= input(32);
output(2, 161) <= input(0);
output(2, 162) <= input(1);
output(2, 163) <= input(2);
output(2, 164) <= input(3);
output(2, 165) <= input(4);
output(2, 166) <= input(5);
output(2, 167) <= input(6);
output(2, 168) <= input(7);
output(2, 169) <= input(8);
output(2, 170) <= input(9);
output(2, 171) <= input(10);
output(2, 172) <= input(11);
output(2, 173) <= input(12);
output(2, 174) <= input(13);
output(2, 175) <= input(14);
output(2, 176) <= input(32);
output(2, 177) <= input(0);
output(2, 178) <= input(1);
output(2, 179) <= input(2);
output(2, 180) <= input(3);
output(2, 181) <= input(4);
output(2, 182) <= input(5);
output(2, 183) <= input(6);
output(2, 184) <= input(7);
output(2, 185) <= input(8);
output(2, 186) <= input(9);
output(2, 187) <= input(10);
output(2, 188) <= input(11);
output(2, 189) <= input(12);
output(2, 190) <= input(13);
output(2, 191) <= input(14);
output(2, 192) <= input(33);
output(2, 193) <= input(16);
output(2, 194) <= input(17);
output(2, 195) <= input(18);
output(2, 196) <= input(19);
output(2, 197) <= input(20);
output(2, 198) <= input(21);
output(2, 199) <= input(22);
output(2, 200) <= input(23);
output(2, 201) <= input(24);
output(2, 202) <= input(25);
output(2, 203) <= input(26);
output(2, 204) <= input(27);
output(2, 205) <= input(28);
output(2, 206) <= input(29);
output(2, 207) <= input(30);
output(2, 208) <= input(33);
output(2, 209) <= input(16);
output(2, 210) <= input(17);
output(2, 211) <= input(18);
output(2, 212) <= input(19);
output(2, 213) <= input(20);
output(2, 214) <= input(21);
output(2, 215) <= input(22);
output(2, 216) <= input(23);
output(2, 217) <= input(24);
output(2, 218) <= input(25);
output(2, 219) <= input(26);
output(2, 220) <= input(27);
output(2, 221) <= input(28);
output(2, 222) <= input(29);
output(2, 223) <= input(30);
output(2, 224) <= input(33);
output(2, 225) <= input(16);
output(2, 226) <= input(17);
output(2, 227) <= input(18);
output(2, 228) <= input(19);
output(2, 229) <= input(20);
output(2, 230) <= input(21);
output(2, 231) <= input(22);
output(2, 232) <= input(23);
output(2, 233) <= input(24);
output(2, 234) <= input(25);
output(2, 235) <= input(26);
output(2, 236) <= input(27);
output(2, 237) <= input(28);
output(2, 238) <= input(29);
output(2, 239) <= input(30);
output(2, 240) <= input(33);
output(2, 241) <= input(16);
output(2, 242) <= input(17);
output(2, 243) <= input(18);
output(2, 244) <= input(19);
output(2, 245) <= input(20);
output(2, 246) <= input(21);
output(2, 247) <= input(22);
output(2, 248) <= input(23);
output(2, 249) <= input(24);
output(2, 250) <= input(25);
output(2, 251) <= input(26);
output(2, 252) <= input(27);
output(2, 253) <= input(28);
output(2, 254) <= input(29);
output(2, 255) <= input(30);
when "1101" =>
output(0, 0) <= input(0);
output(0, 1) <= input(1);
output(0, 2) <= input(2);
output(0, 3) <= input(3);
output(0, 4) <= input(4);
output(0, 5) <= input(5);
output(0, 6) <= input(6);
output(0, 7) <= input(7);
output(0, 8) <= input(8);
output(0, 9) <= input(9);
output(0, 10) <= input(10);
output(0, 11) <= input(11);
output(0, 12) <= input(12);
output(0, 13) <= input(13);
output(0, 14) <= input(14);
output(0, 15) <= input(15);
output(0, 16) <= input(0);
output(0, 17) <= input(1);
output(0, 18) <= input(2);
output(0, 19) <= input(3);
output(0, 20) <= input(4);
output(0, 21) <= input(5);
output(0, 22) <= input(6);
output(0, 23) <= input(7);
output(0, 24) <= input(8);
output(0, 25) <= input(9);
output(0, 26) <= input(10);
output(0, 27) <= input(11);
output(0, 28) <= input(12);
output(0, 29) <= input(13);
output(0, 30) <= input(14);
output(0, 31) <= input(15);
output(0, 32) <= input(0);
output(0, 33) <= input(1);
output(0, 34) <= input(2);
output(0, 35) <= input(3);
output(0, 36) <= input(4);
output(0, 37) <= input(5);
output(0, 38) <= input(6);
output(0, 39) <= input(7);
output(0, 40) <= input(8);
output(0, 41) <= input(9);
output(0, 42) <= input(10);
output(0, 43) <= input(11);
output(0, 44) <= input(12);
output(0, 45) <= input(13);
output(0, 46) <= input(14);
output(0, 47) <= input(15);
output(0, 48) <= input(0);
output(0, 49) <= input(1);
output(0, 50) <= input(2);
output(0, 51) <= input(3);
output(0, 52) <= input(4);
output(0, 53) <= input(5);
output(0, 54) <= input(6);
output(0, 55) <= input(7);
output(0, 56) <= input(8);
output(0, 57) <= input(9);
output(0, 58) <= input(10);
output(0, 59) <= input(11);
output(0, 60) <= input(12);
output(0, 61) <= input(13);
output(0, 62) <= input(14);
output(0, 63) <= input(15);
output(0, 64) <= input(0);
output(0, 65) <= input(1);
output(0, 66) <= input(2);
output(0, 67) <= input(3);
output(0, 68) <= input(4);
output(0, 69) <= input(5);
output(0, 70) <= input(6);
output(0, 71) <= input(7);
output(0, 72) <= input(8);
output(0, 73) <= input(9);
output(0, 74) <= input(10);
output(0, 75) <= input(11);
output(0, 76) <= input(12);
output(0, 77) <= input(13);
output(0, 78) <= input(14);
output(0, 79) <= input(15);
output(0, 80) <= input(16);
output(0, 81) <= input(17);
output(0, 82) <= input(18);
output(0, 83) <= input(19);
output(0, 84) <= input(20);
output(0, 85) <= input(21);
output(0, 86) <= input(22);
output(0, 87) <= input(23);
output(0, 88) <= input(24);
output(0, 89) <= input(25);
output(0, 90) <= input(26);
output(0, 91) <= input(27);
output(0, 92) <= input(28);
output(0, 93) <= input(29);
output(0, 94) <= input(30);
output(0, 95) <= input(31);
output(0, 96) <= input(16);
output(0, 97) <= input(17);
output(0, 98) <= input(18);
output(0, 99) <= input(19);
output(0, 100) <= input(20);
output(0, 101) <= input(21);
output(0, 102) <= input(22);
output(0, 103) <= input(23);
output(0, 104) <= input(24);
output(0, 105) <= input(25);
output(0, 106) <= input(26);
output(0, 107) <= input(27);
output(0, 108) <= input(28);
output(0, 109) <= input(29);
output(0, 110) <= input(30);
output(0, 111) <= input(31);
output(0, 112) <= input(16);
output(0, 113) <= input(17);
output(0, 114) <= input(18);
output(0, 115) <= input(19);
output(0, 116) <= input(20);
output(0, 117) <= input(21);
output(0, 118) <= input(22);
output(0, 119) <= input(23);
output(0, 120) <= input(24);
output(0, 121) <= input(25);
output(0, 122) <= input(26);
output(0, 123) <= input(27);
output(0, 124) <= input(28);
output(0, 125) <= input(29);
output(0, 126) <= input(30);
output(0, 127) <= input(31);
output(0, 128) <= input(16);
output(0, 129) <= input(17);
output(0, 130) <= input(18);
output(0, 131) <= input(19);
output(0, 132) <= input(20);
output(0, 133) <= input(21);
output(0, 134) <= input(22);
output(0, 135) <= input(23);
output(0, 136) <= input(24);
output(0, 137) <= input(25);
output(0, 138) <= input(26);
output(0, 139) <= input(27);
output(0, 140) <= input(28);
output(0, 141) <= input(29);
output(0, 142) <= input(30);
output(0, 143) <= input(31);
output(0, 144) <= input(16);
output(0, 145) <= input(17);
output(0, 146) <= input(18);
output(0, 147) <= input(19);
output(0, 148) <= input(20);
output(0, 149) <= input(21);
output(0, 150) <= input(22);
output(0, 151) <= input(23);
output(0, 152) <= input(24);
output(0, 153) <= input(25);
output(0, 154) <= input(26);
output(0, 155) <= input(27);
output(0, 156) <= input(28);
output(0, 157) <= input(29);
output(0, 158) <= input(30);
output(0, 159) <= input(31);
output(0, 160) <= input(32);
output(0, 161) <= input(0);
output(0, 162) <= input(1);
output(0, 163) <= input(2);
output(0, 164) <= input(3);
output(0, 165) <= input(4);
output(0, 166) <= input(5);
output(0, 167) <= input(6);
output(0, 168) <= input(7);
output(0, 169) <= input(8);
output(0, 170) <= input(9);
output(0, 171) <= input(10);
output(0, 172) <= input(11);
output(0, 173) <= input(12);
output(0, 174) <= input(13);
output(0, 175) <= input(14);
output(0, 176) <= input(32);
output(0, 177) <= input(0);
output(0, 178) <= input(1);
output(0, 179) <= input(2);
output(0, 180) <= input(3);
output(0, 181) <= input(4);
output(0, 182) <= input(5);
output(0, 183) <= input(6);
output(0, 184) <= input(7);
output(0, 185) <= input(8);
output(0, 186) <= input(9);
output(0, 187) <= input(10);
output(0, 188) <= input(11);
output(0, 189) <= input(12);
output(0, 190) <= input(13);
output(0, 191) <= input(14);
output(0, 192) <= input(32);
output(0, 193) <= input(0);
output(0, 194) <= input(1);
output(0, 195) <= input(2);
output(0, 196) <= input(3);
output(0, 197) <= input(4);
output(0, 198) <= input(5);
output(0, 199) <= input(6);
output(0, 200) <= input(7);
output(0, 201) <= input(8);
output(0, 202) <= input(9);
output(0, 203) <= input(10);
output(0, 204) <= input(11);
output(0, 205) <= input(12);
output(0, 206) <= input(13);
output(0, 207) <= input(14);
output(0, 208) <= input(32);
output(0, 209) <= input(0);
output(0, 210) <= input(1);
output(0, 211) <= input(2);
output(0, 212) <= input(3);
output(0, 213) <= input(4);
output(0, 214) <= input(5);
output(0, 215) <= input(6);
output(0, 216) <= input(7);
output(0, 217) <= input(8);
output(0, 218) <= input(9);
output(0, 219) <= input(10);
output(0, 220) <= input(11);
output(0, 221) <= input(12);
output(0, 222) <= input(13);
output(0, 223) <= input(14);
output(0, 224) <= input(32);
output(0, 225) <= input(0);
output(0, 226) <= input(1);
output(0, 227) <= input(2);
output(0, 228) <= input(3);
output(0, 229) <= input(4);
output(0, 230) <= input(5);
output(0, 231) <= input(6);
output(0, 232) <= input(7);
output(0, 233) <= input(8);
output(0, 234) <= input(9);
output(0, 235) <= input(10);
output(0, 236) <= input(11);
output(0, 237) <= input(12);
output(0, 238) <= input(13);
output(0, 239) <= input(14);
output(0, 240) <= input(32);
output(0, 241) <= input(0);
output(0, 242) <= input(1);
output(0, 243) <= input(2);
output(0, 244) <= input(3);
output(0, 245) <= input(4);
output(0, 246) <= input(5);
output(0, 247) <= input(6);
output(0, 248) <= input(7);
output(0, 249) <= input(8);
output(0, 250) <= input(9);
output(0, 251) <= input(10);
output(0, 252) <= input(11);
output(0, 253) <= input(12);
output(0, 254) <= input(13);
output(0, 255) <= input(14);
output(1, 0) <= input(0);
output(1, 1) <= input(1);
output(1, 2) <= input(2);
output(1, 3) <= input(3);
output(1, 4) <= input(4);
output(1, 5) <= input(5);
output(1, 6) <= input(6);
output(1, 7) <= input(7);
output(1, 8) <= input(8);
output(1, 9) <= input(9);
output(1, 10) <= input(10);
output(1, 11) <= input(11);
output(1, 12) <= input(12);
output(1, 13) <= input(13);
output(1, 14) <= input(14);
output(1, 15) <= input(15);
output(1, 16) <= input(0);
output(1, 17) <= input(1);
output(1, 18) <= input(2);
output(1, 19) <= input(3);
output(1, 20) <= input(4);
output(1, 21) <= input(5);
output(1, 22) <= input(6);
output(1, 23) <= input(7);
output(1, 24) <= input(8);
output(1, 25) <= input(9);
output(1, 26) <= input(10);
output(1, 27) <= input(11);
output(1, 28) <= input(12);
output(1, 29) <= input(13);
output(1, 30) <= input(14);
output(1, 31) <= input(15);
output(1, 32) <= input(0);
output(1, 33) <= input(1);
output(1, 34) <= input(2);
output(1, 35) <= input(3);
output(1, 36) <= input(4);
output(1, 37) <= input(5);
output(1, 38) <= input(6);
output(1, 39) <= input(7);
output(1, 40) <= input(8);
output(1, 41) <= input(9);
output(1, 42) <= input(10);
output(1, 43) <= input(11);
output(1, 44) <= input(12);
output(1, 45) <= input(13);
output(1, 46) <= input(14);
output(1, 47) <= input(15);
output(1, 48) <= input(0);
output(1, 49) <= input(1);
output(1, 50) <= input(2);
output(1, 51) <= input(3);
output(1, 52) <= input(4);
output(1, 53) <= input(5);
output(1, 54) <= input(6);
output(1, 55) <= input(7);
output(1, 56) <= input(8);
output(1, 57) <= input(9);
output(1, 58) <= input(10);
output(1, 59) <= input(11);
output(1, 60) <= input(12);
output(1, 61) <= input(13);
output(1, 62) <= input(14);
output(1, 63) <= input(15);
output(1, 64) <= input(0);
output(1, 65) <= input(1);
output(1, 66) <= input(2);
output(1, 67) <= input(3);
output(1, 68) <= input(4);
output(1, 69) <= input(5);
output(1, 70) <= input(6);
output(1, 71) <= input(7);
output(1, 72) <= input(8);
output(1, 73) <= input(9);
output(1, 74) <= input(10);
output(1, 75) <= input(11);
output(1, 76) <= input(12);
output(1, 77) <= input(13);
output(1, 78) <= input(14);
output(1, 79) <= input(15);
output(1, 80) <= input(0);
output(1, 81) <= input(1);
output(1, 82) <= input(2);
output(1, 83) <= input(3);
output(1, 84) <= input(4);
output(1, 85) <= input(5);
output(1, 86) <= input(6);
output(1, 87) <= input(7);
output(1, 88) <= input(8);
output(1, 89) <= input(9);
output(1, 90) <= input(10);
output(1, 91) <= input(11);
output(1, 92) <= input(12);
output(1, 93) <= input(13);
output(1, 94) <= input(14);
output(1, 95) <= input(15);
output(1, 96) <= input(0);
output(1, 97) <= input(1);
output(1, 98) <= input(2);
output(1, 99) <= input(3);
output(1, 100) <= input(4);
output(1, 101) <= input(5);
output(1, 102) <= input(6);
output(1, 103) <= input(7);
output(1, 104) <= input(8);
output(1, 105) <= input(9);
output(1, 106) <= input(10);
output(1, 107) <= input(11);
output(1, 108) <= input(12);
output(1, 109) <= input(13);
output(1, 110) <= input(14);
output(1, 111) <= input(15);
output(1, 112) <= input(0);
output(1, 113) <= input(1);
output(1, 114) <= input(2);
output(1, 115) <= input(3);
output(1, 116) <= input(4);
output(1, 117) <= input(5);
output(1, 118) <= input(6);
output(1, 119) <= input(7);
output(1, 120) <= input(8);
output(1, 121) <= input(9);
output(1, 122) <= input(10);
output(1, 123) <= input(11);
output(1, 124) <= input(12);
output(1, 125) <= input(13);
output(1, 126) <= input(14);
output(1, 127) <= input(15);
output(1, 128) <= input(16);
output(1, 129) <= input(17);
output(1, 130) <= input(18);
output(1, 131) <= input(19);
output(1, 132) <= input(20);
output(1, 133) <= input(21);
output(1, 134) <= input(22);
output(1, 135) <= input(23);
output(1, 136) <= input(24);
output(1, 137) <= input(25);
output(1, 138) <= input(26);
output(1, 139) <= input(27);
output(1, 140) <= input(28);
output(1, 141) <= input(29);
output(1, 142) <= input(30);
output(1, 143) <= input(31);
output(1, 144) <= input(16);
output(1, 145) <= input(17);
output(1, 146) <= input(18);
output(1, 147) <= input(19);
output(1, 148) <= input(20);
output(1, 149) <= input(21);
output(1, 150) <= input(22);
output(1, 151) <= input(23);
output(1, 152) <= input(24);
output(1, 153) <= input(25);
output(1, 154) <= input(26);
output(1, 155) <= input(27);
output(1, 156) <= input(28);
output(1, 157) <= input(29);
output(1, 158) <= input(30);
output(1, 159) <= input(31);
output(1, 160) <= input(16);
output(1, 161) <= input(17);
output(1, 162) <= input(18);
output(1, 163) <= input(19);
output(1, 164) <= input(20);
output(1, 165) <= input(21);
output(1, 166) <= input(22);
output(1, 167) <= input(23);
output(1, 168) <= input(24);
output(1, 169) <= input(25);
output(1, 170) <= input(26);
output(1, 171) <= input(27);
output(1, 172) <= input(28);
output(1, 173) <= input(29);
output(1, 174) <= input(30);
output(1, 175) <= input(31);
output(1, 176) <= input(16);
output(1, 177) <= input(17);
output(1, 178) <= input(18);
output(1, 179) <= input(19);
output(1, 180) <= input(20);
output(1, 181) <= input(21);
output(1, 182) <= input(22);
output(1, 183) <= input(23);
output(1, 184) <= input(24);
output(1, 185) <= input(25);
output(1, 186) <= input(26);
output(1, 187) <= input(27);
output(1, 188) <= input(28);
output(1, 189) <= input(29);
output(1, 190) <= input(30);
output(1, 191) <= input(31);
output(1, 192) <= input(16);
output(1, 193) <= input(17);
output(1, 194) <= input(18);
output(1, 195) <= input(19);
output(1, 196) <= input(20);
output(1, 197) <= input(21);
output(1, 198) <= input(22);
output(1, 199) <= input(23);
output(1, 200) <= input(24);
output(1, 201) <= input(25);
output(1, 202) <= input(26);
output(1, 203) <= input(27);
output(1, 204) <= input(28);
output(1, 205) <= input(29);
output(1, 206) <= input(30);
output(1, 207) <= input(31);
output(1, 208) <= input(16);
output(1, 209) <= input(17);
output(1, 210) <= input(18);
output(1, 211) <= input(19);
output(1, 212) <= input(20);
output(1, 213) <= input(21);
output(1, 214) <= input(22);
output(1, 215) <= input(23);
output(1, 216) <= input(24);
output(1, 217) <= input(25);
output(1, 218) <= input(26);
output(1, 219) <= input(27);
output(1, 220) <= input(28);
output(1, 221) <= input(29);
output(1, 222) <= input(30);
output(1, 223) <= input(31);
output(1, 224) <= input(16);
output(1, 225) <= input(17);
output(1, 226) <= input(18);
output(1, 227) <= input(19);
output(1, 228) <= input(20);
output(1, 229) <= input(21);
output(1, 230) <= input(22);
output(1, 231) <= input(23);
output(1, 232) <= input(24);
output(1, 233) <= input(25);
output(1, 234) <= input(26);
output(1, 235) <= input(27);
output(1, 236) <= input(28);
output(1, 237) <= input(29);
output(1, 238) <= input(30);
output(1, 239) <= input(31);
output(1, 240) <= input(16);
output(1, 241) <= input(17);
output(1, 242) <= input(18);
output(1, 243) <= input(19);
output(1, 244) <= input(20);
output(1, 245) <= input(21);
output(1, 246) <= input(22);
output(1, 247) <= input(23);
output(1, 248) <= input(24);
output(1, 249) <= input(25);
output(1, 250) <= input(26);
output(1, 251) <= input(27);
output(1, 252) <= input(28);
output(1, 253) <= input(29);
output(1, 254) <= input(30);
output(1, 255) <= input(31);
output(2, 0) <= input(0);
output(2, 1) <= input(1);
output(2, 2) <= input(2);
output(2, 3) <= input(3);
output(2, 4) <= input(4);
output(2, 5) <= input(5);
output(2, 6) <= input(6);
output(2, 7) <= input(7);
output(2, 8) <= input(8);
output(2, 9) <= input(9);
output(2, 10) <= input(10);
output(2, 11) <= input(11);
output(2, 12) <= input(12);
output(2, 13) <= input(13);
output(2, 14) <= input(14);
output(2, 15) <= input(15);
output(2, 16) <= input(0);
output(2, 17) <= input(1);
output(2, 18) <= input(2);
output(2, 19) <= input(3);
output(2, 20) <= input(4);
output(2, 21) <= input(5);
output(2, 22) <= input(6);
output(2, 23) <= input(7);
output(2, 24) <= input(8);
output(2, 25) <= input(9);
output(2, 26) <= input(10);
output(2, 27) <= input(11);
output(2, 28) <= input(12);
output(2, 29) <= input(13);
output(2, 30) <= input(14);
output(2, 31) <= input(15);
output(2, 32) <= input(0);
output(2, 33) <= input(1);
output(2, 34) <= input(2);
output(2, 35) <= input(3);
output(2, 36) <= input(4);
output(2, 37) <= input(5);
output(2, 38) <= input(6);
output(2, 39) <= input(7);
output(2, 40) <= input(8);
output(2, 41) <= input(9);
output(2, 42) <= input(10);
output(2, 43) <= input(11);
output(2, 44) <= input(12);
output(2, 45) <= input(13);
output(2, 46) <= input(14);
output(2, 47) <= input(15);
output(2, 48) <= input(0);
output(2, 49) <= input(1);
output(2, 50) <= input(2);
output(2, 51) <= input(3);
output(2, 52) <= input(4);
output(2, 53) <= input(5);
output(2, 54) <= input(6);
output(2, 55) <= input(7);
output(2, 56) <= input(8);
output(2, 57) <= input(9);
output(2, 58) <= input(10);
output(2, 59) <= input(11);
output(2, 60) <= input(12);
output(2, 61) <= input(13);
output(2, 62) <= input(14);
output(2, 63) <= input(15);
output(2, 64) <= input(0);
output(2, 65) <= input(1);
output(2, 66) <= input(2);
output(2, 67) <= input(3);
output(2, 68) <= input(4);
output(2, 69) <= input(5);
output(2, 70) <= input(6);
output(2, 71) <= input(7);
output(2, 72) <= input(8);
output(2, 73) <= input(9);
output(2, 74) <= input(10);
output(2, 75) <= input(11);
output(2, 76) <= input(12);
output(2, 77) <= input(13);
output(2, 78) <= input(14);
output(2, 79) <= input(15);
output(2, 80) <= input(0);
output(2, 81) <= input(1);
output(2, 82) <= input(2);
output(2, 83) <= input(3);
output(2, 84) <= input(4);
output(2, 85) <= input(5);
output(2, 86) <= input(6);
output(2, 87) <= input(7);
output(2, 88) <= input(8);
output(2, 89) <= input(9);
output(2, 90) <= input(10);
output(2, 91) <= input(11);
output(2, 92) <= input(12);
output(2, 93) <= input(13);
output(2, 94) <= input(14);
output(2, 95) <= input(15);
output(2, 96) <= input(0);
output(2, 97) <= input(1);
output(2, 98) <= input(2);
output(2, 99) <= input(3);
output(2, 100) <= input(4);
output(2, 101) <= input(5);
output(2, 102) <= input(6);
output(2, 103) <= input(7);
output(2, 104) <= input(8);
output(2, 105) <= input(9);
output(2, 106) <= input(10);
output(2, 107) <= input(11);
output(2, 108) <= input(12);
output(2, 109) <= input(13);
output(2, 110) <= input(14);
output(2, 111) <= input(15);
output(2, 112) <= input(0);
output(2, 113) <= input(1);
output(2, 114) <= input(2);
output(2, 115) <= input(3);
output(2, 116) <= input(4);
output(2, 117) <= input(5);
output(2, 118) <= input(6);
output(2, 119) <= input(7);
output(2, 120) <= input(8);
output(2, 121) <= input(9);
output(2, 122) <= input(10);
output(2, 123) <= input(11);
output(2, 124) <= input(12);
output(2, 125) <= input(13);
output(2, 126) <= input(14);
output(2, 127) <= input(15);
output(2, 128) <= input(0);
output(2, 129) <= input(1);
output(2, 130) <= input(2);
output(2, 131) <= input(3);
output(2, 132) <= input(4);
output(2, 133) <= input(5);
output(2, 134) <= input(6);
output(2, 135) <= input(7);
output(2, 136) <= input(8);
output(2, 137) <= input(9);
output(2, 138) <= input(10);
output(2, 139) <= input(11);
output(2, 140) <= input(12);
output(2, 141) <= input(13);
output(2, 142) <= input(14);
output(2, 143) <= input(15);
output(2, 144) <= input(0);
output(2, 145) <= input(1);
output(2, 146) <= input(2);
output(2, 147) <= input(3);
output(2, 148) <= input(4);
output(2, 149) <= input(5);
output(2, 150) <= input(6);
output(2, 151) <= input(7);
output(2, 152) <= input(8);
output(2, 153) <= input(9);
output(2, 154) <= input(10);
output(2, 155) <= input(11);
output(2, 156) <= input(12);
output(2, 157) <= input(13);
output(2, 158) <= input(14);
output(2, 159) <= input(15);
output(2, 160) <= input(0);
output(2, 161) <= input(1);
output(2, 162) <= input(2);
output(2, 163) <= input(3);
output(2, 164) <= input(4);
output(2, 165) <= input(5);
output(2, 166) <= input(6);
output(2, 167) <= input(7);
output(2, 168) <= input(8);
output(2, 169) <= input(9);
output(2, 170) <= input(10);
output(2, 171) <= input(11);
output(2, 172) <= input(12);
output(2, 173) <= input(13);
output(2, 174) <= input(14);
output(2, 175) <= input(15);
output(2, 176) <= input(0);
output(2, 177) <= input(1);
output(2, 178) <= input(2);
output(2, 179) <= input(3);
output(2, 180) <= input(4);
output(2, 181) <= input(5);
output(2, 182) <= input(6);
output(2, 183) <= input(7);
output(2, 184) <= input(8);
output(2, 185) <= input(9);
output(2, 186) <= input(10);
output(2, 187) <= input(11);
output(2, 188) <= input(12);
output(2, 189) <= input(13);
output(2, 190) <= input(14);
output(2, 191) <= input(15);
output(2, 192) <= input(0);
output(2, 193) <= input(1);
output(2, 194) <= input(2);
output(2, 195) <= input(3);
output(2, 196) <= input(4);
output(2, 197) <= input(5);
output(2, 198) <= input(6);
output(2, 199) <= input(7);
output(2, 200) <= input(8);
output(2, 201) <= input(9);
output(2, 202) <= input(10);
output(2, 203) <= input(11);
output(2, 204) <= input(12);
output(2, 205) <= input(13);
output(2, 206) <= input(14);
output(2, 207) <= input(15);
output(2, 208) <= input(0);
output(2, 209) <= input(1);
output(2, 210) <= input(2);
output(2, 211) <= input(3);
output(2, 212) <= input(4);
output(2, 213) <= input(5);
output(2, 214) <= input(6);
output(2, 215) <= input(7);
output(2, 216) <= input(8);
output(2, 217) <= input(9);
output(2, 218) <= input(10);
output(2, 219) <= input(11);
output(2, 220) <= input(12);
output(2, 221) <= input(13);
output(2, 222) <= input(14);
output(2, 223) <= input(15);
output(2, 224) <= input(0);
output(2, 225) <= input(1);
output(2, 226) <= input(2);
output(2, 227) <= input(3);
output(2, 228) <= input(4);
output(2, 229) <= input(5);
output(2, 230) <= input(6);
output(2, 231) <= input(7);
output(2, 232) <= input(8);
output(2, 233) <= input(9);
output(2, 234) <= input(10);
output(2, 235) <= input(11);
output(2, 236) <= input(12);
output(2, 237) <= input(13);
output(2, 238) <= input(14);
output(2, 239) <= input(15);
output(2, 240) <= input(0);
output(2, 241) <= input(1);
output(2, 242) <= input(2);
output(2, 243) <= input(3);
output(2, 244) <= input(4);
output(2, 245) <= input(5);
output(2, 246) <= input(6);
output(2, 247) <= input(7);
output(2, 248) <= input(8);
output(2, 249) <= input(9);
output(2, 250) <= input(10);
output(2, 251) <= input(11);
output(2, 252) <= input(12);
output(2, 253) <= input(13);
output(2, 254) <= input(14);
output(2, 255) <= input(15);
output(3, 0) <= input(17);
output(3, 1) <= input(18);
output(3, 2) <= input(19);
output(3, 3) <= input(20);
output(3, 4) <= input(21);
output(3, 5) <= input(22);
output(3, 6) <= input(23);
output(3, 7) <= input(24);
output(3, 8) <= input(25);
output(3, 9) <= input(26);
output(3, 10) <= input(27);
output(3, 11) <= input(28);
output(3, 12) <= input(29);
output(3, 13) <= input(30);
output(3, 14) <= input(31);
output(3, 15) <= input(33);
output(3, 16) <= input(17);
output(3, 17) <= input(18);
output(3, 18) <= input(19);
output(3, 19) <= input(20);
output(3, 20) <= input(21);
output(3, 21) <= input(22);
output(3, 22) <= input(23);
output(3, 23) <= input(24);
output(3, 24) <= input(25);
output(3, 25) <= input(26);
output(3, 26) <= input(27);
output(3, 27) <= input(28);
output(3, 28) <= input(29);
output(3, 29) <= input(30);
output(3, 30) <= input(31);
output(3, 31) <= input(33);
output(3, 32) <= input(17);
output(3, 33) <= input(18);
output(3, 34) <= input(19);
output(3, 35) <= input(20);
output(3, 36) <= input(21);
output(3, 37) <= input(22);
output(3, 38) <= input(23);
output(3, 39) <= input(24);
output(3, 40) <= input(25);
output(3, 41) <= input(26);
output(3, 42) <= input(27);
output(3, 43) <= input(28);
output(3, 44) <= input(29);
output(3, 45) <= input(30);
output(3, 46) <= input(31);
output(3, 47) <= input(33);
output(3, 48) <= input(17);
output(3, 49) <= input(18);
output(3, 50) <= input(19);
output(3, 51) <= input(20);
output(3, 52) <= input(21);
output(3, 53) <= input(22);
output(3, 54) <= input(23);
output(3, 55) <= input(24);
output(3, 56) <= input(25);
output(3, 57) <= input(26);
output(3, 58) <= input(27);
output(3, 59) <= input(28);
output(3, 60) <= input(29);
output(3, 61) <= input(30);
output(3, 62) <= input(31);
output(3, 63) <= input(33);
output(3, 64) <= input(17);
output(3, 65) <= input(18);
output(3, 66) <= input(19);
output(3, 67) <= input(20);
output(3, 68) <= input(21);
output(3, 69) <= input(22);
output(3, 70) <= input(23);
output(3, 71) <= input(24);
output(3, 72) <= input(25);
output(3, 73) <= input(26);
output(3, 74) <= input(27);
output(3, 75) <= input(28);
output(3, 76) <= input(29);
output(3, 77) <= input(30);
output(3, 78) <= input(31);
output(3, 79) <= input(33);
output(3, 80) <= input(17);
output(3, 81) <= input(18);
output(3, 82) <= input(19);
output(3, 83) <= input(20);
output(3, 84) <= input(21);
output(3, 85) <= input(22);
output(3, 86) <= input(23);
output(3, 87) <= input(24);
output(3, 88) <= input(25);
output(3, 89) <= input(26);
output(3, 90) <= input(27);
output(3, 91) <= input(28);
output(3, 92) <= input(29);
output(3, 93) <= input(30);
output(3, 94) <= input(31);
output(3, 95) <= input(33);
output(3, 96) <= input(17);
output(3, 97) <= input(18);
output(3, 98) <= input(19);
output(3, 99) <= input(20);
output(3, 100) <= input(21);
output(3, 101) <= input(22);
output(3, 102) <= input(23);
output(3, 103) <= input(24);
output(3, 104) <= input(25);
output(3, 105) <= input(26);
output(3, 106) <= input(27);
output(3, 107) <= input(28);
output(3, 108) <= input(29);
output(3, 109) <= input(30);
output(3, 110) <= input(31);
output(3, 111) <= input(33);
output(3, 112) <= input(17);
output(3, 113) <= input(18);
output(3, 114) <= input(19);
output(3, 115) <= input(20);
output(3, 116) <= input(21);
output(3, 117) <= input(22);
output(3, 118) <= input(23);
output(3, 119) <= input(24);
output(3, 120) <= input(25);
output(3, 121) <= input(26);
output(3, 122) <= input(27);
output(3, 123) <= input(28);
output(3, 124) <= input(29);
output(3, 125) <= input(30);
output(3, 126) <= input(31);
output(3, 127) <= input(33);
output(3, 128) <= input(17);
output(3, 129) <= input(18);
output(3, 130) <= input(19);
output(3, 131) <= input(20);
output(3, 132) <= input(21);
output(3, 133) <= input(22);
output(3, 134) <= input(23);
output(3, 135) <= input(24);
output(3, 136) <= input(25);
output(3, 137) <= input(26);
output(3, 138) <= input(27);
output(3, 139) <= input(28);
output(3, 140) <= input(29);
output(3, 141) <= input(30);
output(3, 142) <= input(31);
output(3, 143) <= input(33);
output(3, 144) <= input(17);
output(3, 145) <= input(18);
output(3, 146) <= input(19);
output(3, 147) <= input(20);
output(3, 148) <= input(21);
output(3, 149) <= input(22);
output(3, 150) <= input(23);
output(3, 151) <= input(24);
output(3, 152) <= input(25);
output(3, 153) <= input(26);
output(3, 154) <= input(27);
output(3, 155) <= input(28);
output(3, 156) <= input(29);
output(3, 157) <= input(30);
output(3, 158) <= input(31);
output(3, 159) <= input(33);
output(3, 160) <= input(17);
output(3, 161) <= input(18);
output(3, 162) <= input(19);
output(3, 163) <= input(20);
output(3, 164) <= input(21);
output(3, 165) <= input(22);
output(3, 166) <= input(23);
output(3, 167) <= input(24);
output(3, 168) <= input(25);
output(3, 169) <= input(26);
output(3, 170) <= input(27);
output(3, 171) <= input(28);
output(3, 172) <= input(29);
output(3, 173) <= input(30);
output(3, 174) <= input(31);
output(3, 175) <= input(33);
output(3, 176) <= input(17);
output(3, 177) <= input(18);
output(3, 178) <= input(19);
output(3, 179) <= input(20);
output(3, 180) <= input(21);
output(3, 181) <= input(22);
output(3, 182) <= input(23);
output(3, 183) <= input(24);
output(3, 184) <= input(25);
output(3, 185) <= input(26);
output(3, 186) <= input(27);
output(3, 187) <= input(28);
output(3, 188) <= input(29);
output(3, 189) <= input(30);
output(3, 190) <= input(31);
output(3, 191) <= input(33);
output(3, 192) <= input(17);
output(3, 193) <= input(18);
output(3, 194) <= input(19);
output(3, 195) <= input(20);
output(3, 196) <= input(21);
output(3, 197) <= input(22);
output(3, 198) <= input(23);
output(3, 199) <= input(24);
output(3, 200) <= input(25);
output(3, 201) <= input(26);
output(3, 202) <= input(27);
output(3, 203) <= input(28);
output(3, 204) <= input(29);
output(3, 205) <= input(30);
output(3, 206) <= input(31);
output(3, 207) <= input(33);
output(3, 208) <= input(17);
output(3, 209) <= input(18);
output(3, 210) <= input(19);
output(3, 211) <= input(20);
output(3, 212) <= input(21);
output(3, 213) <= input(22);
output(3, 214) <= input(23);
output(3, 215) <= input(24);
output(3, 216) <= input(25);
output(3, 217) <= input(26);
output(3, 218) <= input(27);
output(3, 219) <= input(28);
output(3, 220) <= input(29);
output(3, 221) <= input(30);
output(3, 222) <= input(31);
output(3, 223) <= input(33);
output(3, 224) <= input(17);
output(3, 225) <= input(18);
output(3, 226) <= input(19);
output(3, 227) <= input(20);
output(3, 228) <= input(21);
output(3, 229) <= input(22);
output(3, 230) <= input(23);
output(3, 231) <= input(24);
output(3, 232) <= input(25);
output(3, 233) <= input(26);
output(3, 234) <= input(27);
output(3, 235) <= input(28);
output(3, 236) <= input(29);
output(3, 237) <= input(30);
output(3, 238) <= input(31);
output(3, 239) <= input(33);
output(3, 240) <= input(17);
output(3, 241) <= input(18);
output(3, 242) <= input(19);
output(3, 243) <= input(20);
output(3, 244) <= input(21);
output(3, 245) <= input(22);
output(3, 246) <= input(23);
output(3, 247) <= input(24);
output(3, 248) <= input(25);
output(3, 249) <= input(26);
output(3, 250) <= input(27);
output(3, 251) <= input(28);
output(3, 252) <= input(29);
output(3, 253) <= input(30);
output(3, 254) <= input(31);
output(3, 255) <= input(33);
output(4, 0) <= input(17);
output(4, 1) <= input(18);
output(4, 2) <= input(19);
output(4, 3) <= input(20);
output(4, 4) <= input(21);
output(4, 5) <= input(22);
output(4, 6) <= input(23);
output(4, 7) <= input(24);
output(4, 8) <= input(25);
output(4, 9) <= input(26);
output(4, 10) <= input(27);
output(4, 11) <= input(28);
output(4, 12) <= input(29);
output(4, 13) <= input(30);
output(4, 14) <= input(31);
output(4, 15) <= input(33);
output(4, 16) <= input(17);
output(4, 17) <= input(18);
output(4, 18) <= input(19);
output(4, 19) <= input(20);
output(4, 20) <= input(21);
output(4, 21) <= input(22);
output(4, 22) <= input(23);
output(4, 23) <= input(24);
output(4, 24) <= input(25);
output(4, 25) <= input(26);
output(4, 26) <= input(27);
output(4, 27) <= input(28);
output(4, 28) <= input(29);
output(4, 29) <= input(30);
output(4, 30) <= input(31);
output(4, 31) <= input(33);
output(4, 32) <= input(17);
output(4, 33) <= input(18);
output(4, 34) <= input(19);
output(4, 35) <= input(20);
output(4, 36) <= input(21);
output(4, 37) <= input(22);
output(4, 38) <= input(23);
output(4, 39) <= input(24);
output(4, 40) <= input(25);
output(4, 41) <= input(26);
output(4, 42) <= input(27);
output(4, 43) <= input(28);
output(4, 44) <= input(29);
output(4, 45) <= input(30);
output(4, 46) <= input(31);
output(4, 47) <= input(33);
output(4, 48) <= input(17);
output(4, 49) <= input(18);
output(4, 50) <= input(19);
output(4, 51) <= input(20);
output(4, 52) <= input(21);
output(4, 53) <= input(22);
output(4, 54) <= input(23);
output(4, 55) <= input(24);
output(4, 56) <= input(25);
output(4, 57) <= input(26);
output(4, 58) <= input(27);
output(4, 59) <= input(28);
output(4, 60) <= input(29);
output(4, 61) <= input(30);
output(4, 62) <= input(31);
output(4, 63) <= input(33);
output(4, 64) <= input(17);
output(4, 65) <= input(18);
output(4, 66) <= input(19);
output(4, 67) <= input(20);
output(4, 68) <= input(21);
output(4, 69) <= input(22);
output(4, 70) <= input(23);
output(4, 71) <= input(24);
output(4, 72) <= input(25);
output(4, 73) <= input(26);
output(4, 74) <= input(27);
output(4, 75) <= input(28);
output(4, 76) <= input(29);
output(4, 77) <= input(30);
output(4, 78) <= input(31);
output(4, 79) <= input(33);
output(4, 80) <= input(17);
output(4, 81) <= input(18);
output(4, 82) <= input(19);
output(4, 83) <= input(20);
output(4, 84) <= input(21);
output(4, 85) <= input(22);
output(4, 86) <= input(23);
output(4, 87) <= input(24);
output(4, 88) <= input(25);
output(4, 89) <= input(26);
output(4, 90) <= input(27);
output(4, 91) <= input(28);
output(4, 92) <= input(29);
output(4, 93) <= input(30);
output(4, 94) <= input(31);
output(4, 95) <= input(33);
output(4, 96) <= input(17);
output(4, 97) <= input(18);
output(4, 98) <= input(19);
output(4, 99) <= input(20);
output(4, 100) <= input(21);
output(4, 101) <= input(22);
output(4, 102) <= input(23);
output(4, 103) <= input(24);
output(4, 104) <= input(25);
output(4, 105) <= input(26);
output(4, 106) <= input(27);
output(4, 107) <= input(28);
output(4, 108) <= input(29);
output(4, 109) <= input(30);
output(4, 110) <= input(31);
output(4, 111) <= input(33);
output(4, 112) <= input(17);
output(4, 113) <= input(18);
output(4, 114) <= input(19);
output(4, 115) <= input(20);
output(4, 116) <= input(21);
output(4, 117) <= input(22);
output(4, 118) <= input(23);
output(4, 119) <= input(24);
output(4, 120) <= input(25);
output(4, 121) <= input(26);
output(4, 122) <= input(27);
output(4, 123) <= input(28);
output(4, 124) <= input(29);
output(4, 125) <= input(30);
output(4, 126) <= input(31);
output(4, 127) <= input(33);
output(4, 128) <= input(17);
output(4, 129) <= input(18);
output(4, 130) <= input(19);
output(4, 131) <= input(20);
output(4, 132) <= input(21);
output(4, 133) <= input(22);
output(4, 134) <= input(23);
output(4, 135) <= input(24);
output(4, 136) <= input(25);
output(4, 137) <= input(26);
output(4, 138) <= input(27);
output(4, 139) <= input(28);
output(4, 140) <= input(29);
output(4, 141) <= input(30);
output(4, 142) <= input(31);
output(4, 143) <= input(33);
output(4, 144) <= input(17);
output(4, 145) <= input(18);
output(4, 146) <= input(19);
output(4, 147) <= input(20);
output(4, 148) <= input(21);
output(4, 149) <= input(22);
output(4, 150) <= input(23);
output(4, 151) <= input(24);
output(4, 152) <= input(25);
output(4, 153) <= input(26);
output(4, 154) <= input(27);
output(4, 155) <= input(28);
output(4, 156) <= input(29);
output(4, 157) <= input(30);
output(4, 158) <= input(31);
output(4, 159) <= input(33);
output(4, 160) <= input(17);
output(4, 161) <= input(18);
output(4, 162) <= input(19);
output(4, 163) <= input(20);
output(4, 164) <= input(21);
output(4, 165) <= input(22);
output(4, 166) <= input(23);
output(4, 167) <= input(24);
output(4, 168) <= input(25);
output(4, 169) <= input(26);
output(4, 170) <= input(27);
output(4, 171) <= input(28);
output(4, 172) <= input(29);
output(4, 173) <= input(30);
output(4, 174) <= input(31);
output(4, 175) <= input(33);
output(4, 176) <= input(17);
output(4, 177) <= input(18);
output(4, 178) <= input(19);
output(4, 179) <= input(20);
output(4, 180) <= input(21);
output(4, 181) <= input(22);
output(4, 182) <= input(23);
output(4, 183) <= input(24);
output(4, 184) <= input(25);
output(4, 185) <= input(26);
output(4, 186) <= input(27);
output(4, 187) <= input(28);
output(4, 188) <= input(29);
output(4, 189) <= input(30);
output(4, 190) <= input(31);
output(4, 191) <= input(33);
output(4, 192) <= input(17);
output(4, 193) <= input(18);
output(4, 194) <= input(19);
output(4, 195) <= input(20);
output(4, 196) <= input(21);
output(4, 197) <= input(22);
output(4, 198) <= input(23);
output(4, 199) <= input(24);
output(4, 200) <= input(25);
output(4, 201) <= input(26);
output(4, 202) <= input(27);
output(4, 203) <= input(28);
output(4, 204) <= input(29);
output(4, 205) <= input(30);
output(4, 206) <= input(31);
output(4, 207) <= input(33);
output(4, 208) <= input(17);
output(4, 209) <= input(18);
output(4, 210) <= input(19);
output(4, 211) <= input(20);
output(4, 212) <= input(21);
output(4, 213) <= input(22);
output(4, 214) <= input(23);
output(4, 215) <= input(24);
output(4, 216) <= input(25);
output(4, 217) <= input(26);
output(4, 218) <= input(27);
output(4, 219) <= input(28);
output(4, 220) <= input(29);
output(4, 221) <= input(30);
output(4, 222) <= input(31);
output(4, 223) <= input(33);
output(4, 224) <= input(17);
output(4, 225) <= input(18);
output(4, 226) <= input(19);
output(4, 227) <= input(20);
output(4, 228) <= input(21);
output(4, 229) <= input(22);
output(4, 230) <= input(23);
output(4, 231) <= input(24);
output(4, 232) <= input(25);
output(4, 233) <= input(26);
output(4, 234) <= input(27);
output(4, 235) <= input(28);
output(4, 236) <= input(29);
output(4, 237) <= input(30);
output(4, 238) <= input(31);
output(4, 239) <= input(33);
output(4, 240) <= input(1);
output(4, 241) <= input(2);
output(4, 242) <= input(3);
output(4, 243) <= input(4);
output(4, 244) <= input(5);
output(4, 245) <= input(6);
output(4, 246) <= input(7);
output(4, 247) <= input(8);
output(4, 248) <= input(9);
output(4, 249) <= input(10);
output(4, 250) <= input(11);
output(4, 251) <= input(12);
output(4, 252) <= input(13);
output(4, 253) <= input(14);
output(4, 254) <= input(15);
output(4, 255) <= input(34);
output(5, 0) <= input(17);
output(5, 1) <= input(18);
output(5, 2) <= input(19);
output(5, 3) <= input(20);
output(5, 4) <= input(21);
output(5, 5) <= input(22);
output(5, 6) <= input(23);
output(5, 7) <= input(24);
output(5, 8) <= input(25);
output(5, 9) <= input(26);
output(5, 10) <= input(27);
output(5, 11) <= input(28);
output(5, 12) <= input(29);
output(5, 13) <= input(30);
output(5, 14) <= input(31);
output(5, 15) <= input(33);
output(5, 16) <= input(17);
output(5, 17) <= input(18);
output(5, 18) <= input(19);
output(5, 19) <= input(20);
output(5, 20) <= input(21);
output(5, 21) <= input(22);
output(5, 22) <= input(23);
output(5, 23) <= input(24);
output(5, 24) <= input(25);
output(5, 25) <= input(26);
output(5, 26) <= input(27);
output(5, 27) <= input(28);
output(5, 28) <= input(29);
output(5, 29) <= input(30);
output(5, 30) <= input(31);
output(5, 31) <= input(33);
output(5, 32) <= input(17);
output(5, 33) <= input(18);
output(5, 34) <= input(19);
output(5, 35) <= input(20);
output(5, 36) <= input(21);
output(5, 37) <= input(22);
output(5, 38) <= input(23);
output(5, 39) <= input(24);
output(5, 40) <= input(25);
output(5, 41) <= input(26);
output(5, 42) <= input(27);
output(5, 43) <= input(28);
output(5, 44) <= input(29);
output(5, 45) <= input(30);
output(5, 46) <= input(31);
output(5, 47) <= input(33);
output(5, 48) <= input(17);
output(5, 49) <= input(18);
output(5, 50) <= input(19);
output(5, 51) <= input(20);
output(5, 52) <= input(21);
output(5, 53) <= input(22);
output(5, 54) <= input(23);
output(5, 55) <= input(24);
output(5, 56) <= input(25);
output(5, 57) <= input(26);
output(5, 58) <= input(27);
output(5, 59) <= input(28);
output(5, 60) <= input(29);
output(5, 61) <= input(30);
output(5, 62) <= input(31);
output(5, 63) <= input(33);
output(5, 64) <= input(17);
output(5, 65) <= input(18);
output(5, 66) <= input(19);
output(5, 67) <= input(20);
output(5, 68) <= input(21);
output(5, 69) <= input(22);
output(5, 70) <= input(23);
output(5, 71) <= input(24);
output(5, 72) <= input(25);
output(5, 73) <= input(26);
output(5, 74) <= input(27);
output(5, 75) <= input(28);
output(5, 76) <= input(29);
output(5, 77) <= input(30);
output(5, 78) <= input(31);
output(5, 79) <= input(33);
output(5, 80) <= input(17);
output(5, 81) <= input(18);
output(5, 82) <= input(19);
output(5, 83) <= input(20);
output(5, 84) <= input(21);
output(5, 85) <= input(22);
output(5, 86) <= input(23);
output(5, 87) <= input(24);
output(5, 88) <= input(25);
output(5, 89) <= input(26);
output(5, 90) <= input(27);
output(5, 91) <= input(28);
output(5, 92) <= input(29);
output(5, 93) <= input(30);
output(5, 94) <= input(31);
output(5, 95) <= input(33);
output(5, 96) <= input(17);
output(5, 97) <= input(18);
output(5, 98) <= input(19);
output(5, 99) <= input(20);
output(5, 100) <= input(21);
output(5, 101) <= input(22);
output(5, 102) <= input(23);
output(5, 103) <= input(24);
output(5, 104) <= input(25);
output(5, 105) <= input(26);
output(5, 106) <= input(27);
output(5, 107) <= input(28);
output(5, 108) <= input(29);
output(5, 109) <= input(30);
output(5, 110) <= input(31);
output(5, 111) <= input(33);
output(5, 112) <= input(1);
output(5, 113) <= input(2);
output(5, 114) <= input(3);
output(5, 115) <= input(4);
output(5, 116) <= input(5);
output(5, 117) <= input(6);
output(5, 118) <= input(7);
output(5, 119) <= input(8);
output(5, 120) <= input(9);
output(5, 121) <= input(10);
output(5, 122) <= input(11);
output(5, 123) <= input(12);
output(5, 124) <= input(13);
output(5, 125) <= input(14);
output(5, 126) <= input(15);
output(5, 127) <= input(34);
output(5, 128) <= input(1);
output(5, 129) <= input(2);
output(5, 130) <= input(3);
output(5, 131) <= input(4);
output(5, 132) <= input(5);
output(5, 133) <= input(6);
output(5, 134) <= input(7);
output(5, 135) <= input(8);
output(5, 136) <= input(9);
output(5, 137) <= input(10);
output(5, 138) <= input(11);
output(5, 139) <= input(12);
output(5, 140) <= input(13);
output(5, 141) <= input(14);
output(5, 142) <= input(15);
output(5, 143) <= input(34);
output(5, 144) <= input(1);
output(5, 145) <= input(2);
output(5, 146) <= input(3);
output(5, 147) <= input(4);
output(5, 148) <= input(5);
output(5, 149) <= input(6);
output(5, 150) <= input(7);
output(5, 151) <= input(8);
output(5, 152) <= input(9);
output(5, 153) <= input(10);
output(5, 154) <= input(11);
output(5, 155) <= input(12);
output(5, 156) <= input(13);
output(5, 157) <= input(14);
output(5, 158) <= input(15);
output(5, 159) <= input(34);
output(5, 160) <= input(1);
output(5, 161) <= input(2);
output(5, 162) <= input(3);
output(5, 163) <= input(4);
output(5, 164) <= input(5);
output(5, 165) <= input(6);
output(5, 166) <= input(7);
output(5, 167) <= input(8);
output(5, 168) <= input(9);
output(5, 169) <= input(10);
output(5, 170) <= input(11);
output(5, 171) <= input(12);
output(5, 172) <= input(13);
output(5, 173) <= input(14);
output(5, 174) <= input(15);
output(5, 175) <= input(34);
output(5, 176) <= input(1);
output(5, 177) <= input(2);
output(5, 178) <= input(3);
output(5, 179) <= input(4);
output(5, 180) <= input(5);
output(5, 181) <= input(6);
output(5, 182) <= input(7);
output(5, 183) <= input(8);
output(5, 184) <= input(9);
output(5, 185) <= input(10);
output(5, 186) <= input(11);
output(5, 187) <= input(12);
output(5, 188) <= input(13);
output(5, 189) <= input(14);
output(5, 190) <= input(15);
output(5, 191) <= input(34);
output(5, 192) <= input(1);
output(5, 193) <= input(2);
output(5, 194) <= input(3);
output(5, 195) <= input(4);
output(5, 196) <= input(5);
output(5, 197) <= input(6);
output(5, 198) <= input(7);
output(5, 199) <= input(8);
output(5, 200) <= input(9);
output(5, 201) <= input(10);
output(5, 202) <= input(11);
output(5, 203) <= input(12);
output(5, 204) <= input(13);
output(5, 205) <= input(14);
output(5, 206) <= input(15);
output(5, 207) <= input(34);
output(5, 208) <= input(1);
output(5, 209) <= input(2);
output(5, 210) <= input(3);
output(5, 211) <= input(4);
output(5, 212) <= input(5);
output(5, 213) <= input(6);
output(5, 214) <= input(7);
output(5, 215) <= input(8);
output(5, 216) <= input(9);
output(5, 217) <= input(10);
output(5, 218) <= input(11);
output(5, 219) <= input(12);
output(5, 220) <= input(13);
output(5, 221) <= input(14);
output(5, 222) <= input(15);
output(5, 223) <= input(34);
output(5, 224) <= input(1);
output(5, 225) <= input(2);
output(5, 226) <= input(3);
output(5, 227) <= input(4);
output(5, 228) <= input(5);
output(5, 229) <= input(6);
output(5, 230) <= input(7);
output(5, 231) <= input(8);
output(5, 232) <= input(9);
output(5, 233) <= input(10);
output(5, 234) <= input(11);
output(5, 235) <= input(12);
output(5, 236) <= input(13);
output(5, 237) <= input(14);
output(5, 238) <= input(15);
output(5, 239) <= input(34);
output(5, 240) <= input(18);
output(5, 241) <= input(19);
output(5, 242) <= input(20);
output(5, 243) <= input(21);
output(5, 244) <= input(22);
output(5, 245) <= input(23);
output(5, 246) <= input(24);
output(5, 247) <= input(25);
output(5, 248) <= input(26);
output(5, 249) <= input(27);
output(5, 250) <= input(28);
output(5, 251) <= input(29);
output(5, 252) <= input(30);
output(5, 253) <= input(31);
output(5, 254) <= input(33);
output(5, 255) <= input(35);
output(6, 0) <= input(17);
output(6, 1) <= input(18);
output(6, 2) <= input(19);
output(6, 3) <= input(20);
output(6, 4) <= input(21);
output(6, 5) <= input(22);
output(6, 6) <= input(23);
output(6, 7) <= input(24);
output(6, 8) <= input(25);
output(6, 9) <= input(26);
output(6, 10) <= input(27);
output(6, 11) <= input(28);
output(6, 12) <= input(29);
output(6, 13) <= input(30);
output(6, 14) <= input(31);
output(6, 15) <= input(33);
output(6, 16) <= input(17);
output(6, 17) <= input(18);
output(6, 18) <= input(19);
output(6, 19) <= input(20);
output(6, 20) <= input(21);
output(6, 21) <= input(22);
output(6, 22) <= input(23);
output(6, 23) <= input(24);
output(6, 24) <= input(25);
output(6, 25) <= input(26);
output(6, 26) <= input(27);
output(6, 27) <= input(28);
output(6, 28) <= input(29);
output(6, 29) <= input(30);
output(6, 30) <= input(31);
output(6, 31) <= input(33);
output(6, 32) <= input(17);
output(6, 33) <= input(18);
output(6, 34) <= input(19);
output(6, 35) <= input(20);
output(6, 36) <= input(21);
output(6, 37) <= input(22);
output(6, 38) <= input(23);
output(6, 39) <= input(24);
output(6, 40) <= input(25);
output(6, 41) <= input(26);
output(6, 42) <= input(27);
output(6, 43) <= input(28);
output(6, 44) <= input(29);
output(6, 45) <= input(30);
output(6, 46) <= input(31);
output(6, 47) <= input(33);
output(6, 48) <= input(17);
output(6, 49) <= input(18);
output(6, 50) <= input(19);
output(6, 51) <= input(20);
output(6, 52) <= input(21);
output(6, 53) <= input(22);
output(6, 54) <= input(23);
output(6, 55) <= input(24);
output(6, 56) <= input(25);
output(6, 57) <= input(26);
output(6, 58) <= input(27);
output(6, 59) <= input(28);
output(6, 60) <= input(29);
output(6, 61) <= input(30);
output(6, 62) <= input(31);
output(6, 63) <= input(33);
output(6, 64) <= input(17);
output(6, 65) <= input(18);
output(6, 66) <= input(19);
output(6, 67) <= input(20);
output(6, 68) <= input(21);
output(6, 69) <= input(22);
output(6, 70) <= input(23);
output(6, 71) <= input(24);
output(6, 72) <= input(25);
output(6, 73) <= input(26);
output(6, 74) <= input(27);
output(6, 75) <= input(28);
output(6, 76) <= input(29);
output(6, 77) <= input(30);
output(6, 78) <= input(31);
output(6, 79) <= input(33);
output(6, 80) <= input(1);
output(6, 81) <= input(2);
output(6, 82) <= input(3);
output(6, 83) <= input(4);
output(6, 84) <= input(5);
output(6, 85) <= input(6);
output(6, 86) <= input(7);
output(6, 87) <= input(8);
output(6, 88) <= input(9);
output(6, 89) <= input(10);
output(6, 90) <= input(11);
output(6, 91) <= input(12);
output(6, 92) <= input(13);
output(6, 93) <= input(14);
output(6, 94) <= input(15);
output(6, 95) <= input(34);
output(6, 96) <= input(1);
output(6, 97) <= input(2);
output(6, 98) <= input(3);
output(6, 99) <= input(4);
output(6, 100) <= input(5);
output(6, 101) <= input(6);
output(6, 102) <= input(7);
output(6, 103) <= input(8);
output(6, 104) <= input(9);
output(6, 105) <= input(10);
output(6, 106) <= input(11);
output(6, 107) <= input(12);
output(6, 108) <= input(13);
output(6, 109) <= input(14);
output(6, 110) <= input(15);
output(6, 111) <= input(34);
output(6, 112) <= input(1);
output(6, 113) <= input(2);
output(6, 114) <= input(3);
output(6, 115) <= input(4);
output(6, 116) <= input(5);
output(6, 117) <= input(6);
output(6, 118) <= input(7);
output(6, 119) <= input(8);
output(6, 120) <= input(9);
output(6, 121) <= input(10);
output(6, 122) <= input(11);
output(6, 123) <= input(12);
output(6, 124) <= input(13);
output(6, 125) <= input(14);
output(6, 126) <= input(15);
output(6, 127) <= input(34);
output(6, 128) <= input(1);
output(6, 129) <= input(2);
output(6, 130) <= input(3);
output(6, 131) <= input(4);
output(6, 132) <= input(5);
output(6, 133) <= input(6);
output(6, 134) <= input(7);
output(6, 135) <= input(8);
output(6, 136) <= input(9);
output(6, 137) <= input(10);
output(6, 138) <= input(11);
output(6, 139) <= input(12);
output(6, 140) <= input(13);
output(6, 141) <= input(14);
output(6, 142) <= input(15);
output(6, 143) <= input(34);
output(6, 144) <= input(1);
output(6, 145) <= input(2);
output(6, 146) <= input(3);
output(6, 147) <= input(4);
output(6, 148) <= input(5);
output(6, 149) <= input(6);
output(6, 150) <= input(7);
output(6, 151) <= input(8);
output(6, 152) <= input(9);
output(6, 153) <= input(10);
output(6, 154) <= input(11);
output(6, 155) <= input(12);
output(6, 156) <= input(13);
output(6, 157) <= input(14);
output(6, 158) <= input(15);
output(6, 159) <= input(34);
output(6, 160) <= input(18);
output(6, 161) <= input(19);
output(6, 162) <= input(20);
output(6, 163) <= input(21);
output(6, 164) <= input(22);
output(6, 165) <= input(23);
output(6, 166) <= input(24);
output(6, 167) <= input(25);
output(6, 168) <= input(26);
output(6, 169) <= input(27);
output(6, 170) <= input(28);
output(6, 171) <= input(29);
output(6, 172) <= input(30);
output(6, 173) <= input(31);
output(6, 174) <= input(33);
output(6, 175) <= input(35);
output(6, 176) <= input(18);
output(6, 177) <= input(19);
output(6, 178) <= input(20);
output(6, 179) <= input(21);
output(6, 180) <= input(22);
output(6, 181) <= input(23);
output(6, 182) <= input(24);
output(6, 183) <= input(25);
output(6, 184) <= input(26);
output(6, 185) <= input(27);
output(6, 186) <= input(28);
output(6, 187) <= input(29);
output(6, 188) <= input(30);
output(6, 189) <= input(31);
output(6, 190) <= input(33);
output(6, 191) <= input(35);
output(6, 192) <= input(18);
output(6, 193) <= input(19);
output(6, 194) <= input(20);
output(6, 195) <= input(21);
output(6, 196) <= input(22);
output(6, 197) <= input(23);
output(6, 198) <= input(24);
output(6, 199) <= input(25);
output(6, 200) <= input(26);
output(6, 201) <= input(27);
output(6, 202) <= input(28);
output(6, 203) <= input(29);
output(6, 204) <= input(30);
output(6, 205) <= input(31);
output(6, 206) <= input(33);
output(6, 207) <= input(35);
output(6, 208) <= input(18);
output(6, 209) <= input(19);
output(6, 210) <= input(20);
output(6, 211) <= input(21);
output(6, 212) <= input(22);
output(6, 213) <= input(23);
output(6, 214) <= input(24);
output(6, 215) <= input(25);
output(6, 216) <= input(26);
output(6, 217) <= input(27);
output(6, 218) <= input(28);
output(6, 219) <= input(29);
output(6, 220) <= input(30);
output(6, 221) <= input(31);
output(6, 222) <= input(33);
output(6, 223) <= input(35);
output(6, 224) <= input(18);
output(6, 225) <= input(19);
output(6, 226) <= input(20);
output(6, 227) <= input(21);
output(6, 228) <= input(22);
output(6, 229) <= input(23);
output(6, 230) <= input(24);
output(6, 231) <= input(25);
output(6, 232) <= input(26);
output(6, 233) <= input(27);
output(6, 234) <= input(28);
output(6, 235) <= input(29);
output(6, 236) <= input(30);
output(6, 237) <= input(31);
output(6, 238) <= input(33);
output(6, 239) <= input(35);
output(6, 240) <= input(2);
output(6, 241) <= input(3);
output(6, 242) <= input(4);
output(6, 243) <= input(5);
output(6, 244) <= input(6);
output(6, 245) <= input(7);
output(6, 246) <= input(8);
output(6, 247) <= input(9);
output(6, 248) <= input(10);
output(6, 249) <= input(11);
output(6, 250) <= input(12);
output(6, 251) <= input(13);
output(6, 252) <= input(14);
output(6, 253) <= input(15);
output(6, 254) <= input(34);
output(6, 255) <= input(36);
output(7, 0) <= input(17);
output(7, 1) <= input(18);
output(7, 2) <= input(19);
output(7, 3) <= input(20);
output(7, 4) <= input(21);
output(7, 5) <= input(22);
output(7, 6) <= input(23);
output(7, 7) <= input(24);
output(7, 8) <= input(25);
output(7, 9) <= input(26);
output(7, 10) <= input(27);
output(7, 11) <= input(28);
output(7, 12) <= input(29);
output(7, 13) <= input(30);
output(7, 14) <= input(31);
output(7, 15) <= input(33);
output(7, 16) <= input(17);
output(7, 17) <= input(18);
output(7, 18) <= input(19);
output(7, 19) <= input(20);
output(7, 20) <= input(21);
output(7, 21) <= input(22);
output(7, 22) <= input(23);
output(7, 23) <= input(24);
output(7, 24) <= input(25);
output(7, 25) <= input(26);
output(7, 26) <= input(27);
output(7, 27) <= input(28);
output(7, 28) <= input(29);
output(7, 29) <= input(30);
output(7, 30) <= input(31);
output(7, 31) <= input(33);
output(7, 32) <= input(17);
output(7, 33) <= input(18);
output(7, 34) <= input(19);
output(7, 35) <= input(20);
output(7, 36) <= input(21);
output(7, 37) <= input(22);
output(7, 38) <= input(23);
output(7, 39) <= input(24);
output(7, 40) <= input(25);
output(7, 41) <= input(26);
output(7, 42) <= input(27);
output(7, 43) <= input(28);
output(7, 44) <= input(29);
output(7, 45) <= input(30);
output(7, 46) <= input(31);
output(7, 47) <= input(33);
output(7, 48) <= input(1);
output(7, 49) <= input(2);
output(7, 50) <= input(3);
output(7, 51) <= input(4);
output(7, 52) <= input(5);
output(7, 53) <= input(6);
output(7, 54) <= input(7);
output(7, 55) <= input(8);
output(7, 56) <= input(9);
output(7, 57) <= input(10);
output(7, 58) <= input(11);
output(7, 59) <= input(12);
output(7, 60) <= input(13);
output(7, 61) <= input(14);
output(7, 62) <= input(15);
output(7, 63) <= input(34);
output(7, 64) <= input(1);
output(7, 65) <= input(2);
output(7, 66) <= input(3);
output(7, 67) <= input(4);
output(7, 68) <= input(5);
output(7, 69) <= input(6);
output(7, 70) <= input(7);
output(7, 71) <= input(8);
output(7, 72) <= input(9);
output(7, 73) <= input(10);
output(7, 74) <= input(11);
output(7, 75) <= input(12);
output(7, 76) <= input(13);
output(7, 77) <= input(14);
output(7, 78) <= input(15);
output(7, 79) <= input(34);
output(7, 80) <= input(1);
output(7, 81) <= input(2);
output(7, 82) <= input(3);
output(7, 83) <= input(4);
output(7, 84) <= input(5);
output(7, 85) <= input(6);
output(7, 86) <= input(7);
output(7, 87) <= input(8);
output(7, 88) <= input(9);
output(7, 89) <= input(10);
output(7, 90) <= input(11);
output(7, 91) <= input(12);
output(7, 92) <= input(13);
output(7, 93) <= input(14);
output(7, 94) <= input(15);
output(7, 95) <= input(34);
output(7, 96) <= input(1);
output(7, 97) <= input(2);
output(7, 98) <= input(3);
output(7, 99) <= input(4);
output(7, 100) <= input(5);
output(7, 101) <= input(6);
output(7, 102) <= input(7);
output(7, 103) <= input(8);
output(7, 104) <= input(9);
output(7, 105) <= input(10);
output(7, 106) <= input(11);
output(7, 107) <= input(12);
output(7, 108) <= input(13);
output(7, 109) <= input(14);
output(7, 110) <= input(15);
output(7, 111) <= input(34);
output(7, 112) <= input(18);
output(7, 113) <= input(19);
output(7, 114) <= input(20);
output(7, 115) <= input(21);
output(7, 116) <= input(22);
output(7, 117) <= input(23);
output(7, 118) <= input(24);
output(7, 119) <= input(25);
output(7, 120) <= input(26);
output(7, 121) <= input(27);
output(7, 122) <= input(28);
output(7, 123) <= input(29);
output(7, 124) <= input(30);
output(7, 125) <= input(31);
output(7, 126) <= input(33);
output(7, 127) <= input(35);
output(7, 128) <= input(18);
output(7, 129) <= input(19);
output(7, 130) <= input(20);
output(7, 131) <= input(21);
output(7, 132) <= input(22);
output(7, 133) <= input(23);
output(7, 134) <= input(24);
output(7, 135) <= input(25);
output(7, 136) <= input(26);
output(7, 137) <= input(27);
output(7, 138) <= input(28);
output(7, 139) <= input(29);
output(7, 140) <= input(30);
output(7, 141) <= input(31);
output(7, 142) <= input(33);
output(7, 143) <= input(35);
output(7, 144) <= input(18);
output(7, 145) <= input(19);
output(7, 146) <= input(20);
output(7, 147) <= input(21);
output(7, 148) <= input(22);
output(7, 149) <= input(23);
output(7, 150) <= input(24);
output(7, 151) <= input(25);
output(7, 152) <= input(26);
output(7, 153) <= input(27);
output(7, 154) <= input(28);
output(7, 155) <= input(29);
output(7, 156) <= input(30);
output(7, 157) <= input(31);
output(7, 158) <= input(33);
output(7, 159) <= input(35);
output(7, 160) <= input(18);
output(7, 161) <= input(19);
output(7, 162) <= input(20);
output(7, 163) <= input(21);
output(7, 164) <= input(22);
output(7, 165) <= input(23);
output(7, 166) <= input(24);
output(7, 167) <= input(25);
output(7, 168) <= input(26);
output(7, 169) <= input(27);
output(7, 170) <= input(28);
output(7, 171) <= input(29);
output(7, 172) <= input(30);
output(7, 173) <= input(31);
output(7, 174) <= input(33);
output(7, 175) <= input(35);
output(7, 176) <= input(2);
output(7, 177) <= input(3);
output(7, 178) <= input(4);
output(7, 179) <= input(5);
output(7, 180) <= input(6);
output(7, 181) <= input(7);
output(7, 182) <= input(8);
output(7, 183) <= input(9);
output(7, 184) <= input(10);
output(7, 185) <= input(11);
output(7, 186) <= input(12);
output(7, 187) <= input(13);
output(7, 188) <= input(14);
output(7, 189) <= input(15);
output(7, 190) <= input(34);
output(7, 191) <= input(36);
output(7, 192) <= input(2);
output(7, 193) <= input(3);
output(7, 194) <= input(4);
output(7, 195) <= input(5);
output(7, 196) <= input(6);
output(7, 197) <= input(7);
output(7, 198) <= input(8);
output(7, 199) <= input(9);
output(7, 200) <= input(10);
output(7, 201) <= input(11);
output(7, 202) <= input(12);
output(7, 203) <= input(13);
output(7, 204) <= input(14);
output(7, 205) <= input(15);
output(7, 206) <= input(34);
output(7, 207) <= input(36);
output(7, 208) <= input(2);
output(7, 209) <= input(3);
output(7, 210) <= input(4);
output(7, 211) <= input(5);
output(7, 212) <= input(6);
output(7, 213) <= input(7);
output(7, 214) <= input(8);
output(7, 215) <= input(9);
output(7, 216) <= input(10);
output(7, 217) <= input(11);
output(7, 218) <= input(12);
output(7, 219) <= input(13);
output(7, 220) <= input(14);
output(7, 221) <= input(15);
output(7, 222) <= input(34);
output(7, 223) <= input(36);
output(7, 224) <= input(2);
output(7, 225) <= input(3);
output(7, 226) <= input(4);
output(7, 227) <= input(5);
output(7, 228) <= input(6);
output(7, 229) <= input(7);
output(7, 230) <= input(8);
output(7, 231) <= input(9);
output(7, 232) <= input(10);
output(7, 233) <= input(11);
output(7, 234) <= input(12);
output(7, 235) <= input(13);
output(7, 236) <= input(14);
output(7, 237) <= input(15);
output(7, 238) <= input(34);
output(7, 239) <= input(36);
output(7, 240) <= input(19);
output(7, 241) <= input(20);
output(7, 242) <= input(21);
output(7, 243) <= input(22);
output(7, 244) <= input(23);
output(7, 245) <= input(24);
output(7, 246) <= input(25);
output(7, 247) <= input(26);
output(7, 248) <= input(27);
output(7, 249) <= input(28);
output(7, 250) <= input(29);
output(7, 251) <= input(30);
output(7, 252) <= input(31);
output(7, 253) <= input(33);
output(7, 254) <= input(35);
output(7, 255) <= input(37);
when "1110" =>
output(0, 0) <= input(0);
output(0, 1) <= input(1);
output(0, 2) <= input(2);
output(0, 3) <= input(3);
output(0, 4) <= input(4);
output(0, 5) <= input(5);
output(0, 6) <= input(6);
output(0, 7) <= input(7);
output(0, 8) <= input(8);
output(0, 9) <= input(9);
output(0, 10) <= input(10);
output(0, 11) <= input(11);
output(0, 12) <= input(12);
output(0, 13) <= input(13);
output(0, 14) <= input(14);
output(0, 15) <= input(15);
output(0, 16) <= input(0);
output(0, 17) <= input(1);
output(0, 18) <= input(2);
output(0, 19) <= input(3);
output(0, 20) <= input(4);
output(0, 21) <= input(5);
output(0, 22) <= input(6);
output(0, 23) <= input(7);
output(0, 24) <= input(8);
output(0, 25) <= input(9);
output(0, 26) <= input(10);
output(0, 27) <= input(11);
output(0, 28) <= input(12);
output(0, 29) <= input(13);
output(0, 30) <= input(14);
output(0, 31) <= input(15);
output(0, 32) <= input(16);
output(0, 33) <= input(17);
output(0, 34) <= input(18);
output(0, 35) <= input(19);
output(0, 36) <= input(20);
output(0, 37) <= input(21);
output(0, 38) <= input(22);
output(0, 39) <= input(23);
output(0, 40) <= input(24);
output(0, 41) <= input(25);
output(0, 42) <= input(26);
output(0, 43) <= input(27);
output(0, 44) <= input(28);
output(0, 45) <= input(29);
output(0, 46) <= input(30);
output(0, 47) <= input(31);
output(0, 48) <= input(16);
output(0, 49) <= input(17);
output(0, 50) <= input(18);
output(0, 51) <= input(19);
output(0, 52) <= input(20);
output(0, 53) <= input(21);
output(0, 54) <= input(22);
output(0, 55) <= input(23);
output(0, 56) <= input(24);
output(0, 57) <= input(25);
output(0, 58) <= input(26);
output(0, 59) <= input(27);
output(0, 60) <= input(28);
output(0, 61) <= input(29);
output(0, 62) <= input(30);
output(0, 63) <= input(31);
output(0, 64) <= input(16);
output(0, 65) <= input(17);
output(0, 66) <= input(18);
output(0, 67) <= input(19);
output(0, 68) <= input(20);
output(0, 69) <= input(21);
output(0, 70) <= input(22);
output(0, 71) <= input(23);
output(0, 72) <= input(24);
output(0, 73) <= input(25);
output(0, 74) <= input(26);
output(0, 75) <= input(27);
output(0, 76) <= input(28);
output(0, 77) <= input(29);
output(0, 78) <= input(30);
output(0, 79) <= input(31);
output(0, 80) <= input(1);
output(0, 81) <= input(2);
output(0, 82) <= input(3);
output(0, 83) <= input(4);
output(0, 84) <= input(5);
output(0, 85) <= input(6);
output(0, 86) <= input(7);
output(0, 87) <= input(8);
output(0, 88) <= input(9);
output(0, 89) <= input(10);
output(0, 90) <= input(11);
output(0, 91) <= input(12);
output(0, 92) <= input(13);
output(0, 93) <= input(14);
output(0, 94) <= input(15);
output(0, 95) <= input(32);
output(0, 96) <= input(1);
output(0, 97) <= input(2);
output(0, 98) <= input(3);
output(0, 99) <= input(4);
output(0, 100) <= input(5);
output(0, 101) <= input(6);
output(0, 102) <= input(7);
output(0, 103) <= input(8);
output(0, 104) <= input(9);
output(0, 105) <= input(10);
output(0, 106) <= input(11);
output(0, 107) <= input(12);
output(0, 108) <= input(13);
output(0, 109) <= input(14);
output(0, 110) <= input(15);
output(0, 111) <= input(32);
output(0, 112) <= input(17);
output(0, 113) <= input(18);
output(0, 114) <= input(19);
output(0, 115) <= input(20);
output(0, 116) <= input(21);
output(0, 117) <= input(22);
output(0, 118) <= input(23);
output(0, 119) <= input(24);
output(0, 120) <= input(25);
output(0, 121) <= input(26);
output(0, 122) <= input(27);
output(0, 123) <= input(28);
output(0, 124) <= input(29);
output(0, 125) <= input(30);
output(0, 126) <= input(31);
output(0, 127) <= input(33);
output(0, 128) <= input(17);
output(0, 129) <= input(18);
output(0, 130) <= input(19);
output(0, 131) <= input(20);
output(0, 132) <= input(21);
output(0, 133) <= input(22);
output(0, 134) <= input(23);
output(0, 135) <= input(24);
output(0, 136) <= input(25);
output(0, 137) <= input(26);
output(0, 138) <= input(27);
output(0, 139) <= input(28);
output(0, 140) <= input(29);
output(0, 141) <= input(30);
output(0, 142) <= input(31);
output(0, 143) <= input(33);
output(0, 144) <= input(17);
output(0, 145) <= input(18);
output(0, 146) <= input(19);
output(0, 147) <= input(20);
output(0, 148) <= input(21);
output(0, 149) <= input(22);
output(0, 150) <= input(23);
output(0, 151) <= input(24);
output(0, 152) <= input(25);
output(0, 153) <= input(26);
output(0, 154) <= input(27);
output(0, 155) <= input(28);
output(0, 156) <= input(29);
output(0, 157) <= input(30);
output(0, 158) <= input(31);
output(0, 159) <= input(33);
output(0, 160) <= input(2);
output(0, 161) <= input(3);
output(0, 162) <= input(4);
output(0, 163) <= input(5);
output(0, 164) <= input(6);
output(0, 165) <= input(7);
output(0, 166) <= input(8);
output(0, 167) <= input(9);
output(0, 168) <= input(10);
output(0, 169) <= input(11);
output(0, 170) <= input(12);
output(0, 171) <= input(13);
output(0, 172) <= input(14);
output(0, 173) <= input(15);
output(0, 174) <= input(32);
output(0, 175) <= input(34);
output(0, 176) <= input(2);
output(0, 177) <= input(3);
output(0, 178) <= input(4);
output(0, 179) <= input(5);
output(0, 180) <= input(6);
output(0, 181) <= input(7);
output(0, 182) <= input(8);
output(0, 183) <= input(9);
output(0, 184) <= input(10);
output(0, 185) <= input(11);
output(0, 186) <= input(12);
output(0, 187) <= input(13);
output(0, 188) <= input(14);
output(0, 189) <= input(15);
output(0, 190) <= input(32);
output(0, 191) <= input(34);
output(0, 192) <= input(2);
output(0, 193) <= input(3);
output(0, 194) <= input(4);
output(0, 195) <= input(5);
output(0, 196) <= input(6);
output(0, 197) <= input(7);
output(0, 198) <= input(8);
output(0, 199) <= input(9);
output(0, 200) <= input(10);
output(0, 201) <= input(11);
output(0, 202) <= input(12);
output(0, 203) <= input(13);
output(0, 204) <= input(14);
output(0, 205) <= input(15);
output(0, 206) <= input(32);
output(0, 207) <= input(34);
output(0, 208) <= input(18);
output(0, 209) <= input(19);
output(0, 210) <= input(20);
output(0, 211) <= input(21);
output(0, 212) <= input(22);
output(0, 213) <= input(23);
output(0, 214) <= input(24);
output(0, 215) <= input(25);
output(0, 216) <= input(26);
output(0, 217) <= input(27);
output(0, 218) <= input(28);
output(0, 219) <= input(29);
output(0, 220) <= input(30);
output(0, 221) <= input(31);
output(0, 222) <= input(33);
output(0, 223) <= input(35);
output(0, 224) <= input(18);
output(0, 225) <= input(19);
output(0, 226) <= input(20);
output(0, 227) <= input(21);
output(0, 228) <= input(22);
output(0, 229) <= input(23);
output(0, 230) <= input(24);
output(0, 231) <= input(25);
output(0, 232) <= input(26);
output(0, 233) <= input(27);
output(0, 234) <= input(28);
output(0, 235) <= input(29);
output(0, 236) <= input(30);
output(0, 237) <= input(31);
output(0, 238) <= input(33);
output(0, 239) <= input(35);
output(0, 240) <= input(3);
output(0, 241) <= input(4);
output(0, 242) <= input(5);
output(0, 243) <= input(6);
output(0, 244) <= input(7);
output(0, 245) <= input(8);
output(0, 246) <= input(9);
output(0, 247) <= input(10);
output(0, 248) <= input(11);
output(0, 249) <= input(12);
output(0, 250) <= input(13);
output(0, 251) <= input(14);
output(0, 252) <= input(15);
output(0, 253) <= input(32);
output(0, 254) <= input(34);
output(0, 255) <= input(36);
output(1, 0) <= input(0);
output(1, 1) <= input(1);
output(1, 2) <= input(2);
output(1, 3) <= input(3);
output(1, 4) <= input(4);
output(1, 5) <= input(5);
output(1, 6) <= input(6);
output(1, 7) <= input(7);
output(1, 8) <= input(8);
output(1, 9) <= input(9);
output(1, 10) <= input(10);
output(1, 11) <= input(11);
output(1, 12) <= input(12);
output(1, 13) <= input(13);
output(1, 14) <= input(14);
output(1, 15) <= input(15);
output(1, 16) <= input(16);
output(1, 17) <= input(17);
output(1, 18) <= input(18);
output(1, 19) <= input(19);
output(1, 20) <= input(20);
output(1, 21) <= input(21);
output(1, 22) <= input(22);
output(1, 23) <= input(23);
output(1, 24) <= input(24);
output(1, 25) <= input(25);
output(1, 26) <= input(26);
output(1, 27) <= input(27);
output(1, 28) <= input(28);
output(1, 29) <= input(29);
output(1, 30) <= input(30);
output(1, 31) <= input(31);
output(1, 32) <= input(16);
output(1, 33) <= input(17);
output(1, 34) <= input(18);
output(1, 35) <= input(19);
output(1, 36) <= input(20);
output(1, 37) <= input(21);
output(1, 38) <= input(22);
output(1, 39) <= input(23);
output(1, 40) <= input(24);
output(1, 41) <= input(25);
output(1, 42) <= input(26);
output(1, 43) <= input(27);
output(1, 44) <= input(28);
output(1, 45) <= input(29);
output(1, 46) <= input(30);
output(1, 47) <= input(31);
output(1, 48) <= input(1);
output(1, 49) <= input(2);
output(1, 50) <= input(3);
output(1, 51) <= input(4);
output(1, 52) <= input(5);
output(1, 53) <= input(6);
output(1, 54) <= input(7);
output(1, 55) <= input(8);
output(1, 56) <= input(9);
output(1, 57) <= input(10);
output(1, 58) <= input(11);
output(1, 59) <= input(12);
output(1, 60) <= input(13);
output(1, 61) <= input(14);
output(1, 62) <= input(15);
output(1, 63) <= input(32);
output(1, 64) <= input(1);
output(1, 65) <= input(2);
output(1, 66) <= input(3);
output(1, 67) <= input(4);
output(1, 68) <= input(5);
output(1, 69) <= input(6);
output(1, 70) <= input(7);
output(1, 71) <= input(8);
output(1, 72) <= input(9);
output(1, 73) <= input(10);
output(1, 74) <= input(11);
output(1, 75) <= input(12);
output(1, 76) <= input(13);
output(1, 77) <= input(14);
output(1, 78) <= input(15);
output(1, 79) <= input(32);
output(1, 80) <= input(17);
output(1, 81) <= input(18);
output(1, 82) <= input(19);
output(1, 83) <= input(20);
output(1, 84) <= input(21);
output(1, 85) <= input(22);
output(1, 86) <= input(23);
output(1, 87) <= input(24);
output(1, 88) <= input(25);
output(1, 89) <= input(26);
output(1, 90) <= input(27);
output(1, 91) <= input(28);
output(1, 92) <= input(29);
output(1, 93) <= input(30);
output(1, 94) <= input(31);
output(1, 95) <= input(33);
output(1, 96) <= input(17);
output(1, 97) <= input(18);
output(1, 98) <= input(19);
output(1, 99) <= input(20);
output(1, 100) <= input(21);
output(1, 101) <= input(22);
output(1, 102) <= input(23);
output(1, 103) <= input(24);
output(1, 104) <= input(25);
output(1, 105) <= input(26);
output(1, 106) <= input(27);
output(1, 107) <= input(28);
output(1, 108) <= input(29);
output(1, 109) <= input(30);
output(1, 110) <= input(31);
output(1, 111) <= input(33);
output(1, 112) <= input(2);
output(1, 113) <= input(3);
output(1, 114) <= input(4);
output(1, 115) <= input(5);
output(1, 116) <= input(6);
output(1, 117) <= input(7);
output(1, 118) <= input(8);
output(1, 119) <= input(9);
output(1, 120) <= input(10);
output(1, 121) <= input(11);
output(1, 122) <= input(12);
output(1, 123) <= input(13);
output(1, 124) <= input(14);
output(1, 125) <= input(15);
output(1, 126) <= input(32);
output(1, 127) <= input(34);
output(1, 128) <= input(2);
output(1, 129) <= input(3);
output(1, 130) <= input(4);
output(1, 131) <= input(5);
output(1, 132) <= input(6);
output(1, 133) <= input(7);
output(1, 134) <= input(8);
output(1, 135) <= input(9);
output(1, 136) <= input(10);
output(1, 137) <= input(11);
output(1, 138) <= input(12);
output(1, 139) <= input(13);
output(1, 140) <= input(14);
output(1, 141) <= input(15);
output(1, 142) <= input(32);
output(1, 143) <= input(34);
output(1, 144) <= input(18);
output(1, 145) <= input(19);
output(1, 146) <= input(20);
output(1, 147) <= input(21);
output(1, 148) <= input(22);
output(1, 149) <= input(23);
output(1, 150) <= input(24);
output(1, 151) <= input(25);
output(1, 152) <= input(26);
output(1, 153) <= input(27);
output(1, 154) <= input(28);
output(1, 155) <= input(29);
output(1, 156) <= input(30);
output(1, 157) <= input(31);
output(1, 158) <= input(33);
output(1, 159) <= input(35);
output(1, 160) <= input(18);
output(1, 161) <= input(19);
output(1, 162) <= input(20);
output(1, 163) <= input(21);
output(1, 164) <= input(22);
output(1, 165) <= input(23);
output(1, 166) <= input(24);
output(1, 167) <= input(25);
output(1, 168) <= input(26);
output(1, 169) <= input(27);
output(1, 170) <= input(28);
output(1, 171) <= input(29);
output(1, 172) <= input(30);
output(1, 173) <= input(31);
output(1, 174) <= input(33);
output(1, 175) <= input(35);
output(1, 176) <= input(3);
output(1, 177) <= input(4);
output(1, 178) <= input(5);
output(1, 179) <= input(6);
output(1, 180) <= input(7);
output(1, 181) <= input(8);
output(1, 182) <= input(9);
output(1, 183) <= input(10);
output(1, 184) <= input(11);
output(1, 185) <= input(12);
output(1, 186) <= input(13);
output(1, 187) <= input(14);
output(1, 188) <= input(15);
output(1, 189) <= input(32);
output(1, 190) <= input(34);
output(1, 191) <= input(36);
output(1, 192) <= input(3);
output(1, 193) <= input(4);
output(1, 194) <= input(5);
output(1, 195) <= input(6);
output(1, 196) <= input(7);
output(1, 197) <= input(8);
output(1, 198) <= input(9);
output(1, 199) <= input(10);
output(1, 200) <= input(11);
output(1, 201) <= input(12);
output(1, 202) <= input(13);
output(1, 203) <= input(14);
output(1, 204) <= input(15);
output(1, 205) <= input(32);
output(1, 206) <= input(34);
output(1, 207) <= input(36);
output(1, 208) <= input(19);
output(1, 209) <= input(20);
output(1, 210) <= input(21);
output(1, 211) <= input(22);
output(1, 212) <= input(23);
output(1, 213) <= input(24);
output(1, 214) <= input(25);
output(1, 215) <= input(26);
output(1, 216) <= input(27);
output(1, 217) <= input(28);
output(1, 218) <= input(29);
output(1, 219) <= input(30);
output(1, 220) <= input(31);
output(1, 221) <= input(33);
output(1, 222) <= input(35);
output(1, 223) <= input(37);
output(1, 224) <= input(19);
output(1, 225) <= input(20);
output(1, 226) <= input(21);
output(1, 227) <= input(22);
output(1, 228) <= input(23);
output(1, 229) <= input(24);
output(1, 230) <= input(25);
output(1, 231) <= input(26);
output(1, 232) <= input(27);
output(1, 233) <= input(28);
output(1, 234) <= input(29);
output(1, 235) <= input(30);
output(1, 236) <= input(31);
output(1, 237) <= input(33);
output(1, 238) <= input(35);
output(1, 239) <= input(37);
output(1, 240) <= input(4);
output(1, 241) <= input(5);
output(1, 242) <= input(6);
output(1, 243) <= input(7);
output(1, 244) <= input(8);
output(1, 245) <= input(9);
output(1, 246) <= input(10);
output(1, 247) <= input(11);
output(1, 248) <= input(12);
output(1, 249) <= input(13);
output(1, 250) <= input(14);
output(1, 251) <= input(15);
output(1, 252) <= input(32);
output(1, 253) <= input(34);
output(1, 254) <= input(36);
output(1, 255) <= input(38);
output(2, 0) <= input(0);
output(2, 1) <= input(1);
output(2, 2) <= input(2);
output(2, 3) <= input(3);
output(2, 4) <= input(4);
output(2, 5) <= input(5);
output(2, 6) <= input(6);
output(2, 7) <= input(7);
output(2, 8) <= input(8);
output(2, 9) <= input(9);
output(2, 10) <= input(10);
output(2, 11) <= input(11);
output(2, 12) <= input(12);
output(2, 13) <= input(13);
output(2, 14) <= input(14);
output(2, 15) <= input(15);
output(2, 16) <= input(16);
output(2, 17) <= input(17);
output(2, 18) <= input(18);
output(2, 19) <= input(19);
output(2, 20) <= input(20);
output(2, 21) <= input(21);
output(2, 22) <= input(22);
output(2, 23) <= input(23);
output(2, 24) <= input(24);
output(2, 25) <= input(25);
output(2, 26) <= input(26);
output(2, 27) <= input(27);
output(2, 28) <= input(28);
output(2, 29) <= input(29);
output(2, 30) <= input(30);
output(2, 31) <= input(31);
output(2, 32) <= input(16);
output(2, 33) <= input(17);
output(2, 34) <= input(18);
output(2, 35) <= input(19);
output(2, 36) <= input(20);
output(2, 37) <= input(21);
output(2, 38) <= input(22);
output(2, 39) <= input(23);
output(2, 40) <= input(24);
output(2, 41) <= input(25);
output(2, 42) <= input(26);
output(2, 43) <= input(27);
output(2, 44) <= input(28);
output(2, 45) <= input(29);
output(2, 46) <= input(30);
output(2, 47) <= input(31);
output(2, 48) <= input(1);
output(2, 49) <= input(2);
output(2, 50) <= input(3);
output(2, 51) <= input(4);
output(2, 52) <= input(5);
output(2, 53) <= input(6);
output(2, 54) <= input(7);
output(2, 55) <= input(8);
output(2, 56) <= input(9);
output(2, 57) <= input(10);
output(2, 58) <= input(11);
output(2, 59) <= input(12);
output(2, 60) <= input(13);
output(2, 61) <= input(14);
output(2, 62) <= input(15);
output(2, 63) <= input(32);
output(2, 64) <= input(17);
output(2, 65) <= input(18);
output(2, 66) <= input(19);
output(2, 67) <= input(20);
output(2, 68) <= input(21);
output(2, 69) <= input(22);
output(2, 70) <= input(23);
output(2, 71) <= input(24);
output(2, 72) <= input(25);
output(2, 73) <= input(26);
output(2, 74) <= input(27);
output(2, 75) <= input(28);
output(2, 76) <= input(29);
output(2, 77) <= input(30);
output(2, 78) <= input(31);
output(2, 79) <= input(33);
output(2, 80) <= input(17);
output(2, 81) <= input(18);
output(2, 82) <= input(19);
output(2, 83) <= input(20);
output(2, 84) <= input(21);
output(2, 85) <= input(22);
output(2, 86) <= input(23);
output(2, 87) <= input(24);
output(2, 88) <= input(25);
output(2, 89) <= input(26);
output(2, 90) <= input(27);
output(2, 91) <= input(28);
output(2, 92) <= input(29);
output(2, 93) <= input(30);
output(2, 94) <= input(31);
output(2, 95) <= input(33);
output(2, 96) <= input(2);
output(2, 97) <= input(3);
output(2, 98) <= input(4);
output(2, 99) <= input(5);
output(2, 100) <= input(6);
output(2, 101) <= input(7);
output(2, 102) <= input(8);
output(2, 103) <= input(9);
output(2, 104) <= input(10);
output(2, 105) <= input(11);
output(2, 106) <= input(12);
output(2, 107) <= input(13);
output(2, 108) <= input(14);
output(2, 109) <= input(15);
output(2, 110) <= input(32);
output(2, 111) <= input(34);
output(2, 112) <= input(18);
output(2, 113) <= input(19);
output(2, 114) <= input(20);
output(2, 115) <= input(21);
output(2, 116) <= input(22);
output(2, 117) <= input(23);
output(2, 118) <= input(24);
output(2, 119) <= input(25);
output(2, 120) <= input(26);
output(2, 121) <= input(27);
output(2, 122) <= input(28);
output(2, 123) <= input(29);
output(2, 124) <= input(30);
output(2, 125) <= input(31);
output(2, 126) <= input(33);
output(2, 127) <= input(35);
output(2, 128) <= input(18);
output(2, 129) <= input(19);
output(2, 130) <= input(20);
output(2, 131) <= input(21);
output(2, 132) <= input(22);
output(2, 133) <= input(23);
output(2, 134) <= input(24);
output(2, 135) <= input(25);
output(2, 136) <= input(26);
output(2, 137) <= input(27);
output(2, 138) <= input(28);
output(2, 139) <= input(29);
output(2, 140) <= input(30);
output(2, 141) <= input(31);
output(2, 142) <= input(33);
output(2, 143) <= input(35);
output(2, 144) <= input(3);
output(2, 145) <= input(4);
output(2, 146) <= input(5);
output(2, 147) <= input(6);
output(2, 148) <= input(7);
output(2, 149) <= input(8);
output(2, 150) <= input(9);
output(2, 151) <= input(10);
output(2, 152) <= input(11);
output(2, 153) <= input(12);
output(2, 154) <= input(13);
output(2, 155) <= input(14);
output(2, 156) <= input(15);
output(2, 157) <= input(32);
output(2, 158) <= input(34);
output(2, 159) <= input(36);
output(2, 160) <= input(3);
output(2, 161) <= input(4);
output(2, 162) <= input(5);
output(2, 163) <= input(6);
output(2, 164) <= input(7);
output(2, 165) <= input(8);
output(2, 166) <= input(9);
output(2, 167) <= input(10);
output(2, 168) <= input(11);
output(2, 169) <= input(12);
output(2, 170) <= input(13);
output(2, 171) <= input(14);
output(2, 172) <= input(15);
output(2, 173) <= input(32);
output(2, 174) <= input(34);
output(2, 175) <= input(36);
output(2, 176) <= input(19);
output(2, 177) <= input(20);
output(2, 178) <= input(21);
output(2, 179) <= input(22);
output(2, 180) <= input(23);
output(2, 181) <= input(24);
output(2, 182) <= input(25);
output(2, 183) <= input(26);
output(2, 184) <= input(27);
output(2, 185) <= input(28);
output(2, 186) <= input(29);
output(2, 187) <= input(30);
output(2, 188) <= input(31);
output(2, 189) <= input(33);
output(2, 190) <= input(35);
output(2, 191) <= input(37);
output(2, 192) <= input(4);
output(2, 193) <= input(5);
output(2, 194) <= input(6);
output(2, 195) <= input(7);
output(2, 196) <= input(8);
output(2, 197) <= input(9);
output(2, 198) <= input(10);
output(2, 199) <= input(11);
output(2, 200) <= input(12);
output(2, 201) <= input(13);
output(2, 202) <= input(14);
output(2, 203) <= input(15);
output(2, 204) <= input(32);
output(2, 205) <= input(34);
output(2, 206) <= input(36);
output(2, 207) <= input(38);
output(2, 208) <= input(4);
output(2, 209) <= input(5);
output(2, 210) <= input(6);
output(2, 211) <= input(7);
output(2, 212) <= input(8);
output(2, 213) <= input(9);
output(2, 214) <= input(10);
output(2, 215) <= input(11);
output(2, 216) <= input(12);
output(2, 217) <= input(13);
output(2, 218) <= input(14);
output(2, 219) <= input(15);
output(2, 220) <= input(32);
output(2, 221) <= input(34);
output(2, 222) <= input(36);
output(2, 223) <= input(38);
output(2, 224) <= input(20);
output(2, 225) <= input(21);
output(2, 226) <= input(22);
output(2, 227) <= input(23);
output(2, 228) <= input(24);
output(2, 229) <= input(25);
output(2, 230) <= input(26);
output(2, 231) <= input(27);
output(2, 232) <= input(28);
output(2, 233) <= input(29);
output(2, 234) <= input(30);
output(2, 235) <= input(31);
output(2, 236) <= input(33);
output(2, 237) <= input(35);
output(2, 238) <= input(37);
output(2, 239) <= input(39);
output(2, 240) <= input(5);
output(2, 241) <= input(6);
output(2, 242) <= input(7);
output(2, 243) <= input(8);
output(2, 244) <= input(9);
output(2, 245) <= input(10);
output(2, 246) <= input(11);
output(2, 247) <= input(12);
output(2, 248) <= input(13);
output(2, 249) <= input(14);
output(2, 250) <= input(15);
output(2, 251) <= input(32);
output(2, 252) <= input(34);
output(2, 253) <= input(36);
output(2, 254) <= input(38);
output(2, 255) <= input(40);
output(3, 0) <= input(0);
output(3, 1) <= input(1);
output(3, 2) <= input(2);
output(3, 3) <= input(3);
output(3, 4) <= input(4);
output(3, 5) <= input(5);
output(3, 6) <= input(6);
output(3, 7) <= input(7);
output(3, 8) <= input(8);
output(3, 9) <= input(9);
output(3, 10) <= input(10);
output(3, 11) <= input(11);
output(3, 12) <= input(12);
output(3, 13) <= input(13);
output(3, 14) <= input(14);
output(3, 15) <= input(15);
output(3, 16) <= input(16);
output(3, 17) <= input(17);
output(3, 18) <= input(18);
output(3, 19) <= input(19);
output(3, 20) <= input(20);
output(3, 21) <= input(21);
output(3, 22) <= input(22);
output(3, 23) <= input(23);
output(3, 24) <= input(24);
output(3, 25) <= input(25);
output(3, 26) <= input(26);
output(3, 27) <= input(27);
output(3, 28) <= input(28);
output(3, 29) <= input(29);
output(3, 30) <= input(30);
output(3, 31) <= input(31);
output(3, 32) <= input(1);
output(3, 33) <= input(2);
output(3, 34) <= input(3);
output(3, 35) <= input(4);
output(3, 36) <= input(5);
output(3, 37) <= input(6);
output(3, 38) <= input(7);
output(3, 39) <= input(8);
output(3, 40) <= input(9);
output(3, 41) <= input(10);
output(3, 42) <= input(11);
output(3, 43) <= input(12);
output(3, 44) <= input(13);
output(3, 45) <= input(14);
output(3, 46) <= input(15);
output(3, 47) <= input(32);
output(3, 48) <= input(17);
output(3, 49) <= input(18);
output(3, 50) <= input(19);
output(3, 51) <= input(20);
output(3, 52) <= input(21);
output(3, 53) <= input(22);
output(3, 54) <= input(23);
output(3, 55) <= input(24);
output(3, 56) <= input(25);
output(3, 57) <= input(26);
output(3, 58) <= input(27);
output(3, 59) <= input(28);
output(3, 60) <= input(29);
output(3, 61) <= input(30);
output(3, 62) <= input(31);
output(3, 63) <= input(33);
output(3, 64) <= input(17);
output(3, 65) <= input(18);
output(3, 66) <= input(19);
output(3, 67) <= input(20);
output(3, 68) <= input(21);
output(3, 69) <= input(22);
output(3, 70) <= input(23);
output(3, 71) <= input(24);
output(3, 72) <= input(25);
output(3, 73) <= input(26);
output(3, 74) <= input(27);
output(3, 75) <= input(28);
output(3, 76) <= input(29);
output(3, 77) <= input(30);
output(3, 78) <= input(31);
output(3, 79) <= input(33);
output(3, 80) <= input(2);
output(3, 81) <= input(3);
output(3, 82) <= input(4);
output(3, 83) <= input(5);
output(3, 84) <= input(6);
output(3, 85) <= input(7);
output(3, 86) <= input(8);
output(3, 87) <= input(9);
output(3, 88) <= input(10);
output(3, 89) <= input(11);
output(3, 90) <= input(12);
output(3, 91) <= input(13);
output(3, 92) <= input(14);
output(3, 93) <= input(15);
output(3, 94) <= input(32);
output(3, 95) <= input(34);
output(3, 96) <= input(18);
output(3, 97) <= input(19);
output(3, 98) <= input(20);
output(3, 99) <= input(21);
output(3, 100) <= input(22);
output(3, 101) <= input(23);
output(3, 102) <= input(24);
output(3, 103) <= input(25);
output(3, 104) <= input(26);
output(3, 105) <= input(27);
output(3, 106) <= input(28);
output(3, 107) <= input(29);
output(3, 108) <= input(30);
output(3, 109) <= input(31);
output(3, 110) <= input(33);
output(3, 111) <= input(35);
output(3, 112) <= input(3);
output(3, 113) <= input(4);
output(3, 114) <= input(5);
output(3, 115) <= input(6);
output(3, 116) <= input(7);
output(3, 117) <= input(8);
output(3, 118) <= input(9);
output(3, 119) <= input(10);
output(3, 120) <= input(11);
output(3, 121) <= input(12);
output(3, 122) <= input(13);
output(3, 123) <= input(14);
output(3, 124) <= input(15);
output(3, 125) <= input(32);
output(3, 126) <= input(34);
output(3, 127) <= input(36);
output(3, 128) <= input(3);
output(3, 129) <= input(4);
output(3, 130) <= input(5);
output(3, 131) <= input(6);
output(3, 132) <= input(7);
output(3, 133) <= input(8);
output(3, 134) <= input(9);
output(3, 135) <= input(10);
output(3, 136) <= input(11);
output(3, 137) <= input(12);
output(3, 138) <= input(13);
output(3, 139) <= input(14);
output(3, 140) <= input(15);
output(3, 141) <= input(32);
output(3, 142) <= input(34);
output(3, 143) <= input(36);
output(3, 144) <= input(19);
output(3, 145) <= input(20);
output(3, 146) <= input(21);
output(3, 147) <= input(22);
output(3, 148) <= input(23);
output(3, 149) <= input(24);
output(3, 150) <= input(25);
output(3, 151) <= input(26);
output(3, 152) <= input(27);
output(3, 153) <= input(28);
output(3, 154) <= input(29);
output(3, 155) <= input(30);
output(3, 156) <= input(31);
output(3, 157) <= input(33);
output(3, 158) <= input(35);
output(3, 159) <= input(37);
output(3, 160) <= input(4);
output(3, 161) <= input(5);
output(3, 162) <= input(6);
output(3, 163) <= input(7);
output(3, 164) <= input(8);
output(3, 165) <= input(9);
output(3, 166) <= input(10);
output(3, 167) <= input(11);
output(3, 168) <= input(12);
output(3, 169) <= input(13);
output(3, 170) <= input(14);
output(3, 171) <= input(15);
output(3, 172) <= input(32);
output(3, 173) <= input(34);
output(3, 174) <= input(36);
output(3, 175) <= input(38);
output(3, 176) <= input(20);
output(3, 177) <= input(21);
output(3, 178) <= input(22);
output(3, 179) <= input(23);
output(3, 180) <= input(24);
output(3, 181) <= input(25);
output(3, 182) <= input(26);
output(3, 183) <= input(27);
output(3, 184) <= input(28);
output(3, 185) <= input(29);
output(3, 186) <= input(30);
output(3, 187) <= input(31);
output(3, 188) <= input(33);
output(3, 189) <= input(35);
output(3, 190) <= input(37);
output(3, 191) <= input(39);
output(3, 192) <= input(20);
output(3, 193) <= input(21);
output(3, 194) <= input(22);
output(3, 195) <= input(23);
output(3, 196) <= input(24);
output(3, 197) <= input(25);
output(3, 198) <= input(26);
output(3, 199) <= input(27);
output(3, 200) <= input(28);
output(3, 201) <= input(29);
output(3, 202) <= input(30);
output(3, 203) <= input(31);
output(3, 204) <= input(33);
output(3, 205) <= input(35);
output(3, 206) <= input(37);
output(3, 207) <= input(39);
output(3, 208) <= input(5);
output(3, 209) <= input(6);
output(3, 210) <= input(7);
output(3, 211) <= input(8);
output(3, 212) <= input(9);
output(3, 213) <= input(10);
output(3, 214) <= input(11);
output(3, 215) <= input(12);
output(3, 216) <= input(13);
output(3, 217) <= input(14);
output(3, 218) <= input(15);
output(3, 219) <= input(32);
output(3, 220) <= input(34);
output(3, 221) <= input(36);
output(3, 222) <= input(38);
output(3, 223) <= input(40);
output(3, 224) <= input(21);
output(3, 225) <= input(22);
output(3, 226) <= input(23);
output(3, 227) <= input(24);
output(3, 228) <= input(25);
output(3, 229) <= input(26);
output(3, 230) <= input(27);
output(3, 231) <= input(28);
output(3, 232) <= input(29);
output(3, 233) <= input(30);
output(3, 234) <= input(31);
output(3, 235) <= input(33);
output(3, 236) <= input(35);
output(3, 237) <= input(37);
output(3, 238) <= input(39);
output(3, 239) <= input(41);
output(3, 240) <= input(6);
output(3, 241) <= input(7);
output(3, 242) <= input(8);
output(3, 243) <= input(9);
output(3, 244) <= input(10);
output(3, 245) <= input(11);
output(3, 246) <= input(12);
output(3, 247) <= input(13);
output(3, 248) <= input(14);
output(3, 249) <= input(15);
output(3, 250) <= input(32);
output(3, 251) <= input(34);
output(3, 252) <= input(36);
output(3, 253) <= input(38);
output(3, 254) <= input(40);
output(3, 255) <= input(42);
output(4, 0) <= input(0);
output(4, 1) <= input(1);
output(4, 2) <= input(2);
output(4, 3) <= input(3);
output(4, 4) <= input(4);
output(4, 5) <= input(5);
output(4, 6) <= input(6);
output(4, 7) <= input(7);
output(4, 8) <= input(8);
output(4, 9) <= input(9);
output(4, 10) <= input(10);
output(4, 11) <= input(11);
output(4, 12) <= input(12);
output(4, 13) <= input(13);
output(4, 14) <= input(14);
output(4, 15) <= input(15);
output(4, 16) <= input(16);
output(4, 17) <= input(17);
output(4, 18) <= input(18);
output(4, 19) <= input(19);
output(4, 20) <= input(20);
output(4, 21) <= input(21);
output(4, 22) <= input(22);
output(4, 23) <= input(23);
output(4, 24) <= input(24);
output(4, 25) <= input(25);
output(4, 26) <= input(26);
output(4, 27) <= input(27);
output(4, 28) <= input(28);
output(4, 29) <= input(29);
output(4, 30) <= input(30);
output(4, 31) <= input(31);
output(4, 32) <= input(1);
output(4, 33) <= input(2);
output(4, 34) <= input(3);
output(4, 35) <= input(4);
output(4, 36) <= input(5);
output(4, 37) <= input(6);
output(4, 38) <= input(7);
output(4, 39) <= input(8);
output(4, 40) <= input(9);
output(4, 41) <= input(10);
output(4, 42) <= input(11);
output(4, 43) <= input(12);
output(4, 44) <= input(13);
output(4, 45) <= input(14);
output(4, 46) <= input(15);
output(4, 47) <= input(32);
output(4, 48) <= input(17);
output(4, 49) <= input(18);
output(4, 50) <= input(19);
output(4, 51) <= input(20);
output(4, 52) <= input(21);
output(4, 53) <= input(22);
output(4, 54) <= input(23);
output(4, 55) <= input(24);
output(4, 56) <= input(25);
output(4, 57) <= input(26);
output(4, 58) <= input(27);
output(4, 59) <= input(28);
output(4, 60) <= input(29);
output(4, 61) <= input(30);
output(4, 62) <= input(31);
output(4, 63) <= input(33);
output(4, 64) <= input(2);
output(4, 65) <= input(3);
output(4, 66) <= input(4);
output(4, 67) <= input(5);
output(4, 68) <= input(6);
output(4, 69) <= input(7);
output(4, 70) <= input(8);
output(4, 71) <= input(9);
output(4, 72) <= input(10);
output(4, 73) <= input(11);
output(4, 74) <= input(12);
output(4, 75) <= input(13);
output(4, 76) <= input(14);
output(4, 77) <= input(15);
output(4, 78) <= input(32);
output(4, 79) <= input(34);
output(4, 80) <= input(18);
output(4, 81) <= input(19);
output(4, 82) <= input(20);
output(4, 83) <= input(21);
output(4, 84) <= input(22);
output(4, 85) <= input(23);
output(4, 86) <= input(24);
output(4, 87) <= input(25);
output(4, 88) <= input(26);
output(4, 89) <= input(27);
output(4, 90) <= input(28);
output(4, 91) <= input(29);
output(4, 92) <= input(30);
output(4, 93) <= input(31);
output(4, 94) <= input(33);
output(4, 95) <= input(35);
output(4, 96) <= input(3);
output(4, 97) <= input(4);
output(4, 98) <= input(5);
output(4, 99) <= input(6);
output(4, 100) <= input(7);
output(4, 101) <= input(8);
output(4, 102) <= input(9);
output(4, 103) <= input(10);
output(4, 104) <= input(11);
output(4, 105) <= input(12);
output(4, 106) <= input(13);
output(4, 107) <= input(14);
output(4, 108) <= input(15);
output(4, 109) <= input(32);
output(4, 110) <= input(34);
output(4, 111) <= input(36);
output(4, 112) <= input(19);
output(4, 113) <= input(20);
output(4, 114) <= input(21);
output(4, 115) <= input(22);
output(4, 116) <= input(23);
output(4, 117) <= input(24);
output(4, 118) <= input(25);
output(4, 119) <= input(26);
output(4, 120) <= input(27);
output(4, 121) <= input(28);
output(4, 122) <= input(29);
output(4, 123) <= input(30);
output(4, 124) <= input(31);
output(4, 125) <= input(33);
output(4, 126) <= input(35);
output(4, 127) <= input(37);
output(4, 128) <= input(19);
output(4, 129) <= input(20);
output(4, 130) <= input(21);
output(4, 131) <= input(22);
output(4, 132) <= input(23);
output(4, 133) <= input(24);
output(4, 134) <= input(25);
output(4, 135) <= input(26);
output(4, 136) <= input(27);
output(4, 137) <= input(28);
output(4, 138) <= input(29);
output(4, 139) <= input(30);
output(4, 140) <= input(31);
output(4, 141) <= input(33);
output(4, 142) <= input(35);
output(4, 143) <= input(37);
output(4, 144) <= input(4);
output(4, 145) <= input(5);
output(4, 146) <= input(6);
output(4, 147) <= input(7);
output(4, 148) <= input(8);
output(4, 149) <= input(9);
output(4, 150) <= input(10);
output(4, 151) <= input(11);
output(4, 152) <= input(12);
output(4, 153) <= input(13);
output(4, 154) <= input(14);
output(4, 155) <= input(15);
output(4, 156) <= input(32);
output(4, 157) <= input(34);
output(4, 158) <= input(36);
output(4, 159) <= input(38);
output(4, 160) <= input(20);
output(4, 161) <= input(21);
output(4, 162) <= input(22);
output(4, 163) <= input(23);
output(4, 164) <= input(24);
output(4, 165) <= input(25);
output(4, 166) <= input(26);
output(4, 167) <= input(27);
output(4, 168) <= input(28);
output(4, 169) <= input(29);
output(4, 170) <= input(30);
output(4, 171) <= input(31);
output(4, 172) <= input(33);
output(4, 173) <= input(35);
output(4, 174) <= input(37);
output(4, 175) <= input(39);
output(4, 176) <= input(5);
output(4, 177) <= input(6);
output(4, 178) <= input(7);
output(4, 179) <= input(8);
output(4, 180) <= input(9);
output(4, 181) <= input(10);
output(4, 182) <= input(11);
output(4, 183) <= input(12);
output(4, 184) <= input(13);
output(4, 185) <= input(14);
output(4, 186) <= input(15);
output(4, 187) <= input(32);
output(4, 188) <= input(34);
output(4, 189) <= input(36);
output(4, 190) <= input(38);
output(4, 191) <= input(40);
output(4, 192) <= input(21);
output(4, 193) <= input(22);
output(4, 194) <= input(23);
output(4, 195) <= input(24);
output(4, 196) <= input(25);
output(4, 197) <= input(26);
output(4, 198) <= input(27);
output(4, 199) <= input(28);
output(4, 200) <= input(29);
output(4, 201) <= input(30);
output(4, 202) <= input(31);
output(4, 203) <= input(33);
output(4, 204) <= input(35);
output(4, 205) <= input(37);
output(4, 206) <= input(39);
output(4, 207) <= input(41);
output(4, 208) <= input(6);
output(4, 209) <= input(7);
output(4, 210) <= input(8);
output(4, 211) <= input(9);
output(4, 212) <= input(10);
output(4, 213) <= input(11);
output(4, 214) <= input(12);
output(4, 215) <= input(13);
output(4, 216) <= input(14);
output(4, 217) <= input(15);
output(4, 218) <= input(32);
output(4, 219) <= input(34);
output(4, 220) <= input(36);
output(4, 221) <= input(38);
output(4, 222) <= input(40);
output(4, 223) <= input(42);
output(4, 224) <= input(22);
output(4, 225) <= input(23);
output(4, 226) <= input(24);
output(4, 227) <= input(25);
output(4, 228) <= input(26);
output(4, 229) <= input(27);
output(4, 230) <= input(28);
output(4, 231) <= input(29);
output(4, 232) <= input(30);
output(4, 233) <= input(31);
output(4, 234) <= input(33);
output(4, 235) <= input(35);
output(4, 236) <= input(37);
output(4, 237) <= input(39);
output(4, 238) <= input(41);
output(4, 239) <= input(43);
output(4, 240) <= input(7);
output(4, 241) <= input(8);
output(4, 242) <= input(9);
output(4, 243) <= input(10);
output(4, 244) <= input(11);
output(4, 245) <= input(12);
output(4, 246) <= input(13);
output(4, 247) <= input(14);
output(4, 248) <= input(15);
output(4, 249) <= input(32);
output(4, 250) <= input(34);
output(4, 251) <= input(36);
output(4, 252) <= input(38);
output(4, 253) <= input(40);
output(4, 254) <= input(42);
output(4, 255) <= input(44);
output(5, 0) <= input(16);
output(5, 1) <= input(17);
output(5, 2) <= input(18);
output(5, 3) <= input(19);
output(5, 4) <= input(20);
output(5, 5) <= input(21);
output(5, 6) <= input(22);
output(5, 7) <= input(23);
output(5, 8) <= input(24);
output(5, 9) <= input(25);
output(5, 10) <= input(26);
output(5, 11) <= input(27);
output(5, 12) <= input(28);
output(5, 13) <= input(29);
output(5, 14) <= input(30);
output(5, 15) <= input(31);
output(5, 16) <= input(1);
output(5, 17) <= input(2);
output(5, 18) <= input(3);
output(5, 19) <= input(4);
output(5, 20) <= input(5);
output(5, 21) <= input(6);
output(5, 22) <= input(7);
output(5, 23) <= input(8);
output(5, 24) <= input(9);
output(5, 25) <= input(10);
output(5, 26) <= input(11);
output(5, 27) <= input(12);
output(5, 28) <= input(13);
output(5, 29) <= input(14);
output(5, 30) <= input(15);
output(5, 31) <= input(32);
output(5, 32) <= input(17);
output(5, 33) <= input(18);
output(5, 34) <= input(19);
output(5, 35) <= input(20);
output(5, 36) <= input(21);
output(5, 37) <= input(22);
output(5, 38) <= input(23);
output(5, 39) <= input(24);
output(5, 40) <= input(25);
output(5, 41) <= input(26);
output(5, 42) <= input(27);
output(5, 43) <= input(28);
output(5, 44) <= input(29);
output(5, 45) <= input(30);
output(5, 46) <= input(31);
output(5, 47) <= input(33);
output(5, 48) <= input(2);
output(5, 49) <= input(3);
output(5, 50) <= input(4);
output(5, 51) <= input(5);
output(5, 52) <= input(6);
output(5, 53) <= input(7);
output(5, 54) <= input(8);
output(5, 55) <= input(9);
output(5, 56) <= input(10);
output(5, 57) <= input(11);
output(5, 58) <= input(12);
output(5, 59) <= input(13);
output(5, 60) <= input(14);
output(5, 61) <= input(15);
output(5, 62) <= input(32);
output(5, 63) <= input(34);
output(5, 64) <= input(18);
output(5, 65) <= input(19);
output(5, 66) <= input(20);
output(5, 67) <= input(21);
output(5, 68) <= input(22);
output(5, 69) <= input(23);
output(5, 70) <= input(24);
output(5, 71) <= input(25);
output(5, 72) <= input(26);
output(5, 73) <= input(27);
output(5, 74) <= input(28);
output(5, 75) <= input(29);
output(5, 76) <= input(30);
output(5, 77) <= input(31);
output(5, 78) <= input(33);
output(5, 79) <= input(35);
output(5, 80) <= input(3);
output(5, 81) <= input(4);
output(5, 82) <= input(5);
output(5, 83) <= input(6);
output(5, 84) <= input(7);
output(5, 85) <= input(8);
output(5, 86) <= input(9);
output(5, 87) <= input(10);
output(5, 88) <= input(11);
output(5, 89) <= input(12);
output(5, 90) <= input(13);
output(5, 91) <= input(14);
output(5, 92) <= input(15);
output(5, 93) <= input(32);
output(5, 94) <= input(34);
output(5, 95) <= input(36);
output(5, 96) <= input(19);
output(5, 97) <= input(20);
output(5, 98) <= input(21);
output(5, 99) <= input(22);
output(5, 100) <= input(23);
output(5, 101) <= input(24);
output(5, 102) <= input(25);
output(5, 103) <= input(26);
output(5, 104) <= input(27);
output(5, 105) <= input(28);
output(5, 106) <= input(29);
output(5, 107) <= input(30);
output(5, 108) <= input(31);
output(5, 109) <= input(33);
output(5, 110) <= input(35);
output(5, 111) <= input(37);
output(5, 112) <= input(4);
output(5, 113) <= input(5);
output(5, 114) <= input(6);
output(5, 115) <= input(7);
output(5, 116) <= input(8);
output(5, 117) <= input(9);
output(5, 118) <= input(10);
output(5, 119) <= input(11);
output(5, 120) <= input(12);
output(5, 121) <= input(13);
output(5, 122) <= input(14);
output(5, 123) <= input(15);
output(5, 124) <= input(32);
output(5, 125) <= input(34);
output(5, 126) <= input(36);
output(5, 127) <= input(38);
output(5, 128) <= input(20);
output(5, 129) <= input(21);
output(5, 130) <= input(22);
output(5, 131) <= input(23);
output(5, 132) <= input(24);
output(5, 133) <= input(25);
output(5, 134) <= input(26);
output(5, 135) <= input(27);
output(5, 136) <= input(28);
output(5, 137) <= input(29);
output(5, 138) <= input(30);
output(5, 139) <= input(31);
output(5, 140) <= input(33);
output(5, 141) <= input(35);
output(5, 142) <= input(37);
output(5, 143) <= input(39);
output(5, 144) <= input(5);
output(5, 145) <= input(6);
output(5, 146) <= input(7);
output(5, 147) <= input(8);
output(5, 148) <= input(9);
output(5, 149) <= input(10);
output(5, 150) <= input(11);
output(5, 151) <= input(12);
output(5, 152) <= input(13);
output(5, 153) <= input(14);
output(5, 154) <= input(15);
output(5, 155) <= input(32);
output(5, 156) <= input(34);
output(5, 157) <= input(36);
output(5, 158) <= input(38);
output(5, 159) <= input(40);
output(5, 160) <= input(21);
output(5, 161) <= input(22);
output(5, 162) <= input(23);
output(5, 163) <= input(24);
output(5, 164) <= input(25);
output(5, 165) <= input(26);
output(5, 166) <= input(27);
output(5, 167) <= input(28);
output(5, 168) <= input(29);
output(5, 169) <= input(30);
output(5, 170) <= input(31);
output(5, 171) <= input(33);
output(5, 172) <= input(35);
output(5, 173) <= input(37);
output(5, 174) <= input(39);
output(5, 175) <= input(41);
output(5, 176) <= input(6);
output(5, 177) <= input(7);
output(5, 178) <= input(8);
output(5, 179) <= input(9);
output(5, 180) <= input(10);
output(5, 181) <= input(11);
output(5, 182) <= input(12);
output(5, 183) <= input(13);
output(5, 184) <= input(14);
output(5, 185) <= input(15);
output(5, 186) <= input(32);
output(5, 187) <= input(34);
output(5, 188) <= input(36);
output(5, 189) <= input(38);
output(5, 190) <= input(40);
output(5, 191) <= input(42);
output(5, 192) <= input(22);
output(5, 193) <= input(23);
output(5, 194) <= input(24);
output(5, 195) <= input(25);
output(5, 196) <= input(26);
output(5, 197) <= input(27);
output(5, 198) <= input(28);
output(5, 199) <= input(29);
output(5, 200) <= input(30);
output(5, 201) <= input(31);
output(5, 202) <= input(33);
output(5, 203) <= input(35);
output(5, 204) <= input(37);
output(5, 205) <= input(39);
output(5, 206) <= input(41);
output(5, 207) <= input(43);
output(5, 208) <= input(7);
output(5, 209) <= input(8);
output(5, 210) <= input(9);
output(5, 211) <= input(10);
output(5, 212) <= input(11);
output(5, 213) <= input(12);
output(5, 214) <= input(13);
output(5, 215) <= input(14);
output(5, 216) <= input(15);
output(5, 217) <= input(32);
output(5, 218) <= input(34);
output(5, 219) <= input(36);
output(5, 220) <= input(38);
output(5, 221) <= input(40);
output(5, 222) <= input(42);
output(5, 223) <= input(44);
output(5, 224) <= input(23);
output(5, 225) <= input(24);
output(5, 226) <= input(25);
output(5, 227) <= input(26);
output(5, 228) <= input(27);
output(5, 229) <= input(28);
output(5, 230) <= input(29);
output(5, 231) <= input(30);
output(5, 232) <= input(31);
output(5, 233) <= input(33);
output(5, 234) <= input(35);
output(5, 235) <= input(37);
output(5, 236) <= input(39);
output(5, 237) <= input(41);
output(5, 238) <= input(43);
output(5, 239) <= input(45);
output(5, 240) <= input(8);
output(5, 241) <= input(9);
output(5, 242) <= input(10);
output(5, 243) <= input(11);
output(5, 244) <= input(12);
output(5, 245) <= input(13);
output(5, 246) <= input(14);
output(5, 247) <= input(15);
output(5, 248) <= input(32);
output(5, 249) <= input(34);
output(5, 250) <= input(36);
output(5, 251) <= input(38);
output(5, 252) <= input(40);
output(5, 253) <= input(42);
output(5, 254) <= input(44);
output(5, 255) <= input(46);
when "1111" =>
output(0, 0) <= input(0);
output(0, 1) <= input(1);
output(0, 2) <= input(2);
output(0, 3) <= input(3);
output(0, 4) <= input(4);
output(0, 5) <= input(5);
output(0, 6) <= input(6);
output(0, 7) <= input(7);
output(0, 8) <= input(8);
output(0, 9) <= input(9);
output(0, 10) <= input(10);
output(0, 11) <= input(11);
output(0, 12) <= input(12);
output(0, 13) <= input(13);
output(0, 14) <= input(14);
output(0, 15) <= input(15);
output(0, 16) <= input(16);
output(0, 17) <= input(17);
output(0, 18) <= input(18);
output(0, 19) <= input(19);
output(0, 20) <= input(20);
output(0, 21) <= input(21);
output(0, 22) <= input(22);
output(0, 23) <= input(23);
output(0, 24) <= input(24);
output(0, 25) <= input(25);
output(0, 26) <= input(26);
output(0, 27) <= input(27);
output(0, 28) <= input(28);
output(0, 29) <= input(29);
output(0, 30) <= input(30);
output(0, 31) <= input(31);
output(0, 32) <= input(1);
output(0, 33) <= input(2);
output(0, 34) <= input(3);
output(0, 35) <= input(4);
output(0, 36) <= input(5);
output(0, 37) <= input(6);
output(0, 38) <= input(7);
output(0, 39) <= input(8);
output(0, 40) <= input(9);
output(0, 41) <= input(10);
output(0, 42) <= input(11);
output(0, 43) <= input(12);
output(0, 44) <= input(13);
output(0, 45) <= input(14);
output(0, 46) <= input(15);
output(0, 47) <= input(32);
output(0, 48) <= input(17);
output(0, 49) <= input(18);
output(0, 50) <= input(19);
output(0, 51) <= input(20);
output(0, 52) <= input(21);
output(0, 53) <= input(22);
output(0, 54) <= input(23);
output(0, 55) <= input(24);
output(0, 56) <= input(25);
output(0, 57) <= input(26);
output(0, 58) <= input(27);
output(0, 59) <= input(28);
output(0, 60) <= input(29);
output(0, 61) <= input(30);
output(0, 62) <= input(31);
output(0, 63) <= input(33);
output(0, 64) <= input(2);
output(0, 65) <= input(3);
output(0, 66) <= input(4);
output(0, 67) <= input(5);
output(0, 68) <= input(6);
output(0, 69) <= input(7);
output(0, 70) <= input(8);
output(0, 71) <= input(9);
output(0, 72) <= input(10);
output(0, 73) <= input(11);
output(0, 74) <= input(12);
output(0, 75) <= input(13);
output(0, 76) <= input(14);
output(0, 77) <= input(15);
output(0, 78) <= input(32);
output(0, 79) <= input(34);
output(0, 80) <= input(18);
output(0, 81) <= input(19);
output(0, 82) <= input(20);
output(0, 83) <= input(21);
output(0, 84) <= input(22);
output(0, 85) <= input(23);
output(0, 86) <= input(24);
output(0, 87) <= input(25);
output(0, 88) <= input(26);
output(0, 89) <= input(27);
output(0, 90) <= input(28);
output(0, 91) <= input(29);
output(0, 92) <= input(30);
output(0, 93) <= input(31);
output(0, 94) <= input(33);
output(0, 95) <= input(35);
output(0, 96) <= input(3);
output(0, 97) <= input(4);
output(0, 98) <= input(5);
output(0, 99) <= input(6);
output(0, 100) <= input(7);
output(0, 101) <= input(8);
output(0, 102) <= input(9);
output(0, 103) <= input(10);
output(0, 104) <= input(11);
output(0, 105) <= input(12);
output(0, 106) <= input(13);
output(0, 107) <= input(14);
output(0, 108) <= input(15);
output(0, 109) <= input(32);
output(0, 110) <= input(34);
output(0, 111) <= input(36);
output(0, 112) <= input(4);
output(0, 113) <= input(5);
output(0, 114) <= input(6);
output(0, 115) <= input(7);
output(0, 116) <= input(8);
output(0, 117) <= input(9);
output(0, 118) <= input(10);
output(0, 119) <= input(11);
output(0, 120) <= input(12);
output(0, 121) <= input(13);
output(0, 122) <= input(14);
output(0, 123) <= input(15);
output(0, 124) <= input(32);
output(0, 125) <= input(34);
output(0, 126) <= input(36);
output(0, 127) <= input(37);
output(0, 128) <= input(20);
output(0, 129) <= input(21);
output(0, 130) <= input(22);
output(0, 131) <= input(23);
output(0, 132) <= input(24);
output(0, 133) <= input(25);
output(0, 134) <= input(26);
output(0, 135) <= input(27);
output(0, 136) <= input(28);
output(0, 137) <= input(29);
output(0, 138) <= input(30);
output(0, 139) <= input(31);
output(0, 140) <= input(33);
output(0, 141) <= input(35);
output(0, 142) <= input(38);
output(0, 143) <= input(39);
output(0, 144) <= input(5);
output(0, 145) <= input(6);
output(0, 146) <= input(7);
output(0, 147) <= input(8);
output(0, 148) <= input(9);
output(0, 149) <= input(10);
output(0, 150) <= input(11);
output(0, 151) <= input(12);
output(0, 152) <= input(13);
output(0, 153) <= input(14);
output(0, 154) <= input(15);
output(0, 155) <= input(32);
output(0, 156) <= input(34);
output(0, 157) <= input(36);
output(0, 158) <= input(37);
output(0, 159) <= input(40);
output(0, 160) <= input(21);
output(0, 161) <= input(22);
output(0, 162) <= input(23);
output(0, 163) <= input(24);
output(0, 164) <= input(25);
output(0, 165) <= input(26);
output(0, 166) <= input(27);
output(0, 167) <= input(28);
output(0, 168) <= input(29);
output(0, 169) <= input(30);
output(0, 170) <= input(31);
output(0, 171) <= input(33);
output(0, 172) <= input(35);
output(0, 173) <= input(38);
output(0, 174) <= input(39);
output(0, 175) <= input(41);
output(0, 176) <= input(6);
output(0, 177) <= input(7);
output(0, 178) <= input(8);
output(0, 179) <= input(9);
output(0, 180) <= input(10);
output(0, 181) <= input(11);
output(0, 182) <= input(12);
output(0, 183) <= input(13);
output(0, 184) <= input(14);
output(0, 185) <= input(15);
output(0, 186) <= input(32);
output(0, 187) <= input(34);
output(0, 188) <= input(36);
output(0, 189) <= input(37);
output(0, 190) <= input(40);
output(0, 191) <= input(42);
output(0, 192) <= input(22);
output(0, 193) <= input(23);
output(0, 194) <= input(24);
output(0, 195) <= input(25);
output(0, 196) <= input(26);
output(0, 197) <= input(27);
output(0, 198) <= input(28);
output(0, 199) <= input(29);
output(0, 200) <= input(30);
output(0, 201) <= input(31);
output(0, 202) <= input(33);
output(0, 203) <= input(35);
output(0, 204) <= input(38);
output(0, 205) <= input(39);
output(0, 206) <= input(41);
output(0, 207) <= input(43);
output(0, 208) <= input(7);
output(0, 209) <= input(8);
output(0, 210) <= input(9);
output(0, 211) <= input(10);
output(0, 212) <= input(11);
output(0, 213) <= input(12);
output(0, 214) <= input(13);
output(0, 215) <= input(14);
output(0, 216) <= input(15);
output(0, 217) <= input(32);
output(0, 218) <= input(34);
output(0, 219) <= input(36);
output(0, 220) <= input(37);
output(0, 221) <= input(40);
output(0, 222) <= input(42);
output(0, 223) <= input(44);
output(0, 224) <= input(23);
output(0, 225) <= input(24);
output(0, 226) <= input(25);
output(0, 227) <= input(26);
output(0, 228) <= input(27);
output(0, 229) <= input(28);
output(0, 230) <= input(29);
output(0, 231) <= input(30);
output(0, 232) <= input(31);
output(0, 233) <= input(33);
output(0, 234) <= input(35);
output(0, 235) <= input(38);
output(0, 236) <= input(39);
output(0, 237) <= input(41);
output(0, 238) <= input(43);
output(0, 239) <= input(45);
output(0, 240) <= input(24);
output(0, 241) <= input(25);
output(0, 242) <= input(26);
output(0, 243) <= input(27);
output(0, 244) <= input(28);
output(0, 245) <= input(29);
output(0, 246) <= input(30);
output(0, 247) <= input(31);
output(0, 248) <= input(33);
output(0, 249) <= input(35);
output(0, 250) <= input(38);
output(0, 251) <= input(39);
output(0, 252) <= input(41);
output(0, 253) <= input(43);
output(0, 254) <= input(45);
output(0, 255) <= input(46);
output(1, 0) <= input(0);
output(1, 1) <= input(1);
output(1, 2) <= input(2);
output(1, 3) <= input(3);
output(1, 4) <= input(4);
output(1, 5) <= input(5);
output(1, 6) <= input(6);
output(1, 7) <= input(7);
output(1, 8) <= input(8);
output(1, 9) <= input(9);
output(1, 10) <= input(10);
output(1, 11) <= input(11);
output(1, 12) <= input(12);
output(1, 13) <= input(13);
output(1, 14) <= input(14);
output(1, 15) <= input(15);
output(1, 16) <= input(16);
output(1, 17) <= input(17);
output(1, 18) <= input(18);
output(1, 19) <= input(19);
output(1, 20) <= input(20);
output(1, 21) <= input(21);
output(1, 22) <= input(22);
output(1, 23) <= input(23);
output(1, 24) <= input(24);
output(1, 25) <= input(25);
output(1, 26) <= input(26);
output(1, 27) <= input(27);
output(1, 28) <= input(28);
output(1, 29) <= input(29);
output(1, 30) <= input(30);
output(1, 31) <= input(31);
output(1, 32) <= input(1);
output(1, 33) <= input(2);
output(1, 34) <= input(3);
output(1, 35) <= input(4);
output(1, 36) <= input(5);
output(1, 37) <= input(6);
output(1, 38) <= input(7);
output(1, 39) <= input(8);
output(1, 40) <= input(9);
output(1, 41) <= input(10);
output(1, 42) <= input(11);
output(1, 43) <= input(12);
output(1, 44) <= input(13);
output(1, 45) <= input(14);
output(1, 46) <= input(15);
output(1, 47) <= input(32);
output(1, 48) <= input(2);
output(1, 49) <= input(3);
output(1, 50) <= input(4);
output(1, 51) <= input(5);
output(1, 52) <= input(6);
output(1, 53) <= input(7);
output(1, 54) <= input(8);
output(1, 55) <= input(9);
output(1, 56) <= input(10);
output(1, 57) <= input(11);
output(1, 58) <= input(12);
output(1, 59) <= input(13);
output(1, 60) <= input(14);
output(1, 61) <= input(15);
output(1, 62) <= input(32);
output(1, 63) <= input(34);
output(1, 64) <= input(18);
output(1, 65) <= input(19);
output(1, 66) <= input(20);
output(1, 67) <= input(21);
output(1, 68) <= input(22);
output(1, 69) <= input(23);
output(1, 70) <= input(24);
output(1, 71) <= input(25);
output(1, 72) <= input(26);
output(1, 73) <= input(27);
output(1, 74) <= input(28);
output(1, 75) <= input(29);
output(1, 76) <= input(30);
output(1, 77) <= input(31);
output(1, 78) <= input(33);
output(1, 79) <= input(35);
output(1, 80) <= input(3);
output(1, 81) <= input(4);
output(1, 82) <= input(5);
output(1, 83) <= input(6);
output(1, 84) <= input(7);
output(1, 85) <= input(8);
output(1, 86) <= input(9);
output(1, 87) <= input(10);
output(1, 88) <= input(11);
output(1, 89) <= input(12);
output(1, 90) <= input(13);
output(1, 91) <= input(14);
output(1, 92) <= input(15);
output(1, 93) <= input(32);
output(1, 94) <= input(34);
output(1, 95) <= input(36);
output(1, 96) <= input(19);
output(1, 97) <= input(20);
output(1, 98) <= input(21);
output(1, 99) <= input(22);
output(1, 100) <= input(23);
output(1, 101) <= input(24);
output(1, 102) <= input(25);
output(1, 103) <= input(26);
output(1, 104) <= input(27);
output(1, 105) <= input(28);
output(1, 106) <= input(29);
output(1, 107) <= input(30);
output(1, 108) <= input(31);
output(1, 109) <= input(33);
output(1, 110) <= input(35);
output(1, 111) <= input(38);
output(1, 112) <= input(20);
output(1, 113) <= input(21);
output(1, 114) <= input(22);
output(1, 115) <= input(23);
output(1, 116) <= input(24);
output(1, 117) <= input(25);
output(1, 118) <= input(26);
output(1, 119) <= input(27);
output(1, 120) <= input(28);
output(1, 121) <= input(29);
output(1, 122) <= input(30);
output(1, 123) <= input(31);
output(1, 124) <= input(33);
output(1, 125) <= input(35);
output(1, 126) <= input(38);
output(1, 127) <= input(39);
output(1, 128) <= input(5);
output(1, 129) <= input(6);
output(1, 130) <= input(7);
output(1, 131) <= input(8);
output(1, 132) <= input(9);
output(1, 133) <= input(10);
output(1, 134) <= input(11);
output(1, 135) <= input(12);
output(1, 136) <= input(13);
output(1, 137) <= input(14);
output(1, 138) <= input(15);
output(1, 139) <= input(32);
output(1, 140) <= input(34);
output(1, 141) <= input(36);
output(1, 142) <= input(37);
output(1, 143) <= input(40);
output(1, 144) <= input(21);
output(1, 145) <= input(22);
output(1, 146) <= input(23);
output(1, 147) <= input(24);
output(1, 148) <= input(25);
output(1, 149) <= input(26);
output(1, 150) <= input(27);
output(1, 151) <= input(28);
output(1, 152) <= input(29);
output(1, 153) <= input(30);
output(1, 154) <= input(31);
output(1, 155) <= input(33);
output(1, 156) <= input(35);
output(1, 157) <= input(38);
output(1, 158) <= input(39);
output(1, 159) <= input(41);
output(1, 160) <= input(6);
output(1, 161) <= input(7);
output(1, 162) <= input(8);
output(1, 163) <= input(9);
output(1, 164) <= input(10);
output(1, 165) <= input(11);
output(1, 166) <= input(12);
output(1, 167) <= input(13);
output(1, 168) <= input(14);
output(1, 169) <= input(15);
output(1, 170) <= input(32);
output(1, 171) <= input(34);
output(1, 172) <= input(36);
output(1, 173) <= input(37);
output(1, 174) <= input(40);
output(1, 175) <= input(42);
output(1, 176) <= input(7);
output(1, 177) <= input(8);
output(1, 178) <= input(9);
output(1, 179) <= input(10);
output(1, 180) <= input(11);
output(1, 181) <= input(12);
output(1, 182) <= input(13);
output(1, 183) <= input(14);
output(1, 184) <= input(15);
output(1, 185) <= input(32);
output(1, 186) <= input(34);
output(1, 187) <= input(36);
output(1, 188) <= input(37);
output(1, 189) <= input(40);
output(1, 190) <= input(42);
output(1, 191) <= input(44);
output(1, 192) <= input(23);
output(1, 193) <= input(24);
output(1, 194) <= input(25);
output(1, 195) <= input(26);
output(1, 196) <= input(27);
output(1, 197) <= input(28);
output(1, 198) <= input(29);
output(1, 199) <= input(30);
output(1, 200) <= input(31);
output(1, 201) <= input(33);
output(1, 202) <= input(35);
output(1, 203) <= input(38);
output(1, 204) <= input(39);
output(1, 205) <= input(41);
output(1, 206) <= input(43);
output(1, 207) <= input(45);
output(1, 208) <= input(8);
output(1, 209) <= input(9);
output(1, 210) <= input(10);
output(1, 211) <= input(11);
output(1, 212) <= input(12);
output(1, 213) <= input(13);
output(1, 214) <= input(14);
output(1, 215) <= input(15);
output(1, 216) <= input(32);
output(1, 217) <= input(34);
output(1, 218) <= input(36);
output(1, 219) <= input(37);
output(1, 220) <= input(40);
output(1, 221) <= input(42);
output(1, 222) <= input(44);
output(1, 223) <= input(47);
output(1, 224) <= input(24);
output(1, 225) <= input(25);
output(1, 226) <= input(26);
output(1, 227) <= input(27);
output(1, 228) <= input(28);
output(1, 229) <= input(29);
output(1, 230) <= input(30);
output(1, 231) <= input(31);
output(1, 232) <= input(33);
output(1, 233) <= input(35);
output(1, 234) <= input(38);
output(1, 235) <= input(39);
output(1, 236) <= input(41);
output(1, 237) <= input(43);
output(1, 238) <= input(45);
output(1, 239) <= input(46);
output(1, 240) <= input(25);
output(1, 241) <= input(26);
output(1, 242) <= input(27);
output(1, 243) <= input(28);
output(1, 244) <= input(29);
output(1, 245) <= input(30);
output(1, 246) <= input(31);
output(1, 247) <= input(33);
output(1, 248) <= input(35);
output(1, 249) <= input(38);
output(1, 250) <= input(39);
output(1, 251) <= input(41);
output(1, 252) <= input(43);
output(1, 253) <= input(45);
output(1, 254) <= input(46);
output(1, 255) <= input(48);
output(2, 0) <= input(0);
output(2, 1) <= input(1);
output(2, 2) <= input(2);
output(2, 3) <= input(3);
output(2, 4) <= input(4);
output(2, 5) <= input(5);
output(2, 6) <= input(6);
output(2, 7) <= input(7);
output(2, 8) <= input(8);
output(2, 9) <= input(9);
output(2, 10) <= input(10);
output(2, 11) <= input(11);
output(2, 12) <= input(12);
output(2, 13) <= input(13);
output(2, 14) <= input(14);
output(2, 15) <= input(15);
output(2, 16) <= input(16);
output(2, 17) <= input(17);
output(2, 18) <= input(18);
output(2, 19) <= input(19);
output(2, 20) <= input(20);
output(2, 21) <= input(21);
output(2, 22) <= input(22);
output(2, 23) <= input(23);
output(2, 24) <= input(24);
output(2, 25) <= input(25);
output(2, 26) <= input(26);
output(2, 27) <= input(27);
output(2, 28) <= input(28);
output(2, 29) <= input(29);
output(2, 30) <= input(30);
output(2, 31) <= input(31);
output(2, 32) <= input(17);
output(2, 33) <= input(18);
output(2, 34) <= input(19);
output(2, 35) <= input(20);
output(2, 36) <= input(21);
output(2, 37) <= input(22);
output(2, 38) <= input(23);
output(2, 39) <= input(24);
output(2, 40) <= input(25);
output(2, 41) <= input(26);
output(2, 42) <= input(27);
output(2, 43) <= input(28);
output(2, 44) <= input(29);
output(2, 45) <= input(30);
output(2, 46) <= input(31);
output(2, 47) <= input(33);
output(2, 48) <= input(2);
output(2, 49) <= input(3);
output(2, 50) <= input(4);
output(2, 51) <= input(5);
output(2, 52) <= input(6);
output(2, 53) <= input(7);
output(2, 54) <= input(8);
output(2, 55) <= input(9);
output(2, 56) <= input(10);
output(2, 57) <= input(11);
output(2, 58) <= input(12);
output(2, 59) <= input(13);
output(2, 60) <= input(14);
output(2, 61) <= input(15);
output(2, 62) <= input(32);
output(2, 63) <= input(34);
output(2, 64) <= input(3);
output(2, 65) <= input(4);
output(2, 66) <= input(5);
output(2, 67) <= input(6);
output(2, 68) <= input(7);
output(2, 69) <= input(8);
output(2, 70) <= input(9);
output(2, 71) <= input(10);
output(2, 72) <= input(11);
output(2, 73) <= input(12);
output(2, 74) <= input(13);
output(2, 75) <= input(14);
output(2, 76) <= input(15);
output(2, 77) <= input(32);
output(2, 78) <= input(34);
output(2, 79) <= input(36);
output(2, 80) <= input(19);
output(2, 81) <= input(20);
output(2, 82) <= input(21);
output(2, 83) <= input(22);
output(2, 84) <= input(23);
output(2, 85) <= input(24);
output(2, 86) <= input(25);
output(2, 87) <= input(26);
output(2, 88) <= input(27);
output(2, 89) <= input(28);
output(2, 90) <= input(29);
output(2, 91) <= input(30);
output(2, 92) <= input(31);
output(2, 93) <= input(33);
output(2, 94) <= input(35);
output(2, 95) <= input(38);
output(2, 96) <= input(20);
output(2, 97) <= input(21);
output(2, 98) <= input(22);
output(2, 99) <= input(23);
output(2, 100) <= input(24);
output(2, 101) <= input(25);
output(2, 102) <= input(26);
output(2, 103) <= input(27);
output(2, 104) <= input(28);
output(2, 105) <= input(29);
output(2, 106) <= input(30);
output(2, 107) <= input(31);
output(2, 108) <= input(33);
output(2, 109) <= input(35);
output(2, 110) <= input(38);
output(2, 111) <= input(39);
output(2, 112) <= input(5);
output(2, 113) <= input(6);
output(2, 114) <= input(7);
output(2, 115) <= input(8);
output(2, 116) <= input(9);
output(2, 117) <= input(10);
output(2, 118) <= input(11);
output(2, 119) <= input(12);
output(2, 120) <= input(13);
output(2, 121) <= input(14);
output(2, 122) <= input(15);
output(2, 123) <= input(32);
output(2, 124) <= input(34);
output(2, 125) <= input(36);
output(2, 126) <= input(37);
output(2, 127) <= input(40);
output(2, 128) <= input(21);
output(2, 129) <= input(22);
output(2, 130) <= input(23);
output(2, 131) <= input(24);
output(2, 132) <= input(25);
output(2, 133) <= input(26);
output(2, 134) <= input(27);
output(2, 135) <= input(28);
output(2, 136) <= input(29);
output(2, 137) <= input(30);
output(2, 138) <= input(31);
output(2, 139) <= input(33);
output(2, 140) <= input(35);
output(2, 141) <= input(38);
output(2, 142) <= input(39);
output(2, 143) <= input(41);
output(2, 144) <= input(22);
output(2, 145) <= input(23);
output(2, 146) <= input(24);
output(2, 147) <= input(25);
output(2, 148) <= input(26);
output(2, 149) <= input(27);
output(2, 150) <= input(28);
output(2, 151) <= input(29);
output(2, 152) <= input(30);
output(2, 153) <= input(31);
output(2, 154) <= input(33);
output(2, 155) <= input(35);
output(2, 156) <= input(38);
output(2, 157) <= input(39);
output(2, 158) <= input(41);
output(2, 159) <= input(43);
output(2, 160) <= input(7);
output(2, 161) <= input(8);
output(2, 162) <= input(9);
output(2, 163) <= input(10);
output(2, 164) <= input(11);
output(2, 165) <= input(12);
output(2, 166) <= input(13);
output(2, 167) <= input(14);
output(2, 168) <= input(15);
output(2, 169) <= input(32);
output(2, 170) <= input(34);
output(2, 171) <= input(36);
output(2, 172) <= input(37);
output(2, 173) <= input(40);
output(2, 174) <= input(42);
output(2, 175) <= input(44);
output(2, 176) <= input(8);
output(2, 177) <= input(9);
output(2, 178) <= input(10);
output(2, 179) <= input(11);
output(2, 180) <= input(12);
output(2, 181) <= input(13);
output(2, 182) <= input(14);
output(2, 183) <= input(15);
output(2, 184) <= input(32);
output(2, 185) <= input(34);
output(2, 186) <= input(36);
output(2, 187) <= input(37);
output(2, 188) <= input(40);
output(2, 189) <= input(42);
output(2, 190) <= input(44);
output(2, 191) <= input(47);
output(2, 192) <= input(24);
output(2, 193) <= input(25);
output(2, 194) <= input(26);
output(2, 195) <= input(27);
output(2, 196) <= input(28);
output(2, 197) <= input(29);
output(2, 198) <= input(30);
output(2, 199) <= input(31);
output(2, 200) <= input(33);
output(2, 201) <= input(35);
output(2, 202) <= input(38);
output(2, 203) <= input(39);
output(2, 204) <= input(41);
output(2, 205) <= input(43);
output(2, 206) <= input(45);
output(2, 207) <= input(46);
output(2, 208) <= input(25);
output(2, 209) <= input(26);
output(2, 210) <= input(27);
output(2, 211) <= input(28);
output(2, 212) <= input(29);
output(2, 213) <= input(30);
output(2, 214) <= input(31);
output(2, 215) <= input(33);
output(2, 216) <= input(35);
output(2, 217) <= input(38);
output(2, 218) <= input(39);
output(2, 219) <= input(41);
output(2, 220) <= input(43);
output(2, 221) <= input(45);
output(2, 222) <= input(46);
output(2, 223) <= input(48);
output(2, 224) <= input(10);
output(2, 225) <= input(11);
output(2, 226) <= input(12);
output(2, 227) <= input(13);
output(2, 228) <= input(14);
output(2, 229) <= input(15);
output(2, 230) <= input(32);
output(2, 231) <= input(34);
output(2, 232) <= input(36);
output(2, 233) <= input(37);
output(2, 234) <= input(40);
output(2, 235) <= input(42);
output(2, 236) <= input(44);
output(2, 237) <= input(47);
output(2, 238) <= input(49);
output(2, 239) <= input(50);
output(2, 240) <= input(11);
output(2, 241) <= input(12);
output(2, 242) <= input(13);
output(2, 243) <= input(14);
output(2, 244) <= input(15);
output(2, 245) <= input(32);
output(2, 246) <= input(34);
output(2, 247) <= input(36);
output(2, 248) <= input(37);
output(2, 249) <= input(40);
output(2, 250) <= input(42);
output(2, 251) <= input(44);
output(2, 252) <= input(47);
output(2, 253) <= input(49);
output(2, 254) <= input(50);
output(2, 255) <= input(51);
output(3, 0) <= input(0);
output(3, 1) <= input(1);
output(3, 2) <= input(2);
output(3, 3) <= input(3);
output(3, 4) <= input(4);
output(3, 5) <= input(5);
output(3, 6) <= input(6);
output(3, 7) <= input(7);
output(3, 8) <= input(8);
output(3, 9) <= input(9);
output(3, 10) <= input(10);
output(3, 11) <= input(11);
output(3, 12) <= input(12);
output(3, 13) <= input(13);
output(3, 14) <= input(14);
output(3, 15) <= input(15);
output(3, 16) <= input(1);
output(3, 17) <= input(2);
output(3, 18) <= input(3);
output(3, 19) <= input(4);
output(3, 20) <= input(5);
output(3, 21) <= input(6);
output(3, 22) <= input(7);
output(3, 23) <= input(8);
output(3, 24) <= input(9);
output(3, 25) <= input(10);
output(3, 26) <= input(11);
output(3, 27) <= input(12);
output(3, 28) <= input(13);
output(3, 29) <= input(14);
output(3, 30) <= input(15);
output(3, 31) <= input(32);
output(3, 32) <= input(17);
output(3, 33) <= input(18);
output(3, 34) <= input(19);
output(3, 35) <= input(20);
output(3, 36) <= input(21);
output(3, 37) <= input(22);
output(3, 38) <= input(23);
output(3, 39) <= input(24);
output(3, 40) <= input(25);
output(3, 41) <= input(26);
output(3, 42) <= input(27);
output(3, 43) <= input(28);
output(3, 44) <= input(29);
output(3, 45) <= input(30);
output(3, 46) <= input(31);
output(3, 47) <= input(33);
output(3, 48) <= input(18);
output(3, 49) <= input(19);
output(3, 50) <= input(20);
output(3, 51) <= input(21);
output(3, 52) <= input(22);
output(3, 53) <= input(23);
output(3, 54) <= input(24);
output(3, 55) <= input(25);
output(3, 56) <= input(26);
output(3, 57) <= input(27);
output(3, 58) <= input(28);
output(3, 59) <= input(29);
output(3, 60) <= input(30);
output(3, 61) <= input(31);
output(3, 62) <= input(33);
output(3, 63) <= input(35);
output(3, 64) <= input(19);
output(3, 65) <= input(20);
output(3, 66) <= input(21);
output(3, 67) <= input(22);
output(3, 68) <= input(23);
output(3, 69) <= input(24);
output(3, 70) <= input(25);
output(3, 71) <= input(26);
output(3, 72) <= input(27);
output(3, 73) <= input(28);
output(3, 74) <= input(29);
output(3, 75) <= input(30);
output(3, 76) <= input(31);
output(3, 77) <= input(33);
output(3, 78) <= input(35);
output(3, 79) <= input(38);
output(3, 80) <= input(4);
output(3, 81) <= input(5);
output(3, 82) <= input(6);
output(3, 83) <= input(7);
output(3, 84) <= input(8);
output(3, 85) <= input(9);
output(3, 86) <= input(10);
output(3, 87) <= input(11);
output(3, 88) <= input(12);
output(3, 89) <= input(13);
output(3, 90) <= input(14);
output(3, 91) <= input(15);
output(3, 92) <= input(32);
output(3, 93) <= input(34);
output(3, 94) <= input(36);
output(3, 95) <= input(37);
output(3, 96) <= input(5);
output(3, 97) <= input(6);
output(3, 98) <= input(7);
output(3, 99) <= input(8);
output(3, 100) <= input(9);
output(3, 101) <= input(10);
output(3, 102) <= input(11);
output(3, 103) <= input(12);
output(3, 104) <= input(13);
output(3, 105) <= input(14);
output(3, 106) <= input(15);
output(3, 107) <= input(32);
output(3, 108) <= input(34);
output(3, 109) <= input(36);
output(3, 110) <= input(37);
output(3, 111) <= input(40);
output(3, 112) <= input(6);
output(3, 113) <= input(7);
output(3, 114) <= input(8);
output(3, 115) <= input(9);
output(3, 116) <= input(10);
output(3, 117) <= input(11);
output(3, 118) <= input(12);
output(3, 119) <= input(13);
output(3, 120) <= input(14);
output(3, 121) <= input(15);
output(3, 122) <= input(32);
output(3, 123) <= input(34);
output(3, 124) <= input(36);
output(3, 125) <= input(37);
output(3, 126) <= input(40);
output(3, 127) <= input(42);
output(3, 128) <= input(22);
output(3, 129) <= input(23);
output(3, 130) <= input(24);
output(3, 131) <= input(25);
output(3, 132) <= input(26);
output(3, 133) <= input(27);
output(3, 134) <= input(28);
output(3, 135) <= input(29);
output(3, 136) <= input(30);
output(3, 137) <= input(31);
output(3, 138) <= input(33);
output(3, 139) <= input(35);
output(3, 140) <= input(38);
output(3, 141) <= input(39);
output(3, 142) <= input(41);
output(3, 143) <= input(43);
output(3, 144) <= input(23);
output(3, 145) <= input(24);
output(3, 146) <= input(25);
output(3, 147) <= input(26);
output(3, 148) <= input(27);
output(3, 149) <= input(28);
output(3, 150) <= input(29);
output(3, 151) <= input(30);
output(3, 152) <= input(31);
output(3, 153) <= input(33);
output(3, 154) <= input(35);
output(3, 155) <= input(38);
output(3, 156) <= input(39);
output(3, 157) <= input(41);
output(3, 158) <= input(43);
output(3, 159) <= input(45);
output(3, 160) <= input(8);
output(3, 161) <= input(9);
output(3, 162) <= input(10);
output(3, 163) <= input(11);
output(3, 164) <= input(12);
output(3, 165) <= input(13);
output(3, 166) <= input(14);
output(3, 167) <= input(15);
output(3, 168) <= input(32);
output(3, 169) <= input(34);
output(3, 170) <= input(36);
output(3, 171) <= input(37);
output(3, 172) <= input(40);
output(3, 173) <= input(42);
output(3, 174) <= input(44);
output(3, 175) <= input(47);
output(3, 176) <= input(9);
output(3, 177) <= input(10);
output(3, 178) <= input(11);
output(3, 179) <= input(12);
output(3, 180) <= input(13);
output(3, 181) <= input(14);
output(3, 182) <= input(15);
output(3, 183) <= input(32);
output(3, 184) <= input(34);
output(3, 185) <= input(36);
output(3, 186) <= input(37);
output(3, 187) <= input(40);
output(3, 188) <= input(42);
output(3, 189) <= input(44);
output(3, 190) <= input(47);
output(3, 191) <= input(49);
output(3, 192) <= input(10);
output(3, 193) <= input(11);
output(3, 194) <= input(12);
output(3, 195) <= input(13);
output(3, 196) <= input(14);
output(3, 197) <= input(15);
output(3, 198) <= input(32);
output(3, 199) <= input(34);
output(3, 200) <= input(36);
output(3, 201) <= input(37);
output(3, 202) <= input(40);
output(3, 203) <= input(42);
output(3, 204) <= input(44);
output(3, 205) <= input(47);
output(3, 206) <= input(49);
output(3, 207) <= input(50);
output(3, 208) <= input(26);
output(3, 209) <= input(27);
output(3, 210) <= input(28);
output(3, 211) <= input(29);
output(3, 212) <= input(30);
output(3, 213) <= input(31);
output(3, 214) <= input(33);
output(3, 215) <= input(35);
output(3, 216) <= input(38);
output(3, 217) <= input(39);
output(3, 218) <= input(41);
output(3, 219) <= input(43);
output(3, 220) <= input(45);
output(3, 221) <= input(46);
output(3, 222) <= input(48);
output(3, 223) <= input(52);
output(3, 224) <= input(27);
output(3, 225) <= input(28);
output(3, 226) <= input(29);
output(3, 227) <= input(30);
output(3, 228) <= input(31);
output(3, 229) <= input(33);
output(3, 230) <= input(35);
output(3, 231) <= input(38);
output(3, 232) <= input(39);
output(3, 233) <= input(41);
output(3, 234) <= input(43);
output(3, 235) <= input(45);
output(3, 236) <= input(46);
output(3, 237) <= input(48);
output(3, 238) <= input(52);
output(3, 239) <= input(53);
output(3, 240) <= input(28);
output(3, 241) <= input(29);
output(3, 242) <= input(30);
output(3, 243) <= input(31);
output(3, 244) <= input(33);
output(3, 245) <= input(35);
output(3, 246) <= input(38);
output(3, 247) <= input(39);
output(3, 248) <= input(41);
output(3, 249) <= input(43);
output(3, 250) <= input(45);
output(3, 251) <= input(46);
output(3, 252) <= input(48);
output(3, 253) <= input(52);
output(3, 254) <= input(53);
output(3, 255) <= input(54);
output(4, 0) <= input(0);
output(4, 1) <= input(1);
output(4, 2) <= input(2);
output(4, 3) <= input(3);
output(4, 4) <= input(4);
output(4, 5) <= input(5);
output(4, 6) <= input(6);
output(4, 7) <= input(7);
output(4, 8) <= input(8);
output(4, 9) <= input(9);
output(4, 10) <= input(10);
output(4, 11) <= input(11);
output(4, 12) <= input(12);
output(4, 13) <= input(13);
output(4, 14) <= input(14);
output(4, 15) <= input(15);
output(4, 16) <= input(1);
output(4, 17) <= input(2);
output(4, 18) <= input(3);
output(4, 19) <= input(4);
output(4, 20) <= input(5);
output(4, 21) <= input(6);
output(4, 22) <= input(7);
output(4, 23) <= input(8);
output(4, 24) <= input(9);
output(4, 25) <= input(10);
output(4, 26) <= input(11);
output(4, 27) <= input(12);
output(4, 28) <= input(13);
output(4, 29) <= input(14);
output(4, 30) <= input(15);
output(4, 31) <= input(32);
output(4, 32) <= input(2);
output(4, 33) <= input(3);
output(4, 34) <= input(4);
output(4, 35) <= input(5);
output(4, 36) <= input(6);
output(4, 37) <= input(7);
output(4, 38) <= input(8);
output(4, 39) <= input(9);
output(4, 40) <= input(10);
output(4, 41) <= input(11);
output(4, 42) <= input(12);
output(4, 43) <= input(13);
output(4, 44) <= input(14);
output(4, 45) <= input(15);
output(4, 46) <= input(32);
output(4, 47) <= input(34);
output(4, 48) <= input(3);
output(4, 49) <= input(4);
output(4, 50) <= input(5);
output(4, 51) <= input(6);
output(4, 52) <= input(7);
output(4, 53) <= input(8);
output(4, 54) <= input(9);
output(4, 55) <= input(10);
output(4, 56) <= input(11);
output(4, 57) <= input(12);
output(4, 58) <= input(13);
output(4, 59) <= input(14);
output(4, 60) <= input(15);
output(4, 61) <= input(32);
output(4, 62) <= input(34);
output(4, 63) <= input(36);
output(4, 64) <= input(4);
output(4, 65) <= input(5);
output(4, 66) <= input(6);
output(4, 67) <= input(7);
output(4, 68) <= input(8);
output(4, 69) <= input(9);
output(4, 70) <= input(10);
output(4, 71) <= input(11);
output(4, 72) <= input(12);
output(4, 73) <= input(13);
output(4, 74) <= input(14);
output(4, 75) <= input(15);
output(4, 76) <= input(32);
output(4, 77) <= input(34);
output(4, 78) <= input(36);
output(4, 79) <= input(37);
output(4, 80) <= input(20);
output(4, 81) <= input(21);
output(4, 82) <= input(22);
output(4, 83) <= input(23);
output(4, 84) <= input(24);
output(4, 85) <= input(25);
output(4, 86) <= input(26);
output(4, 87) <= input(27);
output(4, 88) <= input(28);
output(4, 89) <= input(29);
output(4, 90) <= input(30);
output(4, 91) <= input(31);
output(4, 92) <= input(33);
output(4, 93) <= input(35);
output(4, 94) <= input(38);
output(4, 95) <= input(39);
output(4, 96) <= input(21);
output(4, 97) <= input(22);
output(4, 98) <= input(23);
output(4, 99) <= input(24);
output(4, 100) <= input(25);
output(4, 101) <= input(26);
output(4, 102) <= input(27);
output(4, 103) <= input(28);
output(4, 104) <= input(29);
output(4, 105) <= input(30);
output(4, 106) <= input(31);
output(4, 107) <= input(33);
output(4, 108) <= input(35);
output(4, 109) <= input(38);
output(4, 110) <= input(39);
output(4, 111) <= input(41);
output(4, 112) <= input(22);
output(4, 113) <= input(23);
output(4, 114) <= input(24);
output(4, 115) <= input(25);
output(4, 116) <= input(26);
output(4, 117) <= input(27);
output(4, 118) <= input(28);
output(4, 119) <= input(29);
output(4, 120) <= input(30);
output(4, 121) <= input(31);
output(4, 122) <= input(33);
output(4, 123) <= input(35);
output(4, 124) <= input(38);
output(4, 125) <= input(39);
output(4, 126) <= input(41);
output(4, 127) <= input(43);
output(4, 128) <= input(23);
output(4, 129) <= input(24);
output(4, 130) <= input(25);
output(4, 131) <= input(26);
output(4, 132) <= input(27);
output(4, 133) <= input(28);
output(4, 134) <= input(29);
output(4, 135) <= input(30);
output(4, 136) <= input(31);
output(4, 137) <= input(33);
output(4, 138) <= input(35);
output(4, 139) <= input(38);
output(4, 140) <= input(39);
output(4, 141) <= input(41);
output(4, 142) <= input(43);
output(4, 143) <= input(45);
output(4, 144) <= input(24);
output(4, 145) <= input(25);
output(4, 146) <= input(26);
output(4, 147) <= input(27);
output(4, 148) <= input(28);
output(4, 149) <= input(29);
output(4, 150) <= input(30);
output(4, 151) <= input(31);
output(4, 152) <= input(33);
output(4, 153) <= input(35);
output(4, 154) <= input(38);
output(4, 155) <= input(39);
output(4, 156) <= input(41);
output(4, 157) <= input(43);
output(4, 158) <= input(45);
output(4, 159) <= input(46);
output(4, 160) <= input(9);
output(4, 161) <= input(10);
output(4, 162) <= input(11);
output(4, 163) <= input(12);
output(4, 164) <= input(13);
output(4, 165) <= input(14);
output(4, 166) <= input(15);
output(4, 167) <= input(32);
output(4, 168) <= input(34);
output(4, 169) <= input(36);
output(4, 170) <= input(37);
output(4, 171) <= input(40);
output(4, 172) <= input(42);
output(4, 173) <= input(44);
output(4, 174) <= input(47);
output(4, 175) <= input(49);
output(4, 176) <= input(10);
output(4, 177) <= input(11);
output(4, 178) <= input(12);
output(4, 179) <= input(13);
output(4, 180) <= input(14);
output(4, 181) <= input(15);
output(4, 182) <= input(32);
output(4, 183) <= input(34);
output(4, 184) <= input(36);
output(4, 185) <= input(37);
output(4, 186) <= input(40);
output(4, 187) <= input(42);
output(4, 188) <= input(44);
output(4, 189) <= input(47);
output(4, 190) <= input(49);
output(4, 191) <= input(50);
output(4, 192) <= input(11);
output(4, 193) <= input(12);
output(4, 194) <= input(13);
output(4, 195) <= input(14);
output(4, 196) <= input(15);
output(4, 197) <= input(32);
output(4, 198) <= input(34);
output(4, 199) <= input(36);
output(4, 200) <= input(37);
output(4, 201) <= input(40);
output(4, 202) <= input(42);
output(4, 203) <= input(44);
output(4, 204) <= input(47);
output(4, 205) <= input(49);
output(4, 206) <= input(50);
output(4, 207) <= input(51);
output(4, 208) <= input(12);
output(4, 209) <= input(13);
output(4, 210) <= input(14);
output(4, 211) <= input(15);
output(4, 212) <= input(32);
output(4, 213) <= input(34);
output(4, 214) <= input(36);
output(4, 215) <= input(37);
output(4, 216) <= input(40);
output(4, 217) <= input(42);
output(4, 218) <= input(44);
output(4, 219) <= input(47);
output(4, 220) <= input(49);
output(4, 221) <= input(50);
output(4, 222) <= input(51);
output(4, 223) <= input(55);
output(4, 224) <= input(13);
output(4, 225) <= input(14);
output(4, 226) <= input(15);
output(4, 227) <= input(32);
output(4, 228) <= input(34);
output(4, 229) <= input(36);
output(4, 230) <= input(37);
output(4, 231) <= input(40);
output(4, 232) <= input(42);
output(4, 233) <= input(44);
output(4, 234) <= input(47);
output(4, 235) <= input(49);
output(4, 236) <= input(50);
output(4, 237) <= input(51);
output(4, 238) <= input(55);
output(4, 239) <= input(56);
output(4, 240) <= input(14);
output(4, 241) <= input(15);
output(4, 242) <= input(32);
output(4, 243) <= input(34);
output(4, 244) <= input(36);
output(4, 245) <= input(37);
output(4, 246) <= input(40);
output(4, 247) <= input(42);
output(4, 248) <= input(44);
output(4, 249) <= input(47);
output(4, 250) <= input(49);
output(4, 251) <= input(50);
output(4, 252) <= input(51);
output(4, 253) <= input(55);
output(4, 254) <= input(56);
output(4, 255) <= input(57);
output(5, 0) <= input(16);
output(5, 1) <= input(17);
output(5, 2) <= input(18);
output(5, 3) <= input(19);
output(5, 4) <= input(20);
output(5, 5) <= input(21);
output(5, 6) <= input(22);
output(5, 7) <= input(23);
output(5, 8) <= input(24);
output(5, 9) <= input(25);
output(5, 10) <= input(26);
output(5, 11) <= input(27);
output(5, 12) <= input(28);
output(5, 13) <= input(29);
output(5, 14) <= input(30);
output(5, 15) <= input(31);
output(5, 16) <= input(17);
output(5, 17) <= input(18);
output(5, 18) <= input(19);
output(5, 19) <= input(20);
output(5, 20) <= input(21);
output(5, 21) <= input(22);
output(5, 22) <= input(23);
output(5, 23) <= input(24);
output(5, 24) <= input(25);
output(5, 25) <= input(26);
output(5, 26) <= input(27);
output(5, 27) <= input(28);
output(5, 28) <= input(29);
output(5, 29) <= input(30);
output(5, 30) <= input(31);
output(5, 31) <= input(33);
output(5, 32) <= input(18);
output(5, 33) <= input(19);
output(5, 34) <= input(20);
output(5, 35) <= input(21);
output(5, 36) <= input(22);
output(5, 37) <= input(23);
output(5, 38) <= input(24);
output(5, 39) <= input(25);
output(5, 40) <= input(26);
output(5, 41) <= input(27);
output(5, 42) <= input(28);
output(5, 43) <= input(29);
output(5, 44) <= input(30);
output(5, 45) <= input(31);
output(5, 46) <= input(33);
output(5, 47) <= input(35);
output(5, 48) <= input(19);
output(5, 49) <= input(20);
output(5, 50) <= input(21);
output(5, 51) <= input(22);
output(5, 52) <= input(23);
output(5, 53) <= input(24);
output(5, 54) <= input(25);
output(5, 55) <= input(26);
output(5, 56) <= input(27);
output(5, 57) <= input(28);
output(5, 58) <= input(29);
output(5, 59) <= input(30);
output(5, 60) <= input(31);
output(5, 61) <= input(33);
output(5, 62) <= input(35);
output(5, 63) <= input(38);
output(5, 64) <= input(20);
output(5, 65) <= input(21);
output(5, 66) <= input(22);
output(5, 67) <= input(23);
output(5, 68) <= input(24);
output(5, 69) <= input(25);
output(5, 70) <= input(26);
output(5, 71) <= input(27);
output(5, 72) <= input(28);
output(5, 73) <= input(29);
output(5, 74) <= input(30);
output(5, 75) <= input(31);
output(5, 76) <= input(33);
output(5, 77) <= input(35);
output(5, 78) <= input(38);
output(5, 79) <= input(39);
output(5, 80) <= input(21);
output(5, 81) <= input(22);
output(5, 82) <= input(23);
output(5, 83) <= input(24);
output(5, 84) <= input(25);
output(5, 85) <= input(26);
output(5, 86) <= input(27);
output(5, 87) <= input(28);
output(5, 88) <= input(29);
output(5, 89) <= input(30);
output(5, 90) <= input(31);
output(5, 91) <= input(33);
output(5, 92) <= input(35);
output(5, 93) <= input(38);
output(5, 94) <= input(39);
output(5, 95) <= input(41);
output(5, 96) <= input(22);
output(5, 97) <= input(23);
output(5, 98) <= input(24);
output(5, 99) <= input(25);
output(5, 100) <= input(26);
output(5, 101) <= input(27);
output(5, 102) <= input(28);
output(5, 103) <= input(29);
output(5, 104) <= input(30);
output(5, 105) <= input(31);
output(5, 106) <= input(33);
output(5, 107) <= input(35);
output(5, 108) <= input(38);
output(5, 109) <= input(39);
output(5, 110) <= input(41);
output(5, 111) <= input(43);
output(5, 112) <= input(23);
output(5, 113) <= input(24);
output(5, 114) <= input(25);
output(5, 115) <= input(26);
output(5, 116) <= input(27);
output(5, 117) <= input(28);
output(5, 118) <= input(29);
output(5, 119) <= input(30);
output(5, 120) <= input(31);
output(5, 121) <= input(33);
output(5, 122) <= input(35);
output(5, 123) <= input(38);
output(5, 124) <= input(39);
output(5, 125) <= input(41);
output(5, 126) <= input(43);
output(5, 127) <= input(45);
output(5, 128) <= input(24);
output(5, 129) <= input(25);
output(5, 130) <= input(26);
output(5, 131) <= input(27);
output(5, 132) <= input(28);
output(5, 133) <= input(29);
output(5, 134) <= input(30);
output(5, 135) <= input(31);
output(5, 136) <= input(33);
output(5, 137) <= input(35);
output(5, 138) <= input(38);
output(5, 139) <= input(39);
output(5, 140) <= input(41);
output(5, 141) <= input(43);
output(5, 142) <= input(45);
output(5, 143) <= input(46);
output(5, 144) <= input(25);
output(5, 145) <= input(26);
output(5, 146) <= input(27);
output(5, 147) <= input(28);
output(5, 148) <= input(29);
output(5, 149) <= input(30);
output(5, 150) <= input(31);
output(5, 151) <= input(33);
output(5, 152) <= input(35);
output(5, 153) <= input(38);
output(5, 154) <= input(39);
output(5, 155) <= input(41);
output(5, 156) <= input(43);
output(5, 157) <= input(45);
output(5, 158) <= input(46);
output(5, 159) <= input(48);
output(5, 160) <= input(26);
output(5, 161) <= input(27);
output(5, 162) <= input(28);
output(5, 163) <= input(29);
output(5, 164) <= input(30);
output(5, 165) <= input(31);
output(5, 166) <= input(33);
output(5, 167) <= input(35);
output(5, 168) <= input(38);
output(5, 169) <= input(39);
output(5, 170) <= input(41);
output(5, 171) <= input(43);
output(5, 172) <= input(45);
output(5, 173) <= input(46);
output(5, 174) <= input(48);
output(5, 175) <= input(52);
output(5, 176) <= input(27);
output(5, 177) <= input(28);
output(5, 178) <= input(29);
output(5, 179) <= input(30);
output(5, 180) <= input(31);
output(5, 181) <= input(33);
output(5, 182) <= input(35);
output(5, 183) <= input(38);
output(5, 184) <= input(39);
output(5, 185) <= input(41);
output(5, 186) <= input(43);
output(5, 187) <= input(45);
output(5, 188) <= input(46);
output(5, 189) <= input(48);
output(5, 190) <= input(52);
output(5, 191) <= input(53);
output(5, 192) <= input(28);
output(5, 193) <= input(29);
output(5, 194) <= input(30);
output(5, 195) <= input(31);
output(5, 196) <= input(33);
output(5, 197) <= input(35);
output(5, 198) <= input(38);
output(5, 199) <= input(39);
output(5, 200) <= input(41);
output(5, 201) <= input(43);
output(5, 202) <= input(45);
output(5, 203) <= input(46);
output(5, 204) <= input(48);
output(5, 205) <= input(52);
output(5, 206) <= input(53);
output(5, 207) <= input(54);
output(5, 208) <= input(29);
output(5, 209) <= input(30);
output(5, 210) <= input(31);
output(5, 211) <= input(33);
output(5, 212) <= input(35);
output(5, 213) <= input(38);
output(5, 214) <= input(39);
output(5, 215) <= input(41);
output(5, 216) <= input(43);
output(5, 217) <= input(45);
output(5, 218) <= input(46);
output(5, 219) <= input(48);
output(5, 220) <= input(52);
output(5, 221) <= input(53);
output(5, 222) <= input(54);
output(5, 223) <= input(58);
output(5, 224) <= input(30);
output(5, 225) <= input(31);
output(5, 226) <= input(33);
output(5, 227) <= input(35);
output(5, 228) <= input(38);
output(5, 229) <= input(39);
output(5, 230) <= input(41);
output(5, 231) <= input(43);
output(5, 232) <= input(45);
output(5, 233) <= input(46);
output(5, 234) <= input(48);
output(5, 235) <= input(52);
output(5, 236) <= input(53);
output(5, 237) <= input(54);
output(5, 238) <= input(58);
output(5, 239) <= input(59);
output(5, 240) <= input(31);
output(5, 241) <= input(33);
output(5, 242) <= input(35);
output(5, 243) <= input(38);
output(5, 244) <= input(39);
output(5, 245) <= input(41);
output(5, 246) <= input(43);
output(5, 247) <= input(45);
output(5, 248) <= input(46);
output(5, 249) <= input(48);
output(5, 250) <= input(52);
output(5, 251) <= input(53);
output(5, 252) <= input(54);
output(5, 253) <= input(58);
output(5, 254) <= input(59);
output(5, 255) <= input(60);
when others => for i in 0 to 7 loop for j in 0 to 255 loop output(i,j) <= "00000000"; end loop; end loop;
end case;
elsif control = "011" then 
case iteration_control is
when "0000" =>
output(0, 0) <= input(0);
output(0, 1) <= input(1);
output(0, 2) <= input(2);
output(0, 3) <= input(3);
output(0, 4) <= input(4);
output(0, 5) <= input(5);
output(0, 6) <= input(6);
output(0, 7) <= input(7);
output(0, 8) <= input(8);
output(0, 9) <= input(9);
output(0, 10) <= input(10);
output(0, 11) <= input(11);
output(0, 12) <= input(12);
output(0, 13) <= input(13);
output(0, 14) <= input(14);
output(0, 15) <= input(15);
output(0, 16) <= input(1);
output(0, 17) <= input(2);
output(0, 18) <= input(3);
output(0, 19) <= input(4);
output(0, 20) <= input(5);
output(0, 21) <= input(6);
output(0, 22) <= input(7);
output(0, 23) <= input(8);
output(0, 24) <= input(9);
output(0, 25) <= input(10);
output(0, 26) <= input(11);
output(0, 27) <= input(12);
output(0, 28) <= input(13);
output(0, 29) <= input(14);
output(0, 30) <= input(15);
output(0, 31) <= input(16);
output(0, 32) <= input(2);
output(0, 33) <= input(3);
output(0, 34) <= input(4);
output(0, 35) <= input(5);
output(0, 36) <= input(6);
output(0, 37) <= input(7);
output(0, 38) <= input(8);
output(0, 39) <= input(9);
output(0, 40) <= input(10);
output(0, 41) <= input(11);
output(0, 42) <= input(12);
output(0, 43) <= input(13);
output(0, 44) <= input(14);
output(0, 45) <= input(15);
output(0, 46) <= input(16);
output(0, 47) <= input(17);
output(0, 48) <= input(3);
output(0, 49) <= input(4);
output(0, 50) <= input(5);
output(0, 51) <= input(6);
output(0, 52) <= input(7);
output(0, 53) <= input(8);
output(0, 54) <= input(9);
output(0, 55) <= input(10);
output(0, 56) <= input(11);
output(0, 57) <= input(12);
output(0, 58) <= input(13);
output(0, 59) <= input(14);
output(0, 60) <= input(15);
output(0, 61) <= input(16);
output(0, 62) <= input(17);
output(0, 63) <= input(18);
output(0, 64) <= input(4);
output(0, 65) <= input(5);
output(0, 66) <= input(6);
output(0, 67) <= input(7);
output(0, 68) <= input(8);
output(0, 69) <= input(9);
output(0, 70) <= input(10);
output(0, 71) <= input(11);
output(0, 72) <= input(12);
output(0, 73) <= input(13);
output(0, 74) <= input(14);
output(0, 75) <= input(15);
output(0, 76) <= input(16);
output(0, 77) <= input(17);
output(0, 78) <= input(18);
output(0, 79) <= input(19);
output(0, 80) <= input(5);
output(0, 81) <= input(6);
output(0, 82) <= input(7);
output(0, 83) <= input(8);
output(0, 84) <= input(9);
output(0, 85) <= input(10);
output(0, 86) <= input(11);
output(0, 87) <= input(12);
output(0, 88) <= input(13);
output(0, 89) <= input(14);
output(0, 90) <= input(15);
output(0, 91) <= input(16);
output(0, 92) <= input(17);
output(0, 93) <= input(18);
output(0, 94) <= input(19);
output(0, 95) <= input(20);
output(0, 96) <= input(6);
output(0, 97) <= input(7);
output(0, 98) <= input(8);
output(0, 99) <= input(9);
output(0, 100) <= input(10);
output(0, 101) <= input(11);
output(0, 102) <= input(12);
output(0, 103) <= input(13);
output(0, 104) <= input(14);
output(0, 105) <= input(15);
output(0, 106) <= input(16);
output(0, 107) <= input(17);
output(0, 108) <= input(18);
output(0, 109) <= input(19);
output(0, 110) <= input(20);
output(0, 111) <= input(21);
output(0, 112) <= input(7);
output(0, 113) <= input(8);
output(0, 114) <= input(9);
output(0, 115) <= input(10);
output(0, 116) <= input(11);
output(0, 117) <= input(12);
output(0, 118) <= input(13);
output(0, 119) <= input(14);
output(0, 120) <= input(15);
output(0, 121) <= input(16);
output(0, 122) <= input(17);
output(0, 123) <= input(18);
output(0, 124) <= input(19);
output(0, 125) <= input(20);
output(0, 126) <= input(21);
output(0, 127) <= input(22);
output(0, 128) <= input(8);
output(0, 129) <= input(9);
output(0, 130) <= input(10);
output(0, 131) <= input(11);
output(0, 132) <= input(12);
output(0, 133) <= input(13);
output(0, 134) <= input(14);
output(0, 135) <= input(15);
output(0, 136) <= input(16);
output(0, 137) <= input(17);
output(0, 138) <= input(18);
output(0, 139) <= input(19);
output(0, 140) <= input(20);
output(0, 141) <= input(21);
output(0, 142) <= input(22);
output(0, 143) <= input(23);
output(0, 144) <= input(9);
output(0, 145) <= input(10);
output(0, 146) <= input(11);
output(0, 147) <= input(12);
output(0, 148) <= input(13);
output(0, 149) <= input(14);
output(0, 150) <= input(15);
output(0, 151) <= input(16);
output(0, 152) <= input(17);
output(0, 153) <= input(18);
output(0, 154) <= input(19);
output(0, 155) <= input(20);
output(0, 156) <= input(21);
output(0, 157) <= input(22);
output(0, 158) <= input(23);
output(0, 159) <= input(24);
output(0, 160) <= input(10);
output(0, 161) <= input(11);
output(0, 162) <= input(12);
output(0, 163) <= input(13);
output(0, 164) <= input(14);
output(0, 165) <= input(15);
output(0, 166) <= input(16);
output(0, 167) <= input(17);
output(0, 168) <= input(18);
output(0, 169) <= input(19);
output(0, 170) <= input(20);
output(0, 171) <= input(21);
output(0, 172) <= input(22);
output(0, 173) <= input(23);
output(0, 174) <= input(24);
output(0, 175) <= input(25);
output(0, 176) <= input(11);
output(0, 177) <= input(12);
output(0, 178) <= input(13);
output(0, 179) <= input(14);
output(0, 180) <= input(15);
output(0, 181) <= input(16);
output(0, 182) <= input(17);
output(0, 183) <= input(18);
output(0, 184) <= input(19);
output(0, 185) <= input(20);
output(0, 186) <= input(21);
output(0, 187) <= input(22);
output(0, 188) <= input(23);
output(0, 189) <= input(24);
output(0, 190) <= input(25);
output(0, 191) <= input(26);
output(0, 192) <= input(12);
output(0, 193) <= input(13);
output(0, 194) <= input(14);
output(0, 195) <= input(15);
output(0, 196) <= input(16);
output(0, 197) <= input(17);
output(0, 198) <= input(18);
output(0, 199) <= input(19);
output(0, 200) <= input(20);
output(0, 201) <= input(21);
output(0, 202) <= input(22);
output(0, 203) <= input(23);
output(0, 204) <= input(24);
output(0, 205) <= input(25);
output(0, 206) <= input(26);
output(0, 207) <= input(27);
output(0, 208) <= input(13);
output(0, 209) <= input(14);
output(0, 210) <= input(15);
output(0, 211) <= input(16);
output(0, 212) <= input(17);
output(0, 213) <= input(18);
output(0, 214) <= input(19);
output(0, 215) <= input(20);
output(0, 216) <= input(21);
output(0, 217) <= input(22);
output(0, 218) <= input(23);
output(0, 219) <= input(24);
output(0, 220) <= input(25);
output(0, 221) <= input(26);
output(0, 222) <= input(27);
output(0, 223) <= input(28);
output(0, 224) <= input(14);
output(0, 225) <= input(15);
output(0, 226) <= input(16);
output(0, 227) <= input(17);
output(0, 228) <= input(18);
output(0, 229) <= input(19);
output(0, 230) <= input(20);
output(0, 231) <= input(21);
output(0, 232) <= input(22);
output(0, 233) <= input(23);
output(0, 234) <= input(24);
output(0, 235) <= input(25);
output(0, 236) <= input(26);
output(0, 237) <= input(27);
output(0, 238) <= input(28);
output(0, 239) <= input(29);
output(0, 240) <= input(15);
output(0, 241) <= input(16);
output(0, 242) <= input(17);
output(0, 243) <= input(18);
output(0, 244) <= input(19);
output(0, 245) <= input(20);
output(0, 246) <= input(21);
output(0, 247) <= input(22);
output(0, 248) <= input(23);
output(0, 249) <= input(24);
output(0, 250) <= input(25);
output(0, 251) <= input(26);
output(0, 252) <= input(27);
output(0, 253) <= input(28);
output(0, 254) <= input(29);
output(0, 255) <= input(30);
output(1, 0) <= input(31);
output(1, 1) <= input(32);
output(1, 2) <= input(33);
output(1, 3) <= input(34);
output(1, 4) <= input(35);
output(1, 5) <= input(36);
output(1, 6) <= input(37);
output(1, 7) <= input(38);
output(1, 8) <= input(39);
output(1, 9) <= input(40);
output(1, 10) <= input(41);
output(1, 11) <= input(42);
output(1, 12) <= input(43);
output(1, 13) <= input(44);
output(1, 14) <= input(45);
output(1, 15) <= input(46);
output(1, 16) <= input(32);
output(1, 17) <= input(33);
output(1, 18) <= input(34);
output(1, 19) <= input(35);
output(1, 20) <= input(36);
output(1, 21) <= input(37);
output(1, 22) <= input(38);
output(1, 23) <= input(39);
output(1, 24) <= input(40);
output(1, 25) <= input(41);
output(1, 26) <= input(42);
output(1, 27) <= input(43);
output(1, 28) <= input(44);
output(1, 29) <= input(45);
output(1, 30) <= input(46);
output(1, 31) <= input(47);
output(1, 32) <= input(33);
output(1, 33) <= input(34);
output(1, 34) <= input(35);
output(1, 35) <= input(36);
output(1, 36) <= input(37);
output(1, 37) <= input(38);
output(1, 38) <= input(39);
output(1, 39) <= input(40);
output(1, 40) <= input(41);
output(1, 41) <= input(42);
output(1, 42) <= input(43);
output(1, 43) <= input(44);
output(1, 44) <= input(45);
output(1, 45) <= input(46);
output(1, 46) <= input(47);
output(1, 47) <= input(48);
output(1, 48) <= input(34);
output(1, 49) <= input(35);
output(1, 50) <= input(36);
output(1, 51) <= input(37);
output(1, 52) <= input(38);
output(1, 53) <= input(39);
output(1, 54) <= input(40);
output(1, 55) <= input(41);
output(1, 56) <= input(42);
output(1, 57) <= input(43);
output(1, 58) <= input(44);
output(1, 59) <= input(45);
output(1, 60) <= input(46);
output(1, 61) <= input(47);
output(1, 62) <= input(48);
output(1, 63) <= input(49);
output(1, 64) <= input(35);
output(1, 65) <= input(36);
output(1, 66) <= input(37);
output(1, 67) <= input(38);
output(1, 68) <= input(39);
output(1, 69) <= input(40);
output(1, 70) <= input(41);
output(1, 71) <= input(42);
output(1, 72) <= input(43);
output(1, 73) <= input(44);
output(1, 74) <= input(45);
output(1, 75) <= input(46);
output(1, 76) <= input(47);
output(1, 77) <= input(48);
output(1, 78) <= input(49);
output(1, 79) <= input(50);
output(1, 80) <= input(4);
output(1, 81) <= input(5);
output(1, 82) <= input(6);
output(1, 83) <= input(7);
output(1, 84) <= input(8);
output(1, 85) <= input(9);
output(1, 86) <= input(10);
output(1, 87) <= input(11);
output(1, 88) <= input(12);
output(1, 89) <= input(13);
output(1, 90) <= input(14);
output(1, 91) <= input(15);
output(1, 92) <= input(16);
output(1, 93) <= input(17);
output(1, 94) <= input(18);
output(1, 95) <= input(19);
output(1, 96) <= input(5);
output(1, 97) <= input(6);
output(1, 98) <= input(7);
output(1, 99) <= input(8);
output(1, 100) <= input(9);
output(1, 101) <= input(10);
output(1, 102) <= input(11);
output(1, 103) <= input(12);
output(1, 104) <= input(13);
output(1, 105) <= input(14);
output(1, 106) <= input(15);
output(1, 107) <= input(16);
output(1, 108) <= input(17);
output(1, 109) <= input(18);
output(1, 110) <= input(19);
output(1, 111) <= input(20);
output(1, 112) <= input(6);
output(1, 113) <= input(7);
output(1, 114) <= input(8);
output(1, 115) <= input(9);
output(1, 116) <= input(10);
output(1, 117) <= input(11);
output(1, 118) <= input(12);
output(1, 119) <= input(13);
output(1, 120) <= input(14);
output(1, 121) <= input(15);
output(1, 122) <= input(16);
output(1, 123) <= input(17);
output(1, 124) <= input(18);
output(1, 125) <= input(19);
output(1, 126) <= input(20);
output(1, 127) <= input(21);
output(1, 128) <= input(7);
output(1, 129) <= input(8);
output(1, 130) <= input(9);
output(1, 131) <= input(10);
output(1, 132) <= input(11);
output(1, 133) <= input(12);
output(1, 134) <= input(13);
output(1, 135) <= input(14);
output(1, 136) <= input(15);
output(1, 137) <= input(16);
output(1, 138) <= input(17);
output(1, 139) <= input(18);
output(1, 140) <= input(19);
output(1, 141) <= input(20);
output(1, 142) <= input(21);
output(1, 143) <= input(22);
output(1, 144) <= input(8);
output(1, 145) <= input(9);
output(1, 146) <= input(10);
output(1, 147) <= input(11);
output(1, 148) <= input(12);
output(1, 149) <= input(13);
output(1, 150) <= input(14);
output(1, 151) <= input(15);
output(1, 152) <= input(16);
output(1, 153) <= input(17);
output(1, 154) <= input(18);
output(1, 155) <= input(19);
output(1, 156) <= input(20);
output(1, 157) <= input(21);
output(1, 158) <= input(22);
output(1, 159) <= input(23);
output(1, 160) <= input(40);
output(1, 161) <= input(41);
output(1, 162) <= input(42);
output(1, 163) <= input(43);
output(1, 164) <= input(44);
output(1, 165) <= input(45);
output(1, 166) <= input(46);
output(1, 167) <= input(47);
output(1, 168) <= input(48);
output(1, 169) <= input(49);
output(1, 170) <= input(50);
output(1, 171) <= input(51);
output(1, 172) <= input(52);
output(1, 173) <= input(53);
output(1, 174) <= input(54);
output(1, 175) <= input(55);
output(1, 176) <= input(41);
output(1, 177) <= input(42);
output(1, 178) <= input(43);
output(1, 179) <= input(44);
output(1, 180) <= input(45);
output(1, 181) <= input(46);
output(1, 182) <= input(47);
output(1, 183) <= input(48);
output(1, 184) <= input(49);
output(1, 185) <= input(50);
output(1, 186) <= input(51);
output(1, 187) <= input(52);
output(1, 188) <= input(53);
output(1, 189) <= input(54);
output(1, 190) <= input(55);
output(1, 191) <= input(56);
output(1, 192) <= input(42);
output(1, 193) <= input(43);
output(1, 194) <= input(44);
output(1, 195) <= input(45);
output(1, 196) <= input(46);
output(1, 197) <= input(47);
output(1, 198) <= input(48);
output(1, 199) <= input(49);
output(1, 200) <= input(50);
output(1, 201) <= input(51);
output(1, 202) <= input(52);
output(1, 203) <= input(53);
output(1, 204) <= input(54);
output(1, 205) <= input(55);
output(1, 206) <= input(56);
output(1, 207) <= input(57);
output(1, 208) <= input(43);
output(1, 209) <= input(44);
output(1, 210) <= input(45);
output(1, 211) <= input(46);
output(1, 212) <= input(47);
output(1, 213) <= input(48);
output(1, 214) <= input(49);
output(1, 215) <= input(50);
output(1, 216) <= input(51);
output(1, 217) <= input(52);
output(1, 218) <= input(53);
output(1, 219) <= input(54);
output(1, 220) <= input(55);
output(1, 221) <= input(56);
output(1, 222) <= input(57);
output(1, 223) <= input(58);
output(1, 224) <= input(44);
output(1, 225) <= input(45);
output(1, 226) <= input(46);
output(1, 227) <= input(47);
output(1, 228) <= input(48);
output(1, 229) <= input(49);
output(1, 230) <= input(50);
output(1, 231) <= input(51);
output(1, 232) <= input(52);
output(1, 233) <= input(53);
output(1, 234) <= input(54);
output(1, 235) <= input(55);
output(1, 236) <= input(56);
output(1, 237) <= input(57);
output(1, 238) <= input(58);
output(1, 239) <= input(59);
output(1, 240) <= input(45);
output(1, 241) <= input(46);
output(1, 242) <= input(47);
output(1, 243) <= input(48);
output(1, 244) <= input(49);
output(1, 245) <= input(50);
output(1, 246) <= input(51);
output(1, 247) <= input(52);
output(1, 248) <= input(53);
output(1, 249) <= input(54);
output(1, 250) <= input(55);
output(1, 251) <= input(56);
output(1, 252) <= input(57);
output(1, 253) <= input(58);
output(1, 254) <= input(59);
output(1, 255) <= input(60);
output(2, 0) <= input(31);
output(2, 1) <= input(32);
output(2, 2) <= input(33);
output(2, 3) <= input(34);
output(2, 4) <= input(35);
output(2, 5) <= input(36);
output(2, 6) <= input(37);
output(2, 7) <= input(38);
output(2, 8) <= input(39);
output(2, 9) <= input(40);
output(2, 10) <= input(41);
output(2, 11) <= input(42);
output(2, 12) <= input(43);
output(2, 13) <= input(44);
output(2, 14) <= input(45);
output(2, 15) <= input(46);
output(2, 16) <= input(32);
output(2, 17) <= input(33);
output(2, 18) <= input(34);
output(2, 19) <= input(35);
output(2, 20) <= input(36);
output(2, 21) <= input(37);
output(2, 22) <= input(38);
output(2, 23) <= input(39);
output(2, 24) <= input(40);
output(2, 25) <= input(41);
output(2, 26) <= input(42);
output(2, 27) <= input(43);
output(2, 28) <= input(44);
output(2, 29) <= input(45);
output(2, 30) <= input(46);
output(2, 31) <= input(47);
output(2, 32) <= input(1);
output(2, 33) <= input(2);
output(2, 34) <= input(3);
output(2, 35) <= input(4);
output(2, 36) <= input(5);
output(2, 37) <= input(6);
output(2, 38) <= input(7);
output(2, 39) <= input(8);
output(2, 40) <= input(9);
output(2, 41) <= input(10);
output(2, 42) <= input(11);
output(2, 43) <= input(12);
output(2, 44) <= input(13);
output(2, 45) <= input(14);
output(2, 46) <= input(15);
output(2, 47) <= input(16);
output(2, 48) <= input(2);
output(2, 49) <= input(3);
output(2, 50) <= input(4);
output(2, 51) <= input(5);
output(2, 52) <= input(6);
output(2, 53) <= input(7);
output(2, 54) <= input(8);
output(2, 55) <= input(9);
output(2, 56) <= input(10);
output(2, 57) <= input(11);
output(2, 58) <= input(12);
output(2, 59) <= input(13);
output(2, 60) <= input(14);
output(2, 61) <= input(15);
output(2, 62) <= input(16);
output(2, 63) <= input(17);
output(2, 64) <= input(3);
output(2, 65) <= input(4);
output(2, 66) <= input(5);
output(2, 67) <= input(6);
output(2, 68) <= input(7);
output(2, 69) <= input(8);
output(2, 70) <= input(9);
output(2, 71) <= input(10);
output(2, 72) <= input(11);
output(2, 73) <= input(12);
output(2, 74) <= input(13);
output(2, 75) <= input(14);
output(2, 76) <= input(15);
output(2, 77) <= input(16);
output(2, 78) <= input(17);
output(2, 79) <= input(18);
output(2, 80) <= input(35);
output(2, 81) <= input(36);
output(2, 82) <= input(37);
output(2, 83) <= input(38);
output(2, 84) <= input(39);
output(2, 85) <= input(40);
output(2, 86) <= input(41);
output(2, 87) <= input(42);
output(2, 88) <= input(43);
output(2, 89) <= input(44);
output(2, 90) <= input(45);
output(2, 91) <= input(46);
output(2, 92) <= input(47);
output(2, 93) <= input(48);
output(2, 94) <= input(49);
output(2, 95) <= input(50);
output(2, 96) <= input(36);
output(2, 97) <= input(37);
output(2, 98) <= input(38);
output(2, 99) <= input(39);
output(2, 100) <= input(40);
output(2, 101) <= input(41);
output(2, 102) <= input(42);
output(2, 103) <= input(43);
output(2, 104) <= input(44);
output(2, 105) <= input(45);
output(2, 106) <= input(46);
output(2, 107) <= input(47);
output(2, 108) <= input(48);
output(2, 109) <= input(49);
output(2, 110) <= input(50);
output(2, 111) <= input(51);
output(2, 112) <= input(37);
output(2, 113) <= input(38);
output(2, 114) <= input(39);
output(2, 115) <= input(40);
output(2, 116) <= input(41);
output(2, 117) <= input(42);
output(2, 118) <= input(43);
output(2, 119) <= input(44);
output(2, 120) <= input(45);
output(2, 121) <= input(46);
output(2, 122) <= input(47);
output(2, 123) <= input(48);
output(2, 124) <= input(49);
output(2, 125) <= input(50);
output(2, 126) <= input(51);
output(2, 127) <= input(52);
output(2, 128) <= input(6);
output(2, 129) <= input(7);
output(2, 130) <= input(8);
output(2, 131) <= input(9);
output(2, 132) <= input(10);
output(2, 133) <= input(11);
output(2, 134) <= input(12);
output(2, 135) <= input(13);
output(2, 136) <= input(14);
output(2, 137) <= input(15);
output(2, 138) <= input(16);
output(2, 139) <= input(17);
output(2, 140) <= input(18);
output(2, 141) <= input(19);
output(2, 142) <= input(20);
output(2, 143) <= input(21);
output(2, 144) <= input(7);
output(2, 145) <= input(8);
output(2, 146) <= input(9);
output(2, 147) <= input(10);
output(2, 148) <= input(11);
output(2, 149) <= input(12);
output(2, 150) <= input(13);
output(2, 151) <= input(14);
output(2, 152) <= input(15);
output(2, 153) <= input(16);
output(2, 154) <= input(17);
output(2, 155) <= input(18);
output(2, 156) <= input(19);
output(2, 157) <= input(20);
output(2, 158) <= input(21);
output(2, 159) <= input(22);
output(2, 160) <= input(39);
output(2, 161) <= input(40);
output(2, 162) <= input(41);
output(2, 163) <= input(42);
output(2, 164) <= input(43);
output(2, 165) <= input(44);
output(2, 166) <= input(45);
output(2, 167) <= input(46);
output(2, 168) <= input(47);
output(2, 169) <= input(48);
output(2, 170) <= input(49);
output(2, 171) <= input(50);
output(2, 172) <= input(51);
output(2, 173) <= input(52);
output(2, 174) <= input(53);
output(2, 175) <= input(54);
output(2, 176) <= input(40);
output(2, 177) <= input(41);
output(2, 178) <= input(42);
output(2, 179) <= input(43);
output(2, 180) <= input(44);
output(2, 181) <= input(45);
output(2, 182) <= input(46);
output(2, 183) <= input(47);
output(2, 184) <= input(48);
output(2, 185) <= input(49);
output(2, 186) <= input(50);
output(2, 187) <= input(51);
output(2, 188) <= input(52);
output(2, 189) <= input(53);
output(2, 190) <= input(54);
output(2, 191) <= input(55);
output(2, 192) <= input(41);
output(2, 193) <= input(42);
output(2, 194) <= input(43);
output(2, 195) <= input(44);
output(2, 196) <= input(45);
output(2, 197) <= input(46);
output(2, 198) <= input(47);
output(2, 199) <= input(48);
output(2, 200) <= input(49);
output(2, 201) <= input(50);
output(2, 202) <= input(51);
output(2, 203) <= input(52);
output(2, 204) <= input(53);
output(2, 205) <= input(54);
output(2, 206) <= input(55);
output(2, 207) <= input(56);
output(2, 208) <= input(10);
output(2, 209) <= input(11);
output(2, 210) <= input(12);
output(2, 211) <= input(13);
output(2, 212) <= input(14);
output(2, 213) <= input(15);
output(2, 214) <= input(16);
output(2, 215) <= input(17);
output(2, 216) <= input(18);
output(2, 217) <= input(19);
output(2, 218) <= input(20);
output(2, 219) <= input(21);
output(2, 220) <= input(22);
output(2, 221) <= input(23);
output(2, 222) <= input(24);
output(2, 223) <= input(25);
output(2, 224) <= input(11);
output(2, 225) <= input(12);
output(2, 226) <= input(13);
output(2, 227) <= input(14);
output(2, 228) <= input(15);
output(2, 229) <= input(16);
output(2, 230) <= input(17);
output(2, 231) <= input(18);
output(2, 232) <= input(19);
output(2, 233) <= input(20);
output(2, 234) <= input(21);
output(2, 235) <= input(22);
output(2, 236) <= input(23);
output(2, 237) <= input(24);
output(2, 238) <= input(25);
output(2, 239) <= input(26);
output(2, 240) <= input(12);
output(2, 241) <= input(13);
output(2, 242) <= input(14);
output(2, 243) <= input(15);
output(2, 244) <= input(16);
output(2, 245) <= input(17);
output(2, 246) <= input(18);
output(2, 247) <= input(19);
output(2, 248) <= input(20);
output(2, 249) <= input(21);
output(2, 250) <= input(22);
output(2, 251) <= input(23);
output(2, 252) <= input(24);
output(2, 253) <= input(25);
output(2, 254) <= input(26);
output(2, 255) <= input(27);
output(3, 0) <= input(31);
output(3, 1) <= input(32);
output(3, 2) <= input(33);
output(3, 3) <= input(34);
output(3, 4) <= input(35);
output(3, 5) <= input(36);
output(3, 6) <= input(37);
output(3, 7) <= input(38);
output(3, 8) <= input(39);
output(3, 9) <= input(40);
output(3, 10) <= input(41);
output(3, 11) <= input(42);
output(3, 12) <= input(43);
output(3, 13) <= input(44);
output(3, 14) <= input(45);
output(3, 15) <= input(46);
output(3, 16) <= input(0);
output(3, 17) <= input(1);
output(3, 18) <= input(2);
output(3, 19) <= input(3);
output(3, 20) <= input(4);
output(3, 21) <= input(5);
output(3, 22) <= input(6);
output(3, 23) <= input(7);
output(3, 24) <= input(8);
output(3, 25) <= input(9);
output(3, 26) <= input(10);
output(3, 27) <= input(11);
output(3, 28) <= input(12);
output(3, 29) <= input(13);
output(3, 30) <= input(14);
output(3, 31) <= input(15);
output(3, 32) <= input(1);
output(3, 33) <= input(2);
output(3, 34) <= input(3);
output(3, 35) <= input(4);
output(3, 36) <= input(5);
output(3, 37) <= input(6);
output(3, 38) <= input(7);
output(3, 39) <= input(8);
output(3, 40) <= input(9);
output(3, 41) <= input(10);
output(3, 42) <= input(11);
output(3, 43) <= input(12);
output(3, 44) <= input(13);
output(3, 45) <= input(14);
output(3, 46) <= input(15);
output(3, 47) <= input(16);
output(3, 48) <= input(33);
output(3, 49) <= input(34);
output(3, 50) <= input(35);
output(3, 51) <= input(36);
output(3, 52) <= input(37);
output(3, 53) <= input(38);
output(3, 54) <= input(39);
output(3, 55) <= input(40);
output(3, 56) <= input(41);
output(3, 57) <= input(42);
output(3, 58) <= input(43);
output(3, 59) <= input(44);
output(3, 60) <= input(45);
output(3, 61) <= input(46);
output(3, 62) <= input(47);
output(3, 63) <= input(48);
output(3, 64) <= input(34);
output(3, 65) <= input(35);
output(3, 66) <= input(36);
output(3, 67) <= input(37);
output(3, 68) <= input(38);
output(3, 69) <= input(39);
output(3, 70) <= input(40);
output(3, 71) <= input(41);
output(3, 72) <= input(42);
output(3, 73) <= input(43);
output(3, 74) <= input(44);
output(3, 75) <= input(45);
output(3, 76) <= input(46);
output(3, 77) <= input(47);
output(3, 78) <= input(48);
output(3, 79) <= input(49);
output(3, 80) <= input(3);
output(3, 81) <= input(4);
output(3, 82) <= input(5);
output(3, 83) <= input(6);
output(3, 84) <= input(7);
output(3, 85) <= input(8);
output(3, 86) <= input(9);
output(3, 87) <= input(10);
output(3, 88) <= input(11);
output(3, 89) <= input(12);
output(3, 90) <= input(13);
output(3, 91) <= input(14);
output(3, 92) <= input(15);
output(3, 93) <= input(16);
output(3, 94) <= input(17);
output(3, 95) <= input(18);
output(3, 96) <= input(4);
output(3, 97) <= input(5);
output(3, 98) <= input(6);
output(3, 99) <= input(7);
output(3, 100) <= input(8);
output(3, 101) <= input(9);
output(3, 102) <= input(10);
output(3, 103) <= input(11);
output(3, 104) <= input(12);
output(3, 105) <= input(13);
output(3, 106) <= input(14);
output(3, 107) <= input(15);
output(3, 108) <= input(16);
output(3, 109) <= input(17);
output(3, 110) <= input(18);
output(3, 111) <= input(19);
output(3, 112) <= input(36);
output(3, 113) <= input(37);
output(3, 114) <= input(38);
output(3, 115) <= input(39);
output(3, 116) <= input(40);
output(3, 117) <= input(41);
output(3, 118) <= input(42);
output(3, 119) <= input(43);
output(3, 120) <= input(44);
output(3, 121) <= input(45);
output(3, 122) <= input(46);
output(3, 123) <= input(47);
output(3, 124) <= input(48);
output(3, 125) <= input(49);
output(3, 126) <= input(50);
output(3, 127) <= input(51);
output(3, 128) <= input(5);
output(3, 129) <= input(6);
output(3, 130) <= input(7);
output(3, 131) <= input(8);
output(3, 132) <= input(9);
output(3, 133) <= input(10);
output(3, 134) <= input(11);
output(3, 135) <= input(12);
output(3, 136) <= input(13);
output(3, 137) <= input(14);
output(3, 138) <= input(15);
output(3, 139) <= input(16);
output(3, 140) <= input(17);
output(3, 141) <= input(18);
output(3, 142) <= input(19);
output(3, 143) <= input(20);
output(3, 144) <= input(6);
output(3, 145) <= input(7);
output(3, 146) <= input(8);
output(3, 147) <= input(9);
output(3, 148) <= input(10);
output(3, 149) <= input(11);
output(3, 150) <= input(12);
output(3, 151) <= input(13);
output(3, 152) <= input(14);
output(3, 153) <= input(15);
output(3, 154) <= input(16);
output(3, 155) <= input(17);
output(3, 156) <= input(18);
output(3, 157) <= input(19);
output(3, 158) <= input(20);
output(3, 159) <= input(21);
output(3, 160) <= input(38);
output(3, 161) <= input(39);
output(3, 162) <= input(40);
output(3, 163) <= input(41);
output(3, 164) <= input(42);
output(3, 165) <= input(43);
output(3, 166) <= input(44);
output(3, 167) <= input(45);
output(3, 168) <= input(46);
output(3, 169) <= input(47);
output(3, 170) <= input(48);
output(3, 171) <= input(49);
output(3, 172) <= input(50);
output(3, 173) <= input(51);
output(3, 174) <= input(52);
output(3, 175) <= input(53);
output(3, 176) <= input(39);
output(3, 177) <= input(40);
output(3, 178) <= input(41);
output(3, 179) <= input(42);
output(3, 180) <= input(43);
output(3, 181) <= input(44);
output(3, 182) <= input(45);
output(3, 183) <= input(46);
output(3, 184) <= input(47);
output(3, 185) <= input(48);
output(3, 186) <= input(49);
output(3, 187) <= input(50);
output(3, 188) <= input(51);
output(3, 189) <= input(52);
output(3, 190) <= input(53);
output(3, 191) <= input(54);
output(3, 192) <= input(8);
output(3, 193) <= input(9);
output(3, 194) <= input(10);
output(3, 195) <= input(11);
output(3, 196) <= input(12);
output(3, 197) <= input(13);
output(3, 198) <= input(14);
output(3, 199) <= input(15);
output(3, 200) <= input(16);
output(3, 201) <= input(17);
output(3, 202) <= input(18);
output(3, 203) <= input(19);
output(3, 204) <= input(20);
output(3, 205) <= input(21);
output(3, 206) <= input(22);
output(3, 207) <= input(23);
output(3, 208) <= input(9);
output(3, 209) <= input(10);
output(3, 210) <= input(11);
output(3, 211) <= input(12);
output(3, 212) <= input(13);
output(3, 213) <= input(14);
output(3, 214) <= input(15);
output(3, 215) <= input(16);
output(3, 216) <= input(17);
output(3, 217) <= input(18);
output(3, 218) <= input(19);
output(3, 219) <= input(20);
output(3, 220) <= input(21);
output(3, 221) <= input(22);
output(3, 222) <= input(23);
output(3, 223) <= input(24);
output(3, 224) <= input(41);
output(3, 225) <= input(42);
output(3, 226) <= input(43);
output(3, 227) <= input(44);
output(3, 228) <= input(45);
output(3, 229) <= input(46);
output(3, 230) <= input(47);
output(3, 231) <= input(48);
output(3, 232) <= input(49);
output(3, 233) <= input(50);
output(3, 234) <= input(51);
output(3, 235) <= input(52);
output(3, 236) <= input(53);
output(3, 237) <= input(54);
output(3, 238) <= input(55);
output(3, 239) <= input(56);
output(3, 240) <= input(42);
output(3, 241) <= input(43);
output(3, 242) <= input(44);
output(3, 243) <= input(45);
output(3, 244) <= input(46);
output(3, 245) <= input(47);
output(3, 246) <= input(48);
output(3, 247) <= input(49);
output(3, 248) <= input(50);
output(3, 249) <= input(51);
output(3, 250) <= input(52);
output(3, 251) <= input(53);
output(3, 252) <= input(54);
output(3, 253) <= input(55);
output(3, 254) <= input(56);
output(3, 255) <= input(57);
output(4, 0) <= input(31);
output(4, 1) <= input(32);
output(4, 2) <= input(33);
output(4, 3) <= input(34);
output(4, 4) <= input(35);
output(4, 5) <= input(36);
output(4, 6) <= input(37);
output(4, 7) <= input(38);
output(4, 8) <= input(39);
output(4, 9) <= input(40);
output(4, 10) <= input(41);
output(4, 11) <= input(42);
output(4, 12) <= input(43);
output(4, 13) <= input(44);
output(4, 14) <= input(45);
output(4, 15) <= input(46);
output(4, 16) <= input(0);
output(4, 17) <= input(1);
output(4, 18) <= input(2);
output(4, 19) <= input(3);
output(4, 20) <= input(4);
output(4, 21) <= input(5);
output(4, 22) <= input(6);
output(4, 23) <= input(7);
output(4, 24) <= input(8);
output(4, 25) <= input(9);
output(4, 26) <= input(10);
output(4, 27) <= input(11);
output(4, 28) <= input(12);
output(4, 29) <= input(13);
output(4, 30) <= input(14);
output(4, 31) <= input(15);
output(4, 32) <= input(32);
output(4, 33) <= input(33);
output(4, 34) <= input(34);
output(4, 35) <= input(35);
output(4, 36) <= input(36);
output(4, 37) <= input(37);
output(4, 38) <= input(38);
output(4, 39) <= input(39);
output(4, 40) <= input(40);
output(4, 41) <= input(41);
output(4, 42) <= input(42);
output(4, 43) <= input(43);
output(4, 44) <= input(44);
output(4, 45) <= input(45);
output(4, 46) <= input(46);
output(4, 47) <= input(47);
output(4, 48) <= input(33);
output(4, 49) <= input(34);
output(4, 50) <= input(35);
output(4, 51) <= input(36);
output(4, 52) <= input(37);
output(4, 53) <= input(38);
output(4, 54) <= input(39);
output(4, 55) <= input(40);
output(4, 56) <= input(41);
output(4, 57) <= input(42);
output(4, 58) <= input(43);
output(4, 59) <= input(44);
output(4, 60) <= input(45);
output(4, 61) <= input(46);
output(4, 62) <= input(47);
output(4, 63) <= input(48);
output(4, 64) <= input(2);
output(4, 65) <= input(3);
output(4, 66) <= input(4);
output(4, 67) <= input(5);
output(4, 68) <= input(6);
output(4, 69) <= input(7);
output(4, 70) <= input(8);
output(4, 71) <= input(9);
output(4, 72) <= input(10);
output(4, 73) <= input(11);
output(4, 74) <= input(12);
output(4, 75) <= input(13);
output(4, 76) <= input(14);
output(4, 77) <= input(15);
output(4, 78) <= input(16);
output(4, 79) <= input(17);
output(4, 80) <= input(34);
output(4, 81) <= input(35);
output(4, 82) <= input(36);
output(4, 83) <= input(37);
output(4, 84) <= input(38);
output(4, 85) <= input(39);
output(4, 86) <= input(40);
output(4, 87) <= input(41);
output(4, 88) <= input(42);
output(4, 89) <= input(43);
output(4, 90) <= input(44);
output(4, 91) <= input(45);
output(4, 92) <= input(46);
output(4, 93) <= input(47);
output(4, 94) <= input(48);
output(4, 95) <= input(49);
output(4, 96) <= input(3);
output(4, 97) <= input(4);
output(4, 98) <= input(5);
output(4, 99) <= input(6);
output(4, 100) <= input(7);
output(4, 101) <= input(8);
output(4, 102) <= input(9);
output(4, 103) <= input(10);
output(4, 104) <= input(11);
output(4, 105) <= input(12);
output(4, 106) <= input(13);
output(4, 107) <= input(14);
output(4, 108) <= input(15);
output(4, 109) <= input(16);
output(4, 110) <= input(17);
output(4, 111) <= input(18);
output(4, 112) <= input(4);
output(4, 113) <= input(5);
output(4, 114) <= input(6);
output(4, 115) <= input(7);
output(4, 116) <= input(8);
output(4, 117) <= input(9);
output(4, 118) <= input(10);
output(4, 119) <= input(11);
output(4, 120) <= input(12);
output(4, 121) <= input(13);
output(4, 122) <= input(14);
output(4, 123) <= input(15);
output(4, 124) <= input(16);
output(4, 125) <= input(17);
output(4, 126) <= input(18);
output(4, 127) <= input(19);
output(4, 128) <= input(36);
output(4, 129) <= input(37);
output(4, 130) <= input(38);
output(4, 131) <= input(39);
output(4, 132) <= input(40);
output(4, 133) <= input(41);
output(4, 134) <= input(42);
output(4, 135) <= input(43);
output(4, 136) <= input(44);
output(4, 137) <= input(45);
output(4, 138) <= input(46);
output(4, 139) <= input(47);
output(4, 140) <= input(48);
output(4, 141) <= input(49);
output(4, 142) <= input(50);
output(4, 143) <= input(51);
output(4, 144) <= input(5);
output(4, 145) <= input(6);
output(4, 146) <= input(7);
output(4, 147) <= input(8);
output(4, 148) <= input(9);
output(4, 149) <= input(10);
output(4, 150) <= input(11);
output(4, 151) <= input(12);
output(4, 152) <= input(13);
output(4, 153) <= input(14);
output(4, 154) <= input(15);
output(4, 155) <= input(16);
output(4, 156) <= input(17);
output(4, 157) <= input(18);
output(4, 158) <= input(19);
output(4, 159) <= input(20);
output(4, 160) <= input(37);
output(4, 161) <= input(38);
output(4, 162) <= input(39);
output(4, 163) <= input(40);
output(4, 164) <= input(41);
output(4, 165) <= input(42);
output(4, 166) <= input(43);
output(4, 167) <= input(44);
output(4, 168) <= input(45);
output(4, 169) <= input(46);
output(4, 170) <= input(47);
output(4, 171) <= input(48);
output(4, 172) <= input(49);
output(4, 173) <= input(50);
output(4, 174) <= input(51);
output(4, 175) <= input(52);
output(4, 176) <= input(38);
output(4, 177) <= input(39);
output(4, 178) <= input(40);
output(4, 179) <= input(41);
output(4, 180) <= input(42);
output(4, 181) <= input(43);
output(4, 182) <= input(44);
output(4, 183) <= input(45);
output(4, 184) <= input(46);
output(4, 185) <= input(47);
output(4, 186) <= input(48);
output(4, 187) <= input(49);
output(4, 188) <= input(50);
output(4, 189) <= input(51);
output(4, 190) <= input(52);
output(4, 191) <= input(53);
output(4, 192) <= input(7);
output(4, 193) <= input(8);
output(4, 194) <= input(9);
output(4, 195) <= input(10);
output(4, 196) <= input(11);
output(4, 197) <= input(12);
output(4, 198) <= input(13);
output(4, 199) <= input(14);
output(4, 200) <= input(15);
output(4, 201) <= input(16);
output(4, 202) <= input(17);
output(4, 203) <= input(18);
output(4, 204) <= input(19);
output(4, 205) <= input(20);
output(4, 206) <= input(21);
output(4, 207) <= input(22);
output(4, 208) <= input(39);
output(4, 209) <= input(40);
output(4, 210) <= input(41);
output(4, 211) <= input(42);
output(4, 212) <= input(43);
output(4, 213) <= input(44);
output(4, 214) <= input(45);
output(4, 215) <= input(46);
output(4, 216) <= input(47);
output(4, 217) <= input(48);
output(4, 218) <= input(49);
output(4, 219) <= input(50);
output(4, 220) <= input(51);
output(4, 221) <= input(52);
output(4, 222) <= input(53);
output(4, 223) <= input(54);
output(4, 224) <= input(8);
output(4, 225) <= input(9);
output(4, 226) <= input(10);
output(4, 227) <= input(11);
output(4, 228) <= input(12);
output(4, 229) <= input(13);
output(4, 230) <= input(14);
output(4, 231) <= input(15);
output(4, 232) <= input(16);
output(4, 233) <= input(17);
output(4, 234) <= input(18);
output(4, 235) <= input(19);
output(4, 236) <= input(20);
output(4, 237) <= input(21);
output(4, 238) <= input(22);
output(4, 239) <= input(23);
output(4, 240) <= input(9);
output(4, 241) <= input(10);
output(4, 242) <= input(11);
output(4, 243) <= input(12);
output(4, 244) <= input(13);
output(4, 245) <= input(14);
output(4, 246) <= input(15);
output(4, 247) <= input(16);
output(4, 248) <= input(17);
output(4, 249) <= input(18);
output(4, 250) <= input(19);
output(4, 251) <= input(20);
output(4, 252) <= input(21);
output(4, 253) <= input(22);
output(4, 254) <= input(23);
output(4, 255) <= input(24);
output(5, 0) <= input(31);
output(5, 1) <= input(32);
output(5, 2) <= input(33);
output(5, 3) <= input(34);
output(5, 4) <= input(35);
output(5, 5) <= input(36);
output(5, 6) <= input(37);
output(5, 7) <= input(38);
output(5, 8) <= input(39);
output(5, 9) <= input(40);
output(5, 10) <= input(41);
output(5, 11) <= input(42);
output(5, 12) <= input(43);
output(5, 13) <= input(44);
output(5, 14) <= input(45);
output(5, 15) <= input(46);
output(5, 16) <= input(0);
output(5, 17) <= input(1);
output(5, 18) <= input(2);
output(5, 19) <= input(3);
output(5, 20) <= input(4);
output(5, 21) <= input(5);
output(5, 22) <= input(6);
output(5, 23) <= input(7);
output(5, 24) <= input(8);
output(5, 25) <= input(9);
output(5, 26) <= input(10);
output(5, 27) <= input(11);
output(5, 28) <= input(12);
output(5, 29) <= input(13);
output(5, 30) <= input(14);
output(5, 31) <= input(15);
output(5, 32) <= input(32);
output(5, 33) <= input(33);
output(5, 34) <= input(34);
output(5, 35) <= input(35);
output(5, 36) <= input(36);
output(5, 37) <= input(37);
output(5, 38) <= input(38);
output(5, 39) <= input(39);
output(5, 40) <= input(40);
output(5, 41) <= input(41);
output(5, 42) <= input(42);
output(5, 43) <= input(43);
output(5, 44) <= input(44);
output(5, 45) <= input(45);
output(5, 46) <= input(46);
output(5, 47) <= input(47);
output(5, 48) <= input(1);
output(5, 49) <= input(2);
output(5, 50) <= input(3);
output(5, 51) <= input(4);
output(5, 52) <= input(5);
output(5, 53) <= input(6);
output(5, 54) <= input(7);
output(5, 55) <= input(8);
output(5, 56) <= input(9);
output(5, 57) <= input(10);
output(5, 58) <= input(11);
output(5, 59) <= input(12);
output(5, 60) <= input(13);
output(5, 61) <= input(14);
output(5, 62) <= input(15);
output(5, 63) <= input(16);
output(5, 64) <= input(33);
output(5, 65) <= input(34);
output(5, 66) <= input(35);
output(5, 67) <= input(36);
output(5, 68) <= input(37);
output(5, 69) <= input(38);
output(5, 70) <= input(39);
output(5, 71) <= input(40);
output(5, 72) <= input(41);
output(5, 73) <= input(42);
output(5, 74) <= input(43);
output(5, 75) <= input(44);
output(5, 76) <= input(45);
output(5, 77) <= input(46);
output(5, 78) <= input(47);
output(5, 79) <= input(48);
output(5, 80) <= input(2);
output(5, 81) <= input(3);
output(5, 82) <= input(4);
output(5, 83) <= input(5);
output(5, 84) <= input(6);
output(5, 85) <= input(7);
output(5, 86) <= input(8);
output(5, 87) <= input(9);
output(5, 88) <= input(10);
output(5, 89) <= input(11);
output(5, 90) <= input(12);
output(5, 91) <= input(13);
output(5, 92) <= input(14);
output(5, 93) <= input(15);
output(5, 94) <= input(16);
output(5, 95) <= input(17);
output(5, 96) <= input(34);
output(5, 97) <= input(35);
output(5, 98) <= input(36);
output(5, 99) <= input(37);
output(5, 100) <= input(38);
output(5, 101) <= input(39);
output(5, 102) <= input(40);
output(5, 103) <= input(41);
output(5, 104) <= input(42);
output(5, 105) <= input(43);
output(5, 106) <= input(44);
output(5, 107) <= input(45);
output(5, 108) <= input(46);
output(5, 109) <= input(47);
output(5, 110) <= input(48);
output(5, 111) <= input(49);
output(5, 112) <= input(35);
output(5, 113) <= input(36);
output(5, 114) <= input(37);
output(5, 115) <= input(38);
output(5, 116) <= input(39);
output(5, 117) <= input(40);
output(5, 118) <= input(41);
output(5, 119) <= input(42);
output(5, 120) <= input(43);
output(5, 121) <= input(44);
output(5, 122) <= input(45);
output(5, 123) <= input(46);
output(5, 124) <= input(47);
output(5, 125) <= input(48);
output(5, 126) <= input(49);
output(5, 127) <= input(50);
output(5, 128) <= input(4);
output(5, 129) <= input(5);
output(5, 130) <= input(6);
output(5, 131) <= input(7);
output(5, 132) <= input(8);
output(5, 133) <= input(9);
output(5, 134) <= input(10);
output(5, 135) <= input(11);
output(5, 136) <= input(12);
output(5, 137) <= input(13);
output(5, 138) <= input(14);
output(5, 139) <= input(15);
output(5, 140) <= input(16);
output(5, 141) <= input(17);
output(5, 142) <= input(18);
output(5, 143) <= input(19);
output(5, 144) <= input(36);
output(5, 145) <= input(37);
output(5, 146) <= input(38);
output(5, 147) <= input(39);
output(5, 148) <= input(40);
output(5, 149) <= input(41);
output(5, 150) <= input(42);
output(5, 151) <= input(43);
output(5, 152) <= input(44);
output(5, 153) <= input(45);
output(5, 154) <= input(46);
output(5, 155) <= input(47);
output(5, 156) <= input(48);
output(5, 157) <= input(49);
output(5, 158) <= input(50);
output(5, 159) <= input(51);
output(5, 160) <= input(5);
output(5, 161) <= input(6);
output(5, 162) <= input(7);
output(5, 163) <= input(8);
output(5, 164) <= input(9);
output(5, 165) <= input(10);
output(5, 166) <= input(11);
output(5, 167) <= input(12);
output(5, 168) <= input(13);
output(5, 169) <= input(14);
output(5, 170) <= input(15);
output(5, 171) <= input(16);
output(5, 172) <= input(17);
output(5, 173) <= input(18);
output(5, 174) <= input(19);
output(5, 175) <= input(20);
output(5, 176) <= input(37);
output(5, 177) <= input(38);
output(5, 178) <= input(39);
output(5, 179) <= input(40);
output(5, 180) <= input(41);
output(5, 181) <= input(42);
output(5, 182) <= input(43);
output(5, 183) <= input(44);
output(5, 184) <= input(45);
output(5, 185) <= input(46);
output(5, 186) <= input(47);
output(5, 187) <= input(48);
output(5, 188) <= input(49);
output(5, 189) <= input(50);
output(5, 190) <= input(51);
output(5, 191) <= input(52);
output(5, 192) <= input(6);
output(5, 193) <= input(7);
output(5, 194) <= input(8);
output(5, 195) <= input(9);
output(5, 196) <= input(10);
output(5, 197) <= input(11);
output(5, 198) <= input(12);
output(5, 199) <= input(13);
output(5, 200) <= input(14);
output(5, 201) <= input(15);
output(5, 202) <= input(16);
output(5, 203) <= input(17);
output(5, 204) <= input(18);
output(5, 205) <= input(19);
output(5, 206) <= input(20);
output(5, 207) <= input(21);
output(5, 208) <= input(38);
output(5, 209) <= input(39);
output(5, 210) <= input(40);
output(5, 211) <= input(41);
output(5, 212) <= input(42);
output(5, 213) <= input(43);
output(5, 214) <= input(44);
output(5, 215) <= input(45);
output(5, 216) <= input(46);
output(5, 217) <= input(47);
output(5, 218) <= input(48);
output(5, 219) <= input(49);
output(5, 220) <= input(50);
output(5, 221) <= input(51);
output(5, 222) <= input(52);
output(5, 223) <= input(53);
output(5, 224) <= input(7);
output(5, 225) <= input(8);
output(5, 226) <= input(9);
output(5, 227) <= input(10);
output(5, 228) <= input(11);
output(5, 229) <= input(12);
output(5, 230) <= input(13);
output(5, 231) <= input(14);
output(5, 232) <= input(15);
output(5, 233) <= input(16);
output(5, 234) <= input(17);
output(5, 235) <= input(18);
output(5, 236) <= input(19);
output(5, 237) <= input(20);
output(5, 238) <= input(21);
output(5, 239) <= input(22);
output(5, 240) <= input(8);
output(5, 241) <= input(9);
output(5, 242) <= input(10);
output(5, 243) <= input(11);
output(5, 244) <= input(12);
output(5, 245) <= input(13);
output(5, 246) <= input(14);
output(5, 247) <= input(15);
output(5, 248) <= input(16);
output(5, 249) <= input(17);
output(5, 250) <= input(18);
output(5, 251) <= input(19);
output(5, 252) <= input(20);
output(5, 253) <= input(21);
output(5, 254) <= input(22);
output(5, 255) <= input(23);
when "0001" =>
output(0, 0) <= input(0);
output(0, 1) <= input(1);
output(0, 2) <= input(2);
output(0, 3) <= input(3);
output(0, 4) <= input(4);
output(0, 5) <= input(5);
output(0, 6) <= input(6);
output(0, 7) <= input(7);
output(0, 8) <= input(8);
output(0, 9) <= input(9);
output(0, 10) <= input(10);
output(0, 11) <= input(11);
output(0, 12) <= input(12);
output(0, 13) <= input(13);
output(0, 14) <= input(14);
output(0, 15) <= input(15);
output(0, 16) <= input(16);
output(0, 17) <= input(17);
output(0, 18) <= input(18);
output(0, 19) <= input(19);
output(0, 20) <= input(20);
output(0, 21) <= input(21);
output(0, 22) <= input(22);
output(0, 23) <= input(23);
output(0, 24) <= input(24);
output(0, 25) <= input(25);
output(0, 26) <= input(26);
output(0, 27) <= input(27);
output(0, 28) <= input(28);
output(0, 29) <= input(29);
output(0, 30) <= input(30);
output(0, 31) <= input(31);
output(0, 32) <= input(1);
output(0, 33) <= input(2);
output(0, 34) <= input(3);
output(0, 35) <= input(4);
output(0, 36) <= input(5);
output(0, 37) <= input(6);
output(0, 38) <= input(7);
output(0, 39) <= input(8);
output(0, 40) <= input(9);
output(0, 41) <= input(10);
output(0, 42) <= input(11);
output(0, 43) <= input(12);
output(0, 44) <= input(13);
output(0, 45) <= input(14);
output(0, 46) <= input(15);
output(0, 47) <= input(32);
output(0, 48) <= input(17);
output(0, 49) <= input(18);
output(0, 50) <= input(19);
output(0, 51) <= input(20);
output(0, 52) <= input(21);
output(0, 53) <= input(22);
output(0, 54) <= input(23);
output(0, 55) <= input(24);
output(0, 56) <= input(25);
output(0, 57) <= input(26);
output(0, 58) <= input(27);
output(0, 59) <= input(28);
output(0, 60) <= input(29);
output(0, 61) <= input(30);
output(0, 62) <= input(31);
output(0, 63) <= input(33);
output(0, 64) <= input(2);
output(0, 65) <= input(3);
output(0, 66) <= input(4);
output(0, 67) <= input(5);
output(0, 68) <= input(6);
output(0, 69) <= input(7);
output(0, 70) <= input(8);
output(0, 71) <= input(9);
output(0, 72) <= input(10);
output(0, 73) <= input(11);
output(0, 74) <= input(12);
output(0, 75) <= input(13);
output(0, 76) <= input(14);
output(0, 77) <= input(15);
output(0, 78) <= input(32);
output(0, 79) <= input(34);
output(0, 80) <= input(18);
output(0, 81) <= input(19);
output(0, 82) <= input(20);
output(0, 83) <= input(21);
output(0, 84) <= input(22);
output(0, 85) <= input(23);
output(0, 86) <= input(24);
output(0, 87) <= input(25);
output(0, 88) <= input(26);
output(0, 89) <= input(27);
output(0, 90) <= input(28);
output(0, 91) <= input(29);
output(0, 92) <= input(30);
output(0, 93) <= input(31);
output(0, 94) <= input(33);
output(0, 95) <= input(35);
output(0, 96) <= input(3);
output(0, 97) <= input(4);
output(0, 98) <= input(5);
output(0, 99) <= input(6);
output(0, 100) <= input(7);
output(0, 101) <= input(8);
output(0, 102) <= input(9);
output(0, 103) <= input(10);
output(0, 104) <= input(11);
output(0, 105) <= input(12);
output(0, 106) <= input(13);
output(0, 107) <= input(14);
output(0, 108) <= input(15);
output(0, 109) <= input(32);
output(0, 110) <= input(34);
output(0, 111) <= input(36);
output(0, 112) <= input(19);
output(0, 113) <= input(20);
output(0, 114) <= input(21);
output(0, 115) <= input(22);
output(0, 116) <= input(23);
output(0, 117) <= input(24);
output(0, 118) <= input(25);
output(0, 119) <= input(26);
output(0, 120) <= input(27);
output(0, 121) <= input(28);
output(0, 122) <= input(29);
output(0, 123) <= input(30);
output(0, 124) <= input(31);
output(0, 125) <= input(33);
output(0, 126) <= input(35);
output(0, 127) <= input(37);
output(0, 128) <= input(4);
output(0, 129) <= input(5);
output(0, 130) <= input(6);
output(0, 131) <= input(7);
output(0, 132) <= input(8);
output(0, 133) <= input(9);
output(0, 134) <= input(10);
output(0, 135) <= input(11);
output(0, 136) <= input(12);
output(0, 137) <= input(13);
output(0, 138) <= input(14);
output(0, 139) <= input(15);
output(0, 140) <= input(32);
output(0, 141) <= input(34);
output(0, 142) <= input(36);
output(0, 143) <= input(38);
output(0, 144) <= input(20);
output(0, 145) <= input(21);
output(0, 146) <= input(22);
output(0, 147) <= input(23);
output(0, 148) <= input(24);
output(0, 149) <= input(25);
output(0, 150) <= input(26);
output(0, 151) <= input(27);
output(0, 152) <= input(28);
output(0, 153) <= input(29);
output(0, 154) <= input(30);
output(0, 155) <= input(31);
output(0, 156) <= input(33);
output(0, 157) <= input(35);
output(0, 158) <= input(37);
output(0, 159) <= input(39);
output(0, 160) <= input(5);
output(0, 161) <= input(6);
output(0, 162) <= input(7);
output(0, 163) <= input(8);
output(0, 164) <= input(9);
output(0, 165) <= input(10);
output(0, 166) <= input(11);
output(0, 167) <= input(12);
output(0, 168) <= input(13);
output(0, 169) <= input(14);
output(0, 170) <= input(15);
output(0, 171) <= input(32);
output(0, 172) <= input(34);
output(0, 173) <= input(36);
output(0, 174) <= input(38);
output(0, 175) <= input(40);
output(0, 176) <= input(21);
output(0, 177) <= input(22);
output(0, 178) <= input(23);
output(0, 179) <= input(24);
output(0, 180) <= input(25);
output(0, 181) <= input(26);
output(0, 182) <= input(27);
output(0, 183) <= input(28);
output(0, 184) <= input(29);
output(0, 185) <= input(30);
output(0, 186) <= input(31);
output(0, 187) <= input(33);
output(0, 188) <= input(35);
output(0, 189) <= input(37);
output(0, 190) <= input(39);
output(0, 191) <= input(41);
output(0, 192) <= input(6);
output(0, 193) <= input(7);
output(0, 194) <= input(8);
output(0, 195) <= input(9);
output(0, 196) <= input(10);
output(0, 197) <= input(11);
output(0, 198) <= input(12);
output(0, 199) <= input(13);
output(0, 200) <= input(14);
output(0, 201) <= input(15);
output(0, 202) <= input(32);
output(0, 203) <= input(34);
output(0, 204) <= input(36);
output(0, 205) <= input(38);
output(0, 206) <= input(40);
output(0, 207) <= input(42);
output(0, 208) <= input(22);
output(0, 209) <= input(23);
output(0, 210) <= input(24);
output(0, 211) <= input(25);
output(0, 212) <= input(26);
output(0, 213) <= input(27);
output(0, 214) <= input(28);
output(0, 215) <= input(29);
output(0, 216) <= input(30);
output(0, 217) <= input(31);
output(0, 218) <= input(33);
output(0, 219) <= input(35);
output(0, 220) <= input(37);
output(0, 221) <= input(39);
output(0, 222) <= input(41);
output(0, 223) <= input(43);
output(0, 224) <= input(7);
output(0, 225) <= input(8);
output(0, 226) <= input(9);
output(0, 227) <= input(10);
output(0, 228) <= input(11);
output(0, 229) <= input(12);
output(0, 230) <= input(13);
output(0, 231) <= input(14);
output(0, 232) <= input(15);
output(0, 233) <= input(32);
output(0, 234) <= input(34);
output(0, 235) <= input(36);
output(0, 236) <= input(38);
output(0, 237) <= input(40);
output(0, 238) <= input(42);
output(0, 239) <= input(44);
output(0, 240) <= input(23);
output(0, 241) <= input(24);
output(0, 242) <= input(25);
output(0, 243) <= input(26);
output(0, 244) <= input(27);
output(0, 245) <= input(28);
output(0, 246) <= input(29);
output(0, 247) <= input(30);
output(0, 248) <= input(31);
output(0, 249) <= input(33);
output(0, 250) <= input(35);
output(0, 251) <= input(37);
output(0, 252) <= input(39);
output(0, 253) <= input(41);
output(0, 254) <= input(43);
output(0, 255) <= input(45);
output(1, 0) <= input(46);
output(1, 1) <= input(16);
output(1, 2) <= input(17);
output(1, 3) <= input(18);
output(1, 4) <= input(19);
output(1, 5) <= input(20);
output(1, 6) <= input(21);
output(1, 7) <= input(22);
output(1, 8) <= input(23);
output(1, 9) <= input(24);
output(1, 10) <= input(25);
output(1, 11) <= input(26);
output(1, 12) <= input(27);
output(1, 13) <= input(28);
output(1, 14) <= input(29);
output(1, 15) <= input(30);
output(1, 16) <= input(0);
output(1, 17) <= input(1);
output(1, 18) <= input(2);
output(1, 19) <= input(3);
output(1, 20) <= input(4);
output(1, 21) <= input(5);
output(1, 22) <= input(6);
output(1, 23) <= input(7);
output(1, 24) <= input(8);
output(1, 25) <= input(9);
output(1, 26) <= input(10);
output(1, 27) <= input(11);
output(1, 28) <= input(12);
output(1, 29) <= input(13);
output(1, 30) <= input(14);
output(1, 31) <= input(15);
output(1, 32) <= input(16);
output(1, 33) <= input(17);
output(1, 34) <= input(18);
output(1, 35) <= input(19);
output(1, 36) <= input(20);
output(1, 37) <= input(21);
output(1, 38) <= input(22);
output(1, 39) <= input(23);
output(1, 40) <= input(24);
output(1, 41) <= input(25);
output(1, 42) <= input(26);
output(1, 43) <= input(27);
output(1, 44) <= input(28);
output(1, 45) <= input(29);
output(1, 46) <= input(30);
output(1, 47) <= input(31);
output(1, 48) <= input(1);
output(1, 49) <= input(2);
output(1, 50) <= input(3);
output(1, 51) <= input(4);
output(1, 52) <= input(5);
output(1, 53) <= input(6);
output(1, 54) <= input(7);
output(1, 55) <= input(8);
output(1, 56) <= input(9);
output(1, 57) <= input(10);
output(1, 58) <= input(11);
output(1, 59) <= input(12);
output(1, 60) <= input(13);
output(1, 61) <= input(14);
output(1, 62) <= input(15);
output(1, 63) <= input(32);
output(1, 64) <= input(17);
output(1, 65) <= input(18);
output(1, 66) <= input(19);
output(1, 67) <= input(20);
output(1, 68) <= input(21);
output(1, 69) <= input(22);
output(1, 70) <= input(23);
output(1, 71) <= input(24);
output(1, 72) <= input(25);
output(1, 73) <= input(26);
output(1, 74) <= input(27);
output(1, 75) <= input(28);
output(1, 76) <= input(29);
output(1, 77) <= input(30);
output(1, 78) <= input(31);
output(1, 79) <= input(33);
output(1, 80) <= input(2);
output(1, 81) <= input(3);
output(1, 82) <= input(4);
output(1, 83) <= input(5);
output(1, 84) <= input(6);
output(1, 85) <= input(7);
output(1, 86) <= input(8);
output(1, 87) <= input(9);
output(1, 88) <= input(10);
output(1, 89) <= input(11);
output(1, 90) <= input(12);
output(1, 91) <= input(13);
output(1, 92) <= input(14);
output(1, 93) <= input(15);
output(1, 94) <= input(32);
output(1, 95) <= input(34);
output(1, 96) <= input(18);
output(1, 97) <= input(19);
output(1, 98) <= input(20);
output(1, 99) <= input(21);
output(1, 100) <= input(22);
output(1, 101) <= input(23);
output(1, 102) <= input(24);
output(1, 103) <= input(25);
output(1, 104) <= input(26);
output(1, 105) <= input(27);
output(1, 106) <= input(28);
output(1, 107) <= input(29);
output(1, 108) <= input(30);
output(1, 109) <= input(31);
output(1, 110) <= input(33);
output(1, 111) <= input(35);
output(1, 112) <= input(3);
output(1, 113) <= input(4);
output(1, 114) <= input(5);
output(1, 115) <= input(6);
output(1, 116) <= input(7);
output(1, 117) <= input(8);
output(1, 118) <= input(9);
output(1, 119) <= input(10);
output(1, 120) <= input(11);
output(1, 121) <= input(12);
output(1, 122) <= input(13);
output(1, 123) <= input(14);
output(1, 124) <= input(15);
output(1, 125) <= input(32);
output(1, 126) <= input(34);
output(1, 127) <= input(36);
output(1, 128) <= input(3);
output(1, 129) <= input(4);
output(1, 130) <= input(5);
output(1, 131) <= input(6);
output(1, 132) <= input(7);
output(1, 133) <= input(8);
output(1, 134) <= input(9);
output(1, 135) <= input(10);
output(1, 136) <= input(11);
output(1, 137) <= input(12);
output(1, 138) <= input(13);
output(1, 139) <= input(14);
output(1, 140) <= input(15);
output(1, 141) <= input(32);
output(1, 142) <= input(34);
output(1, 143) <= input(36);
output(1, 144) <= input(19);
output(1, 145) <= input(20);
output(1, 146) <= input(21);
output(1, 147) <= input(22);
output(1, 148) <= input(23);
output(1, 149) <= input(24);
output(1, 150) <= input(25);
output(1, 151) <= input(26);
output(1, 152) <= input(27);
output(1, 153) <= input(28);
output(1, 154) <= input(29);
output(1, 155) <= input(30);
output(1, 156) <= input(31);
output(1, 157) <= input(33);
output(1, 158) <= input(35);
output(1, 159) <= input(37);
output(1, 160) <= input(4);
output(1, 161) <= input(5);
output(1, 162) <= input(6);
output(1, 163) <= input(7);
output(1, 164) <= input(8);
output(1, 165) <= input(9);
output(1, 166) <= input(10);
output(1, 167) <= input(11);
output(1, 168) <= input(12);
output(1, 169) <= input(13);
output(1, 170) <= input(14);
output(1, 171) <= input(15);
output(1, 172) <= input(32);
output(1, 173) <= input(34);
output(1, 174) <= input(36);
output(1, 175) <= input(38);
output(1, 176) <= input(20);
output(1, 177) <= input(21);
output(1, 178) <= input(22);
output(1, 179) <= input(23);
output(1, 180) <= input(24);
output(1, 181) <= input(25);
output(1, 182) <= input(26);
output(1, 183) <= input(27);
output(1, 184) <= input(28);
output(1, 185) <= input(29);
output(1, 186) <= input(30);
output(1, 187) <= input(31);
output(1, 188) <= input(33);
output(1, 189) <= input(35);
output(1, 190) <= input(37);
output(1, 191) <= input(39);
output(1, 192) <= input(5);
output(1, 193) <= input(6);
output(1, 194) <= input(7);
output(1, 195) <= input(8);
output(1, 196) <= input(9);
output(1, 197) <= input(10);
output(1, 198) <= input(11);
output(1, 199) <= input(12);
output(1, 200) <= input(13);
output(1, 201) <= input(14);
output(1, 202) <= input(15);
output(1, 203) <= input(32);
output(1, 204) <= input(34);
output(1, 205) <= input(36);
output(1, 206) <= input(38);
output(1, 207) <= input(40);
output(1, 208) <= input(21);
output(1, 209) <= input(22);
output(1, 210) <= input(23);
output(1, 211) <= input(24);
output(1, 212) <= input(25);
output(1, 213) <= input(26);
output(1, 214) <= input(27);
output(1, 215) <= input(28);
output(1, 216) <= input(29);
output(1, 217) <= input(30);
output(1, 218) <= input(31);
output(1, 219) <= input(33);
output(1, 220) <= input(35);
output(1, 221) <= input(37);
output(1, 222) <= input(39);
output(1, 223) <= input(41);
output(1, 224) <= input(6);
output(1, 225) <= input(7);
output(1, 226) <= input(8);
output(1, 227) <= input(9);
output(1, 228) <= input(10);
output(1, 229) <= input(11);
output(1, 230) <= input(12);
output(1, 231) <= input(13);
output(1, 232) <= input(14);
output(1, 233) <= input(15);
output(1, 234) <= input(32);
output(1, 235) <= input(34);
output(1, 236) <= input(36);
output(1, 237) <= input(38);
output(1, 238) <= input(40);
output(1, 239) <= input(42);
output(1, 240) <= input(22);
output(1, 241) <= input(23);
output(1, 242) <= input(24);
output(1, 243) <= input(25);
output(1, 244) <= input(26);
output(1, 245) <= input(27);
output(1, 246) <= input(28);
output(1, 247) <= input(29);
output(1, 248) <= input(30);
output(1, 249) <= input(31);
output(1, 250) <= input(33);
output(1, 251) <= input(35);
output(1, 252) <= input(37);
output(1, 253) <= input(39);
output(1, 254) <= input(41);
output(1, 255) <= input(43);
output(2, 0) <= input(46);
output(2, 1) <= input(16);
output(2, 2) <= input(17);
output(2, 3) <= input(18);
output(2, 4) <= input(19);
output(2, 5) <= input(20);
output(2, 6) <= input(21);
output(2, 7) <= input(22);
output(2, 8) <= input(23);
output(2, 9) <= input(24);
output(2, 10) <= input(25);
output(2, 11) <= input(26);
output(2, 12) <= input(27);
output(2, 13) <= input(28);
output(2, 14) <= input(29);
output(2, 15) <= input(30);
output(2, 16) <= input(0);
output(2, 17) <= input(1);
output(2, 18) <= input(2);
output(2, 19) <= input(3);
output(2, 20) <= input(4);
output(2, 21) <= input(5);
output(2, 22) <= input(6);
output(2, 23) <= input(7);
output(2, 24) <= input(8);
output(2, 25) <= input(9);
output(2, 26) <= input(10);
output(2, 27) <= input(11);
output(2, 28) <= input(12);
output(2, 29) <= input(13);
output(2, 30) <= input(14);
output(2, 31) <= input(15);
output(2, 32) <= input(16);
output(2, 33) <= input(17);
output(2, 34) <= input(18);
output(2, 35) <= input(19);
output(2, 36) <= input(20);
output(2, 37) <= input(21);
output(2, 38) <= input(22);
output(2, 39) <= input(23);
output(2, 40) <= input(24);
output(2, 41) <= input(25);
output(2, 42) <= input(26);
output(2, 43) <= input(27);
output(2, 44) <= input(28);
output(2, 45) <= input(29);
output(2, 46) <= input(30);
output(2, 47) <= input(31);
output(2, 48) <= input(1);
output(2, 49) <= input(2);
output(2, 50) <= input(3);
output(2, 51) <= input(4);
output(2, 52) <= input(5);
output(2, 53) <= input(6);
output(2, 54) <= input(7);
output(2, 55) <= input(8);
output(2, 56) <= input(9);
output(2, 57) <= input(10);
output(2, 58) <= input(11);
output(2, 59) <= input(12);
output(2, 60) <= input(13);
output(2, 61) <= input(14);
output(2, 62) <= input(15);
output(2, 63) <= input(32);
output(2, 64) <= input(1);
output(2, 65) <= input(2);
output(2, 66) <= input(3);
output(2, 67) <= input(4);
output(2, 68) <= input(5);
output(2, 69) <= input(6);
output(2, 70) <= input(7);
output(2, 71) <= input(8);
output(2, 72) <= input(9);
output(2, 73) <= input(10);
output(2, 74) <= input(11);
output(2, 75) <= input(12);
output(2, 76) <= input(13);
output(2, 77) <= input(14);
output(2, 78) <= input(15);
output(2, 79) <= input(32);
output(2, 80) <= input(17);
output(2, 81) <= input(18);
output(2, 82) <= input(19);
output(2, 83) <= input(20);
output(2, 84) <= input(21);
output(2, 85) <= input(22);
output(2, 86) <= input(23);
output(2, 87) <= input(24);
output(2, 88) <= input(25);
output(2, 89) <= input(26);
output(2, 90) <= input(27);
output(2, 91) <= input(28);
output(2, 92) <= input(29);
output(2, 93) <= input(30);
output(2, 94) <= input(31);
output(2, 95) <= input(33);
output(2, 96) <= input(2);
output(2, 97) <= input(3);
output(2, 98) <= input(4);
output(2, 99) <= input(5);
output(2, 100) <= input(6);
output(2, 101) <= input(7);
output(2, 102) <= input(8);
output(2, 103) <= input(9);
output(2, 104) <= input(10);
output(2, 105) <= input(11);
output(2, 106) <= input(12);
output(2, 107) <= input(13);
output(2, 108) <= input(14);
output(2, 109) <= input(15);
output(2, 110) <= input(32);
output(2, 111) <= input(34);
output(2, 112) <= input(18);
output(2, 113) <= input(19);
output(2, 114) <= input(20);
output(2, 115) <= input(21);
output(2, 116) <= input(22);
output(2, 117) <= input(23);
output(2, 118) <= input(24);
output(2, 119) <= input(25);
output(2, 120) <= input(26);
output(2, 121) <= input(27);
output(2, 122) <= input(28);
output(2, 123) <= input(29);
output(2, 124) <= input(30);
output(2, 125) <= input(31);
output(2, 126) <= input(33);
output(2, 127) <= input(35);
output(2, 128) <= input(18);
output(2, 129) <= input(19);
output(2, 130) <= input(20);
output(2, 131) <= input(21);
output(2, 132) <= input(22);
output(2, 133) <= input(23);
output(2, 134) <= input(24);
output(2, 135) <= input(25);
output(2, 136) <= input(26);
output(2, 137) <= input(27);
output(2, 138) <= input(28);
output(2, 139) <= input(29);
output(2, 140) <= input(30);
output(2, 141) <= input(31);
output(2, 142) <= input(33);
output(2, 143) <= input(35);
output(2, 144) <= input(3);
output(2, 145) <= input(4);
output(2, 146) <= input(5);
output(2, 147) <= input(6);
output(2, 148) <= input(7);
output(2, 149) <= input(8);
output(2, 150) <= input(9);
output(2, 151) <= input(10);
output(2, 152) <= input(11);
output(2, 153) <= input(12);
output(2, 154) <= input(13);
output(2, 155) <= input(14);
output(2, 156) <= input(15);
output(2, 157) <= input(32);
output(2, 158) <= input(34);
output(2, 159) <= input(36);
output(2, 160) <= input(19);
output(2, 161) <= input(20);
output(2, 162) <= input(21);
output(2, 163) <= input(22);
output(2, 164) <= input(23);
output(2, 165) <= input(24);
output(2, 166) <= input(25);
output(2, 167) <= input(26);
output(2, 168) <= input(27);
output(2, 169) <= input(28);
output(2, 170) <= input(29);
output(2, 171) <= input(30);
output(2, 172) <= input(31);
output(2, 173) <= input(33);
output(2, 174) <= input(35);
output(2, 175) <= input(37);
output(2, 176) <= input(4);
output(2, 177) <= input(5);
output(2, 178) <= input(6);
output(2, 179) <= input(7);
output(2, 180) <= input(8);
output(2, 181) <= input(9);
output(2, 182) <= input(10);
output(2, 183) <= input(11);
output(2, 184) <= input(12);
output(2, 185) <= input(13);
output(2, 186) <= input(14);
output(2, 187) <= input(15);
output(2, 188) <= input(32);
output(2, 189) <= input(34);
output(2, 190) <= input(36);
output(2, 191) <= input(38);
output(2, 192) <= input(4);
output(2, 193) <= input(5);
output(2, 194) <= input(6);
output(2, 195) <= input(7);
output(2, 196) <= input(8);
output(2, 197) <= input(9);
output(2, 198) <= input(10);
output(2, 199) <= input(11);
output(2, 200) <= input(12);
output(2, 201) <= input(13);
output(2, 202) <= input(14);
output(2, 203) <= input(15);
output(2, 204) <= input(32);
output(2, 205) <= input(34);
output(2, 206) <= input(36);
output(2, 207) <= input(38);
output(2, 208) <= input(20);
output(2, 209) <= input(21);
output(2, 210) <= input(22);
output(2, 211) <= input(23);
output(2, 212) <= input(24);
output(2, 213) <= input(25);
output(2, 214) <= input(26);
output(2, 215) <= input(27);
output(2, 216) <= input(28);
output(2, 217) <= input(29);
output(2, 218) <= input(30);
output(2, 219) <= input(31);
output(2, 220) <= input(33);
output(2, 221) <= input(35);
output(2, 222) <= input(37);
output(2, 223) <= input(39);
output(2, 224) <= input(5);
output(2, 225) <= input(6);
output(2, 226) <= input(7);
output(2, 227) <= input(8);
output(2, 228) <= input(9);
output(2, 229) <= input(10);
output(2, 230) <= input(11);
output(2, 231) <= input(12);
output(2, 232) <= input(13);
output(2, 233) <= input(14);
output(2, 234) <= input(15);
output(2, 235) <= input(32);
output(2, 236) <= input(34);
output(2, 237) <= input(36);
output(2, 238) <= input(38);
output(2, 239) <= input(40);
output(2, 240) <= input(21);
output(2, 241) <= input(22);
output(2, 242) <= input(23);
output(2, 243) <= input(24);
output(2, 244) <= input(25);
output(2, 245) <= input(26);
output(2, 246) <= input(27);
output(2, 247) <= input(28);
output(2, 248) <= input(29);
output(2, 249) <= input(30);
output(2, 250) <= input(31);
output(2, 251) <= input(33);
output(2, 252) <= input(35);
output(2, 253) <= input(37);
output(2, 254) <= input(39);
output(2, 255) <= input(41);
output(3, 0) <= input(46);
output(3, 1) <= input(16);
output(3, 2) <= input(17);
output(3, 3) <= input(18);
output(3, 4) <= input(19);
output(3, 5) <= input(20);
output(3, 6) <= input(21);
output(3, 7) <= input(22);
output(3, 8) <= input(23);
output(3, 9) <= input(24);
output(3, 10) <= input(25);
output(3, 11) <= input(26);
output(3, 12) <= input(27);
output(3, 13) <= input(28);
output(3, 14) <= input(29);
output(3, 15) <= input(30);
output(3, 16) <= input(0);
output(3, 17) <= input(1);
output(3, 18) <= input(2);
output(3, 19) <= input(3);
output(3, 20) <= input(4);
output(3, 21) <= input(5);
output(3, 22) <= input(6);
output(3, 23) <= input(7);
output(3, 24) <= input(8);
output(3, 25) <= input(9);
output(3, 26) <= input(10);
output(3, 27) <= input(11);
output(3, 28) <= input(12);
output(3, 29) <= input(13);
output(3, 30) <= input(14);
output(3, 31) <= input(15);
output(3, 32) <= input(0);
output(3, 33) <= input(1);
output(3, 34) <= input(2);
output(3, 35) <= input(3);
output(3, 36) <= input(4);
output(3, 37) <= input(5);
output(3, 38) <= input(6);
output(3, 39) <= input(7);
output(3, 40) <= input(8);
output(3, 41) <= input(9);
output(3, 42) <= input(10);
output(3, 43) <= input(11);
output(3, 44) <= input(12);
output(3, 45) <= input(13);
output(3, 46) <= input(14);
output(3, 47) <= input(15);
output(3, 48) <= input(16);
output(3, 49) <= input(17);
output(3, 50) <= input(18);
output(3, 51) <= input(19);
output(3, 52) <= input(20);
output(3, 53) <= input(21);
output(3, 54) <= input(22);
output(3, 55) <= input(23);
output(3, 56) <= input(24);
output(3, 57) <= input(25);
output(3, 58) <= input(26);
output(3, 59) <= input(27);
output(3, 60) <= input(28);
output(3, 61) <= input(29);
output(3, 62) <= input(30);
output(3, 63) <= input(31);
output(3, 64) <= input(1);
output(3, 65) <= input(2);
output(3, 66) <= input(3);
output(3, 67) <= input(4);
output(3, 68) <= input(5);
output(3, 69) <= input(6);
output(3, 70) <= input(7);
output(3, 71) <= input(8);
output(3, 72) <= input(9);
output(3, 73) <= input(10);
output(3, 74) <= input(11);
output(3, 75) <= input(12);
output(3, 76) <= input(13);
output(3, 77) <= input(14);
output(3, 78) <= input(15);
output(3, 79) <= input(32);
output(3, 80) <= input(1);
output(3, 81) <= input(2);
output(3, 82) <= input(3);
output(3, 83) <= input(4);
output(3, 84) <= input(5);
output(3, 85) <= input(6);
output(3, 86) <= input(7);
output(3, 87) <= input(8);
output(3, 88) <= input(9);
output(3, 89) <= input(10);
output(3, 90) <= input(11);
output(3, 91) <= input(12);
output(3, 92) <= input(13);
output(3, 93) <= input(14);
output(3, 94) <= input(15);
output(3, 95) <= input(32);
output(3, 96) <= input(17);
output(3, 97) <= input(18);
output(3, 98) <= input(19);
output(3, 99) <= input(20);
output(3, 100) <= input(21);
output(3, 101) <= input(22);
output(3, 102) <= input(23);
output(3, 103) <= input(24);
output(3, 104) <= input(25);
output(3, 105) <= input(26);
output(3, 106) <= input(27);
output(3, 107) <= input(28);
output(3, 108) <= input(29);
output(3, 109) <= input(30);
output(3, 110) <= input(31);
output(3, 111) <= input(33);
output(3, 112) <= input(2);
output(3, 113) <= input(3);
output(3, 114) <= input(4);
output(3, 115) <= input(5);
output(3, 116) <= input(6);
output(3, 117) <= input(7);
output(3, 118) <= input(8);
output(3, 119) <= input(9);
output(3, 120) <= input(10);
output(3, 121) <= input(11);
output(3, 122) <= input(12);
output(3, 123) <= input(13);
output(3, 124) <= input(14);
output(3, 125) <= input(15);
output(3, 126) <= input(32);
output(3, 127) <= input(34);
output(3, 128) <= input(2);
output(3, 129) <= input(3);
output(3, 130) <= input(4);
output(3, 131) <= input(5);
output(3, 132) <= input(6);
output(3, 133) <= input(7);
output(3, 134) <= input(8);
output(3, 135) <= input(9);
output(3, 136) <= input(10);
output(3, 137) <= input(11);
output(3, 138) <= input(12);
output(3, 139) <= input(13);
output(3, 140) <= input(14);
output(3, 141) <= input(15);
output(3, 142) <= input(32);
output(3, 143) <= input(34);
output(3, 144) <= input(18);
output(3, 145) <= input(19);
output(3, 146) <= input(20);
output(3, 147) <= input(21);
output(3, 148) <= input(22);
output(3, 149) <= input(23);
output(3, 150) <= input(24);
output(3, 151) <= input(25);
output(3, 152) <= input(26);
output(3, 153) <= input(27);
output(3, 154) <= input(28);
output(3, 155) <= input(29);
output(3, 156) <= input(30);
output(3, 157) <= input(31);
output(3, 158) <= input(33);
output(3, 159) <= input(35);
output(3, 160) <= input(18);
output(3, 161) <= input(19);
output(3, 162) <= input(20);
output(3, 163) <= input(21);
output(3, 164) <= input(22);
output(3, 165) <= input(23);
output(3, 166) <= input(24);
output(3, 167) <= input(25);
output(3, 168) <= input(26);
output(3, 169) <= input(27);
output(3, 170) <= input(28);
output(3, 171) <= input(29);
output(3, 172) <= input(30);
output(3, 173) <= input(31);
output(3, 174) <= input(33);
output(3, 175) <= input(35);
output(3, 176) <= input(3);
output(3, 177) <= input(4);
output(3, 178) <= input(5);
output(3, 179) <= input(6);
output(3, 180) <= input(7);
output(3, 181) <= input(8);
output(3, 182) <= input(9);
output(3, 183) <= input(10);
output(3, 184) <= input(11);
output(3, 185) <= input(12);
output(3, 186) <= input(13);
output(3, 187) <= input(14);
output(3, 188) <= input(15);
output(3, 189) <= input(32);
output(3, 190) <= input(34);
output(3, 191) <= input(36);
output(3, 192) <= input(19);
output(3, 193) <= input(20);
output(3, 194) <= input(21);
output(3, 195) <= input(22);
output(3, 196) <= input(23);
output(3, 197) <= input(24);
output(3, 198) <= input(25);
output(3, 199) <= input(26);
output(3, 200) <= input(27);
output(3, 201) <= input(28);
output(3, 202) <= input(29);
output(3, 203) <= input(30);
output(3, 204) <= input(31);
output(3, 205) <= input(33);
output(3, 206) <= input(35);
output(3, 207) <= input(37);
output(3, 208) <= input(19);
output(3, 209) <= input(20);
output(3, 210) <= input(21);
output(3, 211) <= input(22);
output(3, 212) <= input(23);
output(3, 213) <= input(24);
output(3, 214) <= input(25);
output(3, 215) <= input(26);
output(3, 216) <= input(27);
output(3, 217) <= input(28);
output(3, 218) <= input(29);
output(3, 219) <= input(30);
output(3, 220) <= input(31);
output(3, 221) <= input(33);
output(3, 222) <= input(35);
output(3, 223) <= input(37);
output(3, 224) <= input(4);
output(3, 225) <= input(5);
output(3, 226) <= input(6);
output(3, 227) <= input(7);
output(3, 228) <= input(8);
output(3, 229) <= input(9);
output(3, 230) <= input(10);
output(3, 231) <= input(11);
output(3, 232) <= input(12);
output(3, 233) <= input(13);
output(3, 234) <= input(14);
output(3, 235) <= input(15);
output(3, 236) <= input(32);
output(3, 237) <= input(34);
output(3, 238) <= input(36);
output(3, 239) <= input(38);
output(3, 240) <= input(20);
output(3, 241) <= input(21);
output(3, 242) <= input(22);
output(3, 243) <= input(23);
output(3, 244) <= input(24);
output(3, 245) <= input(25);
output(3, 246) <= input(26);
output(3, 247) <= input(27);
output(3, 248) <= input(28);
output(3, 249) <= input(29);
output(3, 250) <= input(30);
output(3, 251) <= input(31);
output(3, 252) <= input(33);
output(3, 253) <= input(35);
output(3, 254) <= input(37);
output(3, 255) <= input(39);
output(4, 0) <= input(46);
output(4, 1) <= input(16);
output(4, 2) <= input(17);
output(4, 3) <= input(18);
output(4, 4) <= input(19);
output(4, 5) <= input(20);
output(4, 6) <= input(21);
output(4, 7) <= input(22);
output(4, 8) <= input(23);
output(4, 9) <= input(24);
output(4, 10) <= input(25);
output(4, 11) <= input(26);
output(4, 12) <= input(27);
output(4, 13) <= input(28);
output(4, 14) <= input(29);
output(4, 15) <= input(30);
output(4, 16) <= input(0);
output(4, 17) <= input(1);
output(4, 18) <= input(2);
output(4, 19) <= input(3);
output(4, 20) <= input(4);
output(4, 21) <= input(5);
output(4, 22) <= input(6);
output(4, 23) <= input(7);
output(4, 24) <= input(8);
output(4, 25) <= input(9);
output(4, 26) <= input(10);
output(4, 27) <= input(11);
output(4, 28) <= input(12);
output(4, 29) <= input(13);
output(4, 30) <= input(14);
output(4, 31) <= input(15);
output(4, 32) <= input(0);
output(4, 33) <= input(1);
output(4, 34) <= input(2);
output(4, 35) <= input(3);
output(4, 36) <= input(4);
output(4, 37) <= input(5);
output(4, 38) <= input(6);
output(4, 39) <= input(7);
output(4, 40) <= input(8);
output(4, 41) <= input(9);
output(4, 42) <= input(10);
output(4, 43) <= input(11);
output(4, 44) <= input(12);
output(4, 45) <= input(13);
output(4, 46) <= input(14);
output(4, 47) <= input(15);
output(4, 48) <= input(16);
output(4, 49) <= input(17);
output(4, 50) <= input(18);
output(4, 51) <= input(19);
output(4, 52) <= input(20);
output(4, 53) <= input(21);
output(4, 54) <= input(22);
output(4, 55) <= input(23);
output(4, 56) <= input(24);
output(4, 57) <= input(25);
output(4, 58) <= input(26);
output(4, 59) <= input(27);
output(4, 60) <= input(28);
output(4, 61) <= input(29);
output(4, 62) <= input(30);
output(4, 63) <= input(31);
output(4, 64) <= input(16);
output(4, 65) <= input(17);
output(4, 66) <= input(18);
output(4, 67) <= input(19);
output(4, 68) <= input(20);
output(4, 69) <= input(21);
output(4, 70) <= input(22);
output(4, 71) <= input(23);
output(4, 72) <= input(24);
output(4, 73) <= input(25);
output(4, 74) <= input(26);
output(4, 75) <= input(27);
output(4, 76) <= input(28);
output(4, 77) <= input(29);
output(4, 78) <= input(30);
output(4, 79) <= input(31);
output(4, 80) <= input(1);
output(4, 81) <= input(2);
output(4, 82) <= input(3);
output(4, 83) <= input(4);
output(4, 84) <= input(5);
output(4, 85) <= input(6);
output(4, 86) <= input(7);
output(4, 87) <= input(8);
output(4, 88) <= input(9);
output(4, 89) <= input(10);
output(4, 90) <= input(11);
output(4, 91) <= input(12);
output(4, 92) <= input(13);
output(4, 93) <= input(14);
output(4, 94) <= input(15);
output(4, 95) <= input(32);
output(4, 96) <= input(1);
output(4, 97) <= input(2);
output(4, 98) <= input(3);
output(4, 99) <= input(4);
output(4, 100) <= input(5);
output(4, 101) <= input(6);
output(4, 102) <= input(7);
output(4, 103) <= input(8);
output(4, 104) <= input(9);
output(4, 105) <= input(10);
output(4, 106) <= input(11);
output(4, 107) <= input(12);
output(4, 108) <= input(13);
output(4, 109) <= input(14);
output(4, 110) <= input(15);
output(4, 111) <= input(32);
output(4, 112) <= input(17);
output(4, 113) <= input(18);
output(4, 114) <= input(19);
output(4, 115) <= input(20);
output(4, 116) <= input(21);
output(4, 117) <= input(22);
output(4, 118) <= input(23);
output(4, 119) <= input(24);
output(4, 120) <= input(25);
output(4, 121) <= input(26);
output(4, 122) <= input(27);
output(4, 123) <= input(28);
output(4, 124) <= input(29);
output(4, 125) <= input(30);
output(4, 126) <= input(31);
output(4, 127) <= input(33);
output(4, 128) <= input(17);
output(4, 129) <= input(18);
output(4, 130) <= input(19);
output(4, 131) <= input(20);
output(4, 132) <= input(21);
output(4, 133) <= input(22);
output(4, 134) <= input(23);
output(4, 135) <= input(24);
output(4, 136) <= input(25);
output(4, 137) <= input(26);
output(4, 138) <= input(27);
output(4, 139) <= input(28);
output(4, 140) <= input(29);
output(4, 141) <= input(30);
output(4, 142) <= input(31);
output(4, 143) <= input(33);
output(4, 144) <= input(2);
output(4, 145) <= input(3);
output(4, 146) <= input(4);
output(4, 147) <= input(5);
output(4, 148) <= input(6);
output(4, 149) <= input(7);
output(4, 150) <= input(8);
output(4, 151) <= input(9);
output(4, 152) <= input(10);
output(4, 153) <= input(11);
output(4, 154) <= input(12);
output(4, 155) <= input(13);
output(4, 156) <= input(14);
output(4, 157) <= input(15);
output(4, 158) <= input(32);
output(4, 159) <= input(34);
output(4, 160) <= input(2);
output(4, 161) <= input(3);
output(4, 162) <= input(4);
output(4, 163) <= input(5);
output(4, 164) <= input(6);
output(4, 165) <= input(7);
output(4, 166) <= input(8);
output(4, 167) <= input(9);
output(4, 168) <= input(10);
output(4, 169) <= input(11);
output(4, 170) <= input(12);
output(4, 171) <= input(13);
output(4, 172) <= input(14);
output(4, 173) <= input(15);
output(4, 174) <= input(32);
output(4, 175) <= input(34);
output(4, 176) <= input(18);
output(4, 177) <= input(19);
output(4, 178) <= input(20);
output(4, 179) <= input(21);
output(4, 180) <= input(22);
output(4, 181) <= input(23);
output(4, 182) <= input(24);
output(4, 183) <= input(25);
output(4, 184) <= input(26);
output(4, 185) <= input(27);
output(4, 186) <= input(28);
output(4, 187) <= input(29);
output(4, 188) <= input(30);
output(4, 189) <= input(31);
output(4, 190) <= input(33);
output(4, 191) <= input(35);
output(4, 192) <= input(18);
output(4, 193) <= input(19);
output(4, 194) <= input(20);
output(4, 195) <= input(21);
output(4, 196) <= input(22);
output(4, 197) <= input(23);
output(4, 198) <= input(24);
output(4, 199) <= input(25);
output(4, 200) <= input(26);
output(4, 201) <= input(27);
output(4, 202) <= input(28);
output(4, 203) <= input(29);
output(4, 204) <= input(30);
output(4, 205) <= input(31);
output(4, 206) <= input(33);
output(4, 207) <= input(35);
output(4, 208) <= input(3);
output(4, 209) <= input(4);
output(4, 210) <= input(5);
output(4, 211) <= input(6);
output(4, 212) <= input(7);
output(4, 213) <= input(8);
output(4, 214) <= input(9);
output(4, 215) <= input(10);
output(4, 216) <= input(11);
output(4, 217) <= input(12);
output(4, 218) <= input(13);
output(4, 219) <= input(14);
output(4, 220) <= input(15);
output(4, 221) <= input(32);
output(4, 222) <= input(34);
output(4, 223) <= input(36);
output(4, 224) <= input(3);
output(4, 225) <= input(4);
output(4, 226) <= input(5);
output(4, 227) <= input(6);
output(4, 228) <= input(7);
output(4, 229) <= input(8);
output(4, 230) <= input(9);
output(4, 231) <= input(10);
output(4, 232) <= input(11);
output(4, 233) <= input(12);
output(4, 234) <= input(13);
output(4, 235) <= input(14);
output(4, 236) <= input(15);
output(4, 237) <= input(32);
output(4, 238) <= input(34);
output(4, 239) <= input(36);
output(4, 240) <= input(19);
output(4, 241) <= input(20);
output(4, 242) <= input(21);
output(4, 243) <= input(22);
output(4, 244) <= input(23);
output(4, 245) <= input(24);
output(4, 246) <= input(25);
output(4, 247) <= input(26);
output(4, 248) <= input(27);
output(4, 249) <= input(28);
output(4, 250) <= input(29);
output(4, 251) <= input(30);
output(4, 252) <= input(31);
output(4, 253) <= input(33);
output(4, 254) <= input(35);
output(4, 255) <= input(37);
output(5, 0) <= input(46);
output(5, 1) <= input(16);
output(5, 2) <= input(17);
output(5, 3) <= input(18);
output(5, 4) <= input(19);
output(5, 5) <= input(20);
output(5, 6) <= input(21);
output(5, 7) <= input(22);
output(5, 8) <= input(23);
output(5, 9) <= input(24);
output(5, 10) <= input(25);
output(5, 11) <= input(26);
output(5, 12) <= input(27);
output(5, 13) <= input(28);
output(5, 14) <= input(29);
output(5, 15) <= input(30);
output(5, 16) <= input(46);
output(5, 17) <= input(16);
output(5, 18) <= input(17);
output(5, 19) <= input(18);
output(5, 20) <= input(19);
output(5, 21) <= input(20);
output(5, 22) <= input(21);
output(5, 23) <= input(22);
output(5, 24) <= input(23);
output(5, 25) <= input(24);
output(5, 26) <= input(25);
output(5, 27) <= input(26);
output(5, 28) <= input(27);
output(5, 29) <= input(28);
output(5, 30) <= input(29);
output(5, 31) <= input(30);
output(5, 32) <= input(0);
output(5, 33) <= input(1);
output(5, 34) <= input(2);
output(5, 35) <= input(3);
output(5, 36) <= input(4);
output(5, 37) <= input(5);
output(5, 38) <= input(6);
output(5, 39) <= input(7);
output(5, 40) <= input(8);
output(5, 41) <= input(9);
output(5, 42) <= input(10);
output(5, 43) <= input(11);
output(5, 44) <= input(12);
output(5, 45) <= input(13);
output(5, 46) <= input(14);
output(5, 47) <= input(15);
output(5, 48) <= input(0);
output(5, 49) <= input(1);
output(5, 50) <= input(2);
output(5, 51) <= input(3);
output(5, 52) <= input(4);
output(5, 53) <= input(5);
output(5, 54) <= input(6);
output(5, 55) <= input(7);
output(5, 56) <= input(8);
output(5, 57) <= input(9);
output(5, 58) <= input(10);
output(5, 59) <= input(11);
output(5, 60) <= input(12);
output(5, 61) <= input(13);
output(5, 62) <= input(14);
output(5, 63) <= input(15);
output(5, 64) <= input(0);
output(5, 65) <= input(1);
output(5, 66) <= input(2);
output(5, 67) <= input(3);
output(5, 68) <= input(4);
output(5, 69) <= input(5);
output(5, 70) <= input(6);
output(5, 71) <= input(7);
output(5, 72) <= input(8);
output(5, 73) <= input(9);
output(5, 74) <= input(10);
output(5, 75) <= input(11);
output(5, 76) <= input(12);
output(5, 77) <= input(13);
output(5, 78) <= input(14);
output(5, 79) <= input(15);
output(5, 80) <= input(16);
output(5, 81) <= input(17);
output(5, 82) <= input(18);
output(5, 83) <= input(19);
output(5, 84) <= input(20);
output(5, 85) <= input(21);
output(5, 86) <= input(22);
output(5, 87) <= input(23);
output(5, 88) <= input(24);
output(5, 89) <= input(25);
output(5, 90) <= input(26);
output(5, 91) <= input(27);
output(5, 92) <= input(28);
output(5, 93) <= input(29);
output(5, 94) <= input(30);
output(5, 95) <= input(31);
output(5, 96) <= input(16);
output(5, 97) <= input(17);
output(5, 98) <= input(18);
output(5, 99) <= input(19);
output(5, 100) <= input(20);
output(5, 101) <= input(21);
output(5, 102) <= input(22);
output(5, 103) <= input(23);
output(5, 104) <= input(24);
output(5, 105) <= input(25);
output(5, 106) <= input(26);
output(5, 107) <= input(27);
output(5, 108) <= input(28);
output(5, 109) <= input(29);
output(5, 110) <= input(30);
output(5, 111) <= input(31);
output(5, 112) <= input(1);
output(5, 113) <= input(2);
output(5, 114) <= input(3);
output(5, 115) <= input(4);
output(5, 116) <= input(5);
output(5, 117) <= input(6);
output(5, 118) <= input(7);
output(5, 119) <= input(8);
output(5, 120) <= input(9);
output(5, 121) <= input(10);
output(5, 122) <= input(11);
output(5, 123) <= input(12);
output(5, 124) <= input(13);
output(5, 125) <= input(14);
output(5, 126) <= input(15);
output(5, 127) <= input(32);
output(5, 128) <= input(1);
output(5, 129) <= input(2);
output(5, 130) <= input(3);
output(5, 131) <= input(4);
output(5, 132) <= input(5);
output(5, 133) <= input(6);
output(5, 134) <= input(7);
output(5, 135) <= input(8);
output(5, 136) <= input(9);
output(5, 137) <= input(10);
output(5, 138) <= input(11);
output(5, 139) <= input(12);
output(5, 140) <= input(13);
output(5, 141) <= input(14);
output(5, 142) <= input(15);
output(5, 143) <= input(32);
output(5, 144) <= input(1);
output(5, 145) <= input(2);
output(5, 146) <= input(3);
output(5, 147) <= input(4);
output(5, 148) <= input(5);
output(5, 149) <= input(6);
output(5, 150) <= input(7);
output(5, 151) <= input(8);
output(5, 152) <= input(9);
output(5, 153) <= input(10);
output(5, 154) <= input(11);
output(5, 155) <= input(12);
output(5, 156) <= input(13);
output(5, 157) <= input(14);
output(5, 158) <= input(15);
output(5, 159) <= input(32);
output(5, 160) <= input(17);
output(5, 161) <= input(18);
output(5, 162) <= input(19);
output(5, 163) <= input(20);
output(5, 164) <= input(21);
output(5, 165) <= input(22);
output(5, 166) <= input(23);
output(5, 167) <= input(24);
output(5, 168) <= input(25);
output(5, 169) <= input(26);
output(5, 170) <= input(27);
output(5, 171) <= input(28);
output(5, 172) <= input(29);
output(5, 173) <= input(30);
output(5, 174) <= input(31);
output(5, 175) <= input(33);
output(5, 176) <= input(17);
output(5, 177) <= input(18);
output(5, 178) <= input(19);
output(5, 179) <= input(20);
output(5, 180) <= input(21);
output(5, 181) <= input(22);
output(5, 182) <= input(23);
output(5, 183) <= input(24);
output(5, 184) <= input(25);
output(5, 185) <= input(26);
output(5, 186) <= input(27);
output(5, 187) <= input(28);
output(5, 188) <= input(29);
output(5, 189) <= input(30);
output(5, 190) <= input(31);
output(5, 191) <= input(33);
output(5, 192) <= input(17);
output(5, 193) <= input(18);
output(5, 194) <= input(19);
output(5, 195) <= input(20);
output(5, 196) <= input(21);
output(5, 197) <= input(22);
output(5, 198) <= input(23);
output(5, 199) <= input(24);
output(5, 200) <= input(25);
output(5, 201) <= input(26);
output(5, 202) <= input(27);
output(5, 203) <= input(28);
output(5, 204) <= input(29);
output(5, 205) <= input(30);
output(5, 206) <= input(31);
output(5, 207) <= input(33);
output(5, 208) <= input(2);
output(5, 209) <= input(3);
output(5, 210) <= input(4);
output(5, 211) <= input(5);
output(5, 212) <= input(6);
output(5, 213) <= input(7);
output(5, 214) <= input(8);
output(5, 215) <= input(9);
output(5, 216) <= input(10);
output(5, 217) <= input(11);
output(5, 218) <= input(12);
output(5, 219) <= input(13);
output(5, 220) <= input(14);
output(5, 221) <= input(15);
output(5, 222) <= input(32);
output(5, 223) <= input(34);
output(5, 224) <= input(2);
output(5, 225) <= input(3);
output(5, 226) <= input(4);
output(5, 227) <= input(5);
output(5, 228) <= input(6);
output(5, 229) <= input(7);
output(5, 230) <= input(8);
output(5, 231) <= input(9);
output(5, 232) <= input(10);
output(5, 233) <= input(11);
output(5, 234) <= input(12);
output(5, 235) <= input(13);
output(5, 236) <= input(14);
output(5, 237) <= input(15);
output(5, 238) <= input(32);
output(5, 239) <= input(34);
output(5, 240) <= input(18);
output(5, 241) <= input(19);
output(5, 242) <= input(20);
output(5, 243) <= input(21);
output(5, 244) <= input(22);
output(5, 245) <= input(23);
output(5, 246) <= input(24);
output(5, 247) <= input(25);
output(5, 248) <= input(26);
output(5, 249) <= input(27);
output(5, 250) <= input(28);
output(5, 251) <= input(29);
output(5, 252) <= input(30);
output(5, 253) <= input(31);
output(5, 254) <= input(33);
output(5, 255) <= input(35);
when "0010" =>
output(0, 0) <= input(0);
output(0, 1) <= input(1);
output(0, 2) <= input(2);
output(0, 3) <= input(3);
output(0, 4) <= input(4);
output(0, 5) <= input(5);
output(0, 6) <= input(6);
output(0, 7) <= input(7);
output(0, 8) <= input(8);
output(0, 9) <= input(9);
output(0, 10) <= input(10);
output(0, 11) <= input(11);
output(0, 12) <= input(12);
output(0, 13) <= input(13);
output(0, 14) <= input(14);
output(0, 15) <= input(15);
output(0, 16) <= input(0);
output(0, 17) <= input(1);
output(0, 18) <= input(2);
output(0, 19) <= input(3);
output(0, 20) <= input(4);
output(0, 21) <= input(5);
output(0, 22) <= input(6);
output(0, 23) <= input(7);
output(0, 24) <= input(8);
output(0, 25) <= input(9);
output(0, 26) <= input(10);
output(0, 27) <= input(11);
output(0, 28) <= input(12);
output(0, 29) <= input(13);
output(0, 30) <= input(14);
output(0, 31) <= input(15);
output(0, 32) <= input(0);
output(0, 33) <= input(1);
output(0, 34) <= input(2);
output(0, 35) <= input(3);
output(0, 36) <= input(4);
output(0, 37) <= input(5);
output(0, 38) <= input(6);
output(0, 39) <= input(7);
output(0, 40) <= input(8);
output(0, 41) <= input(9);
output(0, 42) <= input(10);
output(0, 43) <= input(11);
output(0, 44) <= input(12);
output(0, 45) <= input(13);
output(0, 46) <= input(14);
output(0, 47) <= input(15);
output(0, 48) <= input(16);
output(0, 49) <= input(17);
output(0, 50) <= input(18);
output(0, 51) <= input(19);
output(0, 52) <= input(20);
output(0, 53) <= input(21);
output(0, 54) <= input(22);
output(0, 55) <= input(23);
output(0, 56) <= input(24);
output(0, 57) <= input(25);
output(0, 58) <= input(26);
output(0, 59) <= input(27);
output(0, 60) <= input(28);
output(0, 61) <= input(29);
output(0, 62) <= input(30);
output(0, 63) <= input(31);
output(0, 64) <= input(16);
output(0, 65) <= input(17);
output(0, 66) <= input(18);
output(0, 67) <= input(19);
output(0, 68) <= input(20);
output(0, 69) <= input(21);
output(0, 70) <= input(22);
output(0, 71) <= input(23);
output(0, 72) <= input(24);
output(0, 73) <= input(25);
output(0, 74) <= input(26);
output(0, 75) <= input(27);
output(0, 76) <= input(28);
output(0, 77) <= input(29);
output(0, 78) <= input(30);
output(0, 79) <= input(31);
output(0, 80) <= input(16);
output(0, 81) <= input(17);
output(0, 82) <= input(18);
output(0, 83) <= input(19);
output(0, 84) <= input(20);
output(0, 85) <= input(21);
output(0, 86) <= input(22);
output(0, 87) <= input(23);
output(0, 88) <= input(24);
output(0, 89) <= input(25);
output(0, 90) <= input(26);
output(0, 91) <= input(27);
output(0, 92) <= input(28);
output(0, 93) <= input(29);
output(0, 94) <= input(30);
output(0, 95) <= input(31);
output(0, 96) <= input(16);
output(0, 97) <= input(17);
output(0, 98) <= input(18);
output(0, 99) <= input(19);
output(0, 100) <= input(20);
output(0, 101) <= input(21);
output(0, 102) <= input(22);
output(0, 103) <= input(23);
output(0, 104) <= input(24);
output(0, 105) <= input(25);
output(0, 106) <= input(26);
output(0, 107) <= input(27);
output(0, 108) <= input(28);
output(0, 109) <= input(29);
output(0, 110) <= input(30);
output(0, 111) <= input(31);
output(0, 112) <= input(1);
output(0, 113) <= input(2);
output(0, 114) <= input(3);
output(0, 115) <= input(4);
output(0, 116) <= input(5);
output(0, 117) <= input(6);
output(0, 118) <= input(7);
output(0, 119) <= input(8);
output(0, 120) <= input(9);
output(0, 121) <= input(10);
output(0, 122) <= input(11);
output(0, 123) <= input(12);
output(0, 124) <= input(13);
output(0, 125) <= input(14);
output(0, 126) <= input(15);
output(0, 127) <= input(32);
output(0, 128) <= input(1);
output(0, 129) <= input(2);
output(0, 130) <= input(3);
output(0, 131) <= input(4);
output(0, 132) <= input(5);
output(0, 133) <= input(6);
output(0, 134) <= input(7);
output(0, 135) <= input(8);
output(0, 136) <= input(9);
output(0, 137) <= input(10);
output(0, 138) <= input(11);
output(0, 139) <= input(12);
output(0, 140) <= input(13);
output(0, 141) <= input(14);
output(0, 142) <= input(15);
output(0, 143) <= input(32);
output(0, 144) <= input(1);
output(0, 145) <= input(2);
output(0, 146) <= input(3);
output(0, 147) <= input(4);
output(0, 148) <= input(5);
output(0, 149) <= input(6);
output(0, 150) <= input(7);
output(0, 151) <= input(8);
output(0, 152) <= input(9);
output(0, 153) <= input(10);
output(0, 154) <= input(11);
output(0, 155) <= input(12);
output(0, 156) <= input(13);
output(0, 157) <= input(14);
output(0, 158) <= input(15);
output(0, 159) <= input(32);
output(0, 160) <= input(1);
output(0, 161) <= input(2);
output(0, 162) <= input(3);
output(0, 163) <= input(4);
output(0, 164) <= input(5);
output(0, 165) <= input(6);
output(0, 166) <= input(7);
output(0, 167) <= input(8);
output(0, 168) <= input(9);
output(0, 169) <= input(10);
output(0, 170) <= input(11);
output(0, 171) <= input(12);
output(0, 172) <= input(13);
output(0, 173) <= input(14);
output(0, 174) <= input(15);
output(0, 175) <= input(32);
output(0, 176) <= input(17);
output(0, 177) <= input(18);
output(0, 178) <= input(19);
output(0, 179) <= input(20);
output(0, 180) <= input(21);
output(0, 181) <= input(22);
output(0, 182) <= input(23);
output(0, 183) <= input(24);
output(0, 184) <= input(25);
output(0, 185) <= input(26);
output(0, 186) <= input(27);
output(0, 187) <= input(28);
output(0, 188) <= input(29);
output(0, 189) <= input(30);
output(0, 190) <= input(31);
output(0, 191) <= input(33);
output(0, 192) <= input(17);
output(0, 193) <= input(18);
output(0, 194) <= input(19);
output(0, 195) <= input(20);
output(0, 196) <= input(21);
output(0, 197) <= input(22);
output(0, 198) <= input(23);
output(0, 199) <= input(24);
output(0, 200) <= input(25);
output(0, 201) <= input(26);
output(0, 202) <= input(27);
output(0, 203) <= input(28);
output(0, 204) <= input(29);
output(0, 205) <= input(30);
output(0, 206) <= input(31);
output(0, 207) <= input(33);
output(0, 208) <= input(17);
output(0, 209) <= input(18);
output(0, 210) <= input(19);
output(0, 211) <= input(20);
output(0, 212) <= input(21);
output(0, 213) <= input(22);
output(0, 214) <= input(23);
output(0, 215) <= input(24);
output(0, 216) <= input(25);
output(0, 217) <= input(26);
output(0, 218) <= input(27);
output(0, 219) <= input(28);
output(0, 220) <= input(29);
output(0, 221) <= input(30);
output(0, 222) <= input(31);
output(0, 223) <= input(33);
output(0, 224) <= input(17);
output(0, 225) <= input(18);
output(0, 226) <= input(19);
output(0, 227) <= input(20);
output(0, 228) <= input(21);
output(0, 229) <= input(22);
output(0, 230) <= input(23);
output(0, 231) <= input(24);
output(0, 232) <= input(25);
output(0, 233) <= input(26);
output(0, 234) <= input(27);
output(0, 235) <= input(28);
output(0, 236) <= input(29);
output(0, 237) <= input(30);
output(0, 238) <= input(31);
output(0, 239) <= input(33);
output(0, 240) <= input(2);
output(0, 241) <= input(3);
output(0, 242) <= input(4);
output(0, 243) <= input(5);
output(0, 244) <= input(6);
output(0, 245) <= input(7);
output(0, 246) <= input(8);
output(0, 247) <= input(9);
output(0, 248) <= input(10);
output(0, 249) <= input(11);
output(0, 250) <= input(12);
output(0, 251) <= input(13);
output(0, 252) <= input(14);
output(0, 253) <= input(15);
output(0, 254) <= input(32);
output(0, 255) <= input(34);
output(1, 0) <= input(0);
output(1, 1) <= input(1);
output(1, 2) <= input(2);
output(1, 3) <= input(3);
output(1, 4) <= input(4);
output(1, 5) <= input(5);
output(1, 6) <= input(6);
output(1, 7) <= input(7);
output(1, 8) <= input(8);
output(1, 9) <= input(9);
output(1, 10) <= input(10);
output(1, 11) <= input(11);
output(1, 12) <= input(12);
output(1, 13) <= input(13);
output(1, 14) <= input(14);
output(1, 15) <= input(15);
output(1, 16) <= input(0);
output(1, 17) <= input(1);
output(1, 18) <= input(2);
output(1, 19) <= input(3);
output(1, 20) <= input(4);
output(1, 21) <= input(5);
output(1, 22) <= input(6);
output(1, 23) <= input(7);
output(1, 24) <= input(8);
output(1, 25) <= input(9);
output(1, 26) <= input(10);
output(1, 27) <= input(11);
output(1, 28) <= input(12);
output(1, 29) <= input(13);
output(1, 30) <= input(14);
output(1, 31) <= input(15);
output(1, 32) <= input(0);
output(1, 33) <= input(1);
output(1, 34) <= input(2);
output(1, 35) <= input(3);
output(1, 36) <= input(4);
output(1, 37) <= input(5);
output(1, 38) <= input(6);
output(1, 39) <= input(7);
output(1, 40) <= input(8);
output(1, 41) <= input(9);
output(1, 42) <= input(10);
output(1, 43) <= input(11);
output(1, 44) <= input(12);
output(1, 45) <= input(13);
output(1, 46) <= input(14);
output(1, 47) <= input(15);
output(1, 48) <= input(0);
output(1, 49) <= input(1);
output(1, 50) <= input(2);
output(1, 51) <= input(3);
output(1, 52) <= input(4);
output(1, 53) <= input(5);
output(1, 54) <= input(6);
output(1, 55) <= input(7);
output(1, 56) <= input(8);
output(1, 57) <= input(9);
output(1, 58) <= input(10);
output(1, 59) <= input(11);
output(1, 60) <= input(12);
output(1, 61) <= input(13);
output(1, 62) <= input(14);
output(1, 63) <= input(15);
output(1, 64) <= input(0);
output(1, 65) <= input(1);
output(1, 66) <= input(2);
output(1, 67) <= input(3);
output(1, 68) <= input(4);
output(1, 69) <= input(5);
output(1, 70) <= input(6);
output(1, 71) <= input(7);
output(1, 72) <= input(8);
output(1, 73) <= input(9);
output(1, 74) <= input(10);
output(1, 75) <= input(11);
output(1, 76) <= input(12);
output(1, 77) <= input(13);
output(1, 78) <= input(14);
output(1, 79) <= input(15);
output(1, 80) <= input(16);
output(1, 81) <= input(17);
output(1, 82) <= input(18);
output(1, 83) <= input(19);
output(1, 84) <= input(20);
output(1, 85) <= input(21);
output(1, 86) <= input(22);
output(1, 87) <= input(23);
output(1, 88) <= input(24);
output(1, 89) <= input(25);
output(1, 90) <= input(26);
output(1, 91) <= input(27);
output(1, 92) <= input(28);
output(1, 93) <= input(29);
output(1, 94) <= input(30);
output(1, 95) <= input(31);
output(1, 96) <= input(16);
output(1, 97) <= input(17);
output(1, 98) <= input(18);
output(1, 99) <= input(19);
output(1, 100) <= input(20);
output(1, 101) <= input(21);
output(1, 102) <= input(22);
output(1, 103) <= input(23);
output(1, 104) <= input(24);
output(1, 105) <= input(25);
output(1, 106) <= input(26);
output(1, 107) <= input(27);
output(1, 108) <= input(28);
output(1, 109) <= input(29);
output(1, 110) <= input(30);
output(1, 111) <= input(31);
output(1, 112) <= input(16);
output(1, 113) <= input(17);
output(1, 114) <= input(18);
output(1, 115) <= input(19);
output(1, 116) <= input(20);
output(1, 117) <= input(21);
output(1, 118) <= input(22);
output(1, 119) <= input(23);
output(1, 120) <= input(24);
output(1, 121) <= input(25);
output(1, 122) <= input(26);
output(1, 123) <= input(27);
output(1, 124) <= input(28);
output(1, 125) <= input(29);
output(1, 126) <= input(30);
output(1, 127) <= input(31);
output(1, 128) <= input(16);
output(1, 129) <= input(17);
output(1, 130) <= input(18);
output(1, 131) <= input(19);
output(1, 132) <= input(20);
output(1, 133) <= input(21);
output(1, 134) <= input(22);
output(1, 135) <= input(23);
output(1, 136) <= input(24);
output(1, 137) <= input(25);
output(1, 138) <= input(26);
output(1, 139) <= input(27);
output(1, 140) <= input(28);
output(1, 141) <= input(29);
output(1, 142) <= input(30);
output(1, 143) <= input(31);
output(1, 144) <= input(16);
output(1, 145) <= input(17);
output(1, 146) <= input(18);
output(1, 147) <= input(19);
output(1, 148) <= input(20);
output(1, 149) <= input(21);
output(1, 150) <= input(22);
output(1, 151) <= input(23);
output(1, 152) <= input(24);
output(1, 153) <= input(25);
output(1, 154) <= input(26);
output(1, 155) <= input(27);
output(1, 156) <= input(28);
output(1, 157) <= input(29);
output(1, 158) <= input(30);
output(1, 159) <= input(31);
output(1, 160) <= input(1);
output(1, 161) <= input(2);
output(1, 162) <= input(3);
output(1, 163) <= input(4);
output(1, 164) <= input(5);
output(1, 165) <= input(6);
output(1, 166) <= input(7);
output(1, 167) <= input(8);
output(1, 168) <= input(9);
output(1, 169) <= input(10);
output(1, 170) <= input(11);
output(1, 171) <= input(12);
output(1, 172) <= input(13);
output(1, 173) <= input(14);
output(1, 174) <= input(15);
output(1, 175) <= input(32);
output(1, 176) <= input(1);
output(1, 177) <= input(2);
output(1, 178) <= input(3);
output(1, 179) <= input(4);
output(1, 180) <= input(5);
output(1, 181) <= input(6);
output(1, 182) <= input(7);
output(1, 183) <= input(8);
output(1, 184) <= input(9);
output(1, 185) <= input(10);
output(1, 186) <= input(11);
output(1, 187) <= input(12);
output(1, 188) <= input(13);
output(1, 189) <= input(14);
output(1, 190) <= input(15);
output(1, 191) <= input(32);
output(1, 192) <= input(1);
output(1, 193) <= input(2);
output(1, 194) <= input(3);
output(1, 195) <= input(4);
output(1, 196) <= input(5);
output(1, 197) <= input(6);
output(1, 198) <= input(7);
output(1, 199) <= input(8);
output(1, 200) <= input(9);
output(1, 201) <= input(10);
output(1, 202) <= input(11);
output(1, 203) <= input(12);
output(1, 204) <= input(13);
output(1, 205) <= input(14);
output(1, 206) <= input(15);
output(1, 207) <= input(32);
output(1, 208) <= input(1);
output(1, 209) <= input(2);
output(1, 210) <= input(3);
output(1, 211) <= input(4);
output(1, 212) <= input(5);
output(1, 213) <= input(6);
output(1, 214) <= input(7);
output(1, 215) <= input(8);
output(1, 216) <= input(9);
output(1, 217) <= input(10);
output(1, 218) <= input(11);
output(1, 219) <= input(12);
output(1, 220) <= input(13);
output(1, 221) <= input(14);
output(1, 222) <= input(15);
output(1, 223) <= input(32);
output(1, 224) <= input(1);
output(1, 225) <= input(2);
output(1, 226) <= input(3);
output(1, 227) <= input(4);
output(1, 228) <= input(5);
output(1, 229) <= input(6);
output(1, 230) <= input(7);
output(1, 231) <= input(8);
output(1, 232) <= input(9);
output(1, 233) <= input(10);
output(1, 234) <= input(11);
output(1, 235) <= input(12);
output(1, 236) <= input(13);
output(1, 237) <= input(14);
output(1, 238) <= input(15);
output(1, 239) <= input(32);
output(1, 240) <= input(17);
output(1, 241) <= input(18);
output(1, 242) <= input(19);
output(1, 243) <= input(20);
output(1, 244) <= input(21);
output(1, 245) <= input(22);
output(1, 246) <= input(23);
output(1, 247) <= input(24);
output(1, 248) <= input(25);
output(1, 249) <= input(26);
output(1, 250) <= input(27);
output(1, 251) <= input(28);
output(1, 252) <= input(29);
output(1, 253) <= input(30);
output(1, 254) <= input(31);
output(1, 255) <= input(33);
output(2, 0) <= input(0);
output(2, 1) <= input(1);
output(2, 2) <= input(2);
output(2, 3) <= input(3);
output(2, 4) <= input(4);
output(2, 5) <= input(5);
output(2, 6) <= input(6);
output(2, 7) <= input(7);
output(2, 8) <= input(8);
output(2, 9) <= input(9);
output(2, 10) <= input(10);
output(2, 11) <= input(11);
output(2, 12) <= input(12);
output(2, 13) <= input(13);
output(2, 14) <= input(14);
output(2, 15) <= input(15);
output(2, 16) <= input(0);
output(2, 17) <= input(1);
output(2, 18) <= input(2);
output(2, 19) <= input(3);
output(2, 20) <= input(4);
output(2, 21) <= input(5);
output(2, 22) <= input(6);
output(2, 23) <= input(7);
output(2, 24) <= input(8);
output(2, 25) <= input(9);
output(2, 26) <= input(10);
output(2, 27) <= input(11);
output(2, 28) <= input(12);
output(2, 29) <= input(13);
output(2, 30) <= input(14);
output(2, 31) <= input(15);
output(2, 32) <= input(0);
output(2, 33) <= input(1);
output(2, 34) <= input(2);
output(2, 35) <= input(3);
output(2, 36) <= input(4);
output(2, 37) <= input(5);
output(2, 38) <= input(6);
output(2, 39) <= input(7);
output(2, 40) <= input(8);
output(2, 41) <= input(9);
output(2, 42) <= input(10);
output(2, 43) <= input(11);
output(2, 44) <= input(12);
output(2, 45) <= input(13);
output(2, 46) <= input(14);
output(2, 47) <= input(15);
output(2, 48) <= input(0);
output(2, 49) <= input(1);
output(2, 50) <= input(2);
output(2, 51) <= input(3);
output(2, 52) <= input(4);
output(2, 53) <= input(5);
output(2, 54) <= input(6);
output(2, 55) <= input(7);
output(2, 56) <= input(8);
output(2, 57) <= input(9);
output(2, 58) <= input(10);
output(2, 59) <= input(11);
output(2, 60) <= input(12);
output(2, 61) <= input(13);
output(2, 62) <= input(14);
output(2, 63) <= input(15);
output(2, 64) <= input(0);
output(2, 65) <= input(1);
output(2, 66) <= input(2);
output(2, 67) <= input(3);
output(2, 68) <= input(4);
output(2, 69) <= input(5);
output(2, 70) <= input(6);
output(2, 71) <= input(7);
output(2, 72) <= input(8);
output(2, 73) <= input(9);
output(2, 74) <= input(10);
output(2, 75) <= input(11);
output(2, 76) <= input(12);
output(2, 77) <= input(13);
output(2, 78) <= input(14);
output(2, 79) <= input(15);
output(2, 80) <= input(0);
output(2, 81) <= input(1);
output(2, 82) <= input(2);
output(2, 83) <= input(3);
output(2, 84) <= input(4);
output(2, 85) <= input(5);
output(2, 86) <= input(6);
output(2, 87) <= input(7);
output(2, 88) <= input(8);
output(2, 89) <= input(9);
output(2, 90) <= input(10);
output(2, 91) <= input(11);
output(2, 92) <= input(12);
output(2, 93) <= input(13);
output(2, 94) <= input(14);
output(2, 95) <= input(15);
output(2, 96) <= input(0);
output(2, 97) <= input(1);
output(2, 98) <= input(2);
output(2, 99) <= input(3);
output(2, 100) <= input(4);
output(2, 101) <= input(5);
output(2, 102) <= input(6);
output(2, 103) <= input(7);
output(2, 104) <= input(8);
output(2, 105) <= input(9);
output(2, 106) <= input(10);
output(2, 107) <= input(11);
output(2, 108) <= input(12);
output(2, 109) <= input(13);
output(2, 110) <= input(14);
output(2, 111) <= input(15);
output(2, 112) <= input(16);
output(2, 113) <= input(17);
output(2, 114) <= input(18);
output(2, 115) <= input(19);
output(2, 116) <= input(20);
output(2, 117) <= input(21);
output(2, 118) <= input(22);
output(2, 119) <= input(23);
output(2, 120) <= input(24);
output(2, 121) <= input(25);
output(2, 122) <= input(26);
output(2, 123) <= input(27);
output(2, 124) <= input(28);
output(2, 125) <= input(29);
output(2, 126) <= input(30);
output(2, 127) <= input(31);
output(2, 128) <= input(16);
output(2, 129) <= input(17);
output(2, 130) <= input(18);
output(2, 131) <= input(19);
output(2, 132) <= input(20);
output(2, 133) <= input(21);
output(2, 134) <= input(22);
output(2, 135) <= input(23);
output(2, 136) <= input(24);
output(2, 137) <= input(25);
output(2, 138) <= input(26);
output(2, 139) <= input(27);
output(2, 140) <= input(28);
output(2, 141) <= input(29);
output(2, 142) <= input(30);
output(2, 143) <= input(31);
output(2, 144) <= input(16);
output(2, 145) <= input(17);
output(2, 146) <= input(18);
output(2, 147) <= input(19);
output(2, 148) <= input(20);
output(2, 149) <= input(21);
output(2, 150) <= input(22);
output(2, 151) <= input(23);
output(2, 152) <= input(24);
output(2, 153) <= input(25);
output(2, 154) <= input(26);
output(2, 155) <= input(27);
output(2, 156) <= input(28);
output(2, 157) <= input(29);
output(2, 158) <= input(30);
output(2, 159) <= input(31);
output(2, 160) <= input(16);
output(2, 161) <= input(17);
output(2, 162) <= input(18);
output(2, 163) <= input(19);
output(2, 164) <= input(20);
output(2, 165) <= input(21);
output(2, 166) <= input(22);
output(2, 167) <= input(23);
output(2, 168) <= input(24);
output(2, 169) <= input(25);
output(2, 170) <= input(26);
output(2, 171) <= input(27);
output(2, 172) <= input(28);
output(2, 173) <= input(29);
output(2, 174) <= input(30);
output(2, 175) <= input(31);
output(2, 176) <= input(16);
output(2, 177) <= input(17);
output(2, 178) <= input(18);
output(2, 179) <= input(19);
output(2, 180) <= input(20);
output(2, 181) <= input(21);
output(2, 182) <= input(22);
output(2, 183) <= input(23);
output(2, 184) <= input(24);
output(2, 185) <= input(25);
output(2, 186) <= input(26);
output(2, 187) <= input(27);
output(2, 188) <= input(28);
output(2, 189) <= input(29);
output(2, 190) <= input(30);
output(2, 191) <= input(31);
output(2, 192) <= input(16);
output(2, 193) <= input(17);
output(2, 194) <= input(18);
output(2, 195) <= input(19);
output(2, 196) <= input(20);
output(2, 197) <= input(21);
output(2, 198) <= input(22);
output(2, 199) <= input(23);
output(2, 200) <= input(24);
output(2, 201) <= input(25);
output(2, 202) <= input(26);
output(2, 203) <= input(27);
output(2, 204) <= input(28);
output(2, 205) <= input(29);
output(2, 206) <= input(30);
output(2, 207) <= input(31);
output(2, 208) <= input(16);
output(2, 209) <= input(17);
output(2, 210) <= input(18);
output(2, 211) <= input(19);
output(2, 212) <= input(20);
output(2, 213) <= input(21);
output(2, 214) <= input(22);
output(2, 215) <= input(23);
output(2, 216) <= input(24);
output(2, 217) <= input(25);
output(2, 218) <= input(26);
output(2, 219) <= input(27);
output(2, 220) <= input(28);
output(2, 221) <= input(29);
output(2, 222) <= input(30);
output(2, 223) <= input(31);
output(2, 224) <= input(16);
output(2, 225) <= input(17);
output(2, 226) <= input(18);
output(2, 227) <= input(19);
output(2, 228) <= input(20);
output(2, 229) <= input(21);
output(2, 230) <= input(22);
output(2, 231) <= input(23);
output(2, 232) <= input(24);
output(2, 233) <= input(25);
output(2, 234) <= input(26);
output(2, 235) <= input(27);
output(2, 236) <= input(28);
output(2, 237) <= input(29);
output(2, 238) <= input(30);
output(2, 239) <= input(31);
output(2, 240) <= input(1);
output(2, 241) <= input(2);
output(2, 242) <= input(3);
output(2, 243) <= input(4);
output(2, 244) <= input(5);
output(2, 245) <= input(6);
output(2, 246) <= input(7);
output(2, 247) <= input(8);
output(2, 248) <= input(9);
output(2, 249) <= input(10);
output(2, 250) <= input(11);
output(2, 251) <= input(12);
output(2, 252) <= input(13);
output(2, 253) <= input(14);
output(2, 254) <= input(15);
output(2, 255) <= input(32);
output(3, 0) <= input(0);
output(3, 1) <= input(1);
output(3, 2) <= input(2);
output(3, 3) <= input(3);
output(3, 4) <= input(4);
output(3, 5) <= input(5);
output(3, 6) <= input(6);
output(3, 7) <= input(7);
output(3, 8) <= input(8);
output(3, 9) <= input(9);
output(3, 10) <= input(10);
output(3, 11) <= input(11);
output(3, 12) <= input(12);
output(3, 13) <= input(13);
output(3, 14) <= input(14);
output(3, 15) <= input(15);
output(3, 16) <= input(0);
output(3, 17) <= input(1);
output(3, 18) <= input(2);
output(3, 19) <= input(3);
output(3, 20) <= input(4);
output(3, 21) <= input(5);
output(3, 22) <= input(6);
output(3, 23) <= input(7);
output(3, 24) <= input(8);
output(3, 25) <= input(9);
output(3, 26) <= input(10);
output(3, 27) <= input(11);
output(3, 28) <= input(12);
output(3, 29) <= input(13);
output(3, 30) <= input(14);
output(3, 31) <= input(15);
output(3, 32) <= input(0);
output(3, 33) <= input(1);
output(3, 34) <= input(2);
output(3, 35) <= input(3);
output(3, 36) <= input(4);
output(3, 37) <= input(5);
output(3, 38) <= input(6);
output(3, 39) <= input(7);
output(3, 40) <= input(8);
output(3, 41) <= input(9);
output(3, 42) <= input(10);
output(3, 43) <= input(11);
output(3, 44) <= input(12);
output(3, 45) <= input(13);
output(3, 46) <= input(14);
output(3, 47) <= input(15);
output(3, 48) <= input(0);
output(3, 49) <= input(1);
output(3, 50) <= input(2);
output(3, 51) <= input(3);
output(3, 52) <= input(4);
output(3, 53) <= input(5);
output(3, 54) <= input(6);
output(3, 55) <= input(7);
output(3, 56) <= input(8);
output(3, 57) <= input(9);
output(3, 58) <= input(10);
output(3, 59) <= input(11);
output(3, 60) <= input(12);
output(3, 61) <= input(13);
output(3, 62) <= input(14);
output(3, 63) <= input(15);
output(3, 64) <= input(0);
output(3, 65) <= input(1);
output(3, 66) <= input(2);
output(3, 67) <= input(3);
output(3, 68) <= input(4);
output(3, 69) <= input(5);
output(3, 70) <= input(6);
output(3, 71) <= input(7);
output(3, 72) <= input(8);
output(3, 73) <= input(9);
output(3, 74) <= input(10);
output(3, 75) <= input(11);
output(3, 76) <= input(12);
output(3, 77) <= input(13);
output(3, 78) <= input(14);
output(3, 79) <= input(15);
output(3, 80) <= input(0);
output(3, 81) <= input(1);
output(3, 82) <= input(2);
output(3, 83) <= input(3);
output(3, 84) <= input(4);
output(3, 85) <= input(5);
output(3, 86) <= input(6);
output(3, 87) <= input(7);
output(3, 88) <= input(8);
output(3, 89) <= input(9);
output(3, 90) <= input(10);
output(3, 91) <= input(11);
output(3, 92) <= input(12);
output(3, 93) <= input(13);
output(3, 94) <= input(14);
output(3, 95) <= input(15);
output(3, 96) <= input(0);
output(3, 97) <= input(1);
output(3, 98) <= input(2);
output(3, 99) <= input(3);
output(3, 100) <= input(4);
output(3, 101) <= input(5);
output(3, 102) <= input(6);
output(3, 103) <= input(7);
output(3, 104) <= input(8);
output(3, 105) <= input(9);
output(3, 106) <= input(10);
output(3, 107) <= input(11);
output(3, 108) <= input(12);
output(3, 109) <= input(13);
output(3, 110) <= input(14);
output(3, 111) <= input(15);
output(3, 112) <= input(0);
output(3, 113) <= input(1);
output(3, 114) <= input(2);
output(3, 115) <= input(3);
output(3, 116) <= input(4);
output(3, 117) <= input(5);
output(3, 118) <= input(6);
output(3, 119) <= input(7);
output(3, 120) <= input(8);
output(3, 121) <= input(9);
output(3, 122) <= input(10);
output(3, 123) <= input(11);
output(3, 124) <= input(12);
output(3, 125) <= input(13);
output(3, 126) <= input(14);
output(3, 127) <= input(15);
output(3, 128) <= input(0);
output(3, 129) <= input(1);
output(3, 130) <= input(2);
output(3, 131) <= input(3);
output(3, 132) <= input(4);
output(3, 133) <= input(5);
output(3, 134) <= input(6);
output(3, 135) <= input(7);
output(3, 136) <= input(8);
output(3, 137) <= input(9);
output(3, 138) <= input(10);
output(3, 139) <= input(11);
output(3, 140) <= input(12);
output(3, 141) <= input(13);
output(3, 142) <= input(14);
output(3, 143) <= input(15);
output(3, 144) <= input(0);
output(3, 145) <= input(1);
output(3, 146) <= input(2);
output(3, 147) <= input(3);
output(3, 148) <= input(4);
output(3, 149) <= input(5);
output(3, 150) <= input(6);
output(3, 151) <= input(7);
output(3, 152) <= input(8);
output(3, 153) <= input(9);
output(3, 154) <= input(10);
output(3, 155) <= input(11);
output(3, 156) <= input(12);
output(3, 157) <= input(13);
output(3, 158) <= input(14);
output(3, 159) <= input(15);
output(3, 160) <= input(0);
output(3, 161) <= input(1);
output(3, 162) <= input(2);
output(3, 163) <= input(3);
output(3, 164) <= input(4);
output(3, 165) <= input(5);
output(3, 166) <= input(6);
output(3, 167) <= input(7);
output(3, 168) <= input(8);
output(3, 169) <= input(9);
output(3, 170) <= input(10);
output(3, 171) <= input(11);
output(3, 172) <= input(12);
output(3, 173) <= input(13);
output(3, 174) <= input(14);
output(3, 175) <= input(15);
output(3, 176) <= input(0);
output(3, 177) <= input(1);
output(3, 178) <= input(2);
output(3, 179) <= input(3);
output(3, 180) <= input(4);
output(3, 181) <= input(5);
output(3, 182) <= input(6);
output(3, 183) <= input(7);
output(3, 184) <= input(8);
output(3, 185) <= input(9);
output(3, 186) <= input(10);
output(3, 187) <= input(11);
output(3, 188) <= input(12);
output(3, 189) <= input(13);
output(3, 190) <= input(14);
output(3, 191) <= input(15);
output(3, 192) <= input(0);
output(3, 193) <= input(1);
output(3, 194) <= input(2);
output(3, 195) <= input(3);
output(3, 196) <= input(4);
output(3, 197) <= input(5);
output(3, 198) <= input(6);
output(3, 199) <= input(7);
output(3, 200) <= input(8);
output(3, 201) <= input(9);
output(3, 202) <= input(10);
output(3, 203) <= input(11);
output(3, 204) <= input(12);
output(3, 205) <= input(13);
output(3, 206) <= input(14);
output(3, 207) <= input(15);
output(3, 208) <= input(0);
output(3, 209) <= input(1);
output(3, 210) <= input(2);
output(3, 211) <= input(3);
output(3, 212) <= input(4);
output(3, 213) <= input(5);
output(3, 214) <= input(6);
output(3, 215) <= input(7);
output(3, 216) <= input(8);
output(3, 217) <= input(9);
output(3, 218) <= input(10);
output(3, 219) <= input(11);
output(3, 220) <= input(12);
output(3, 221) <= input(13);
output(3, 222) <= input(14);
output(3, 223) <= input(15);
output(3, 224) <= input(0);
output(3, 225) <= input(1);
output(3, 226) <= input(2);
output(3, 227) <= input(3);
output(3, 228) <= input(4);
output(3, 229) <= input(5);
output(3, 230) <= input(6);
output(3, 231) <= input(7);
output(3, 232) <= input(8);
output(3, 233) <= input(9);
output(3, 234) <= input(10);
output(3, 235) <= input(11);
output(3, 236) <= input(12);
output(3, 237) <= input(13);
output(3, 238) <= input(14);
output(3, 239) <= input(15);
output(3, 240) <= input(16);
output(3, 241) <= input(17);
output(3, 242) <= input(18);
output(3, 243) <= input(19);
output(3, 244) <= input(20);
output(3, 245) <= input(21);
output(3, 246) <= input(22);
output(3, 247) <= input(23);
output(3, 248) <= input(24);
output(3, 249) <= input(25);
output(3, 250) <= input(26);
output(3, 251) <= input(27);
output(3, 252) <= input(28);
output(3, 253) <= input(29);
output(3, 254) <= input(30);
output(3, 255) <= input(31);
output(4, 0) <= input(0);
output(4, 1) <= input(1);
output(4, 2) <= input(2);
output(4, 3) <= input(3);
output(4, 4) <= input(4);
output(4, 5) <= input(5);
output(4, 6) <= input(6);
output(4, 7) <= input(7);
output(4, 8) <= input(8);
output(4, 9) <= input(9);
output(4, 10) <= input(10);
output(4, 11) <= input(11);
output(4, 12) <= input(12);
output(4, 13) <= input(13);
output(4, 14) <= input(14);
output(4, 15) <= input(15);
output(4, 16) <= input(0);
output(4, 17) <= input(1);
output(4, 18) <= input(2);
output(4, 19) <= input(3);
output(4, 20) <= input(4);
output(4, 21) <= input(5);
output(4, 22) <= input(6);
output(4, 23) <= input(7);
output(4, 24) <= input(8);
output(4, 25) <= input(9);
output(4, 26) <= input(10);
output(4, 27) <= input(11);
output(4, 28) <= input(12);
output(4, 29) <= input(13);
output(4, 30) <= input(14);
output(4, 31) <= input(15);
output(4, 32) <= input(0);
output(4, 33) <= input(1);
output(4, 34) <= input(2);
output(4, 35) <= input(3);
output(4, 36) <= input(4);
output(4, 37) <= input(5);
output(4, 38) <= input(6);
output(4, 39) <= input(7);
output(4, 40) <= input(8);
output(4, 41) <= input(9);
output(4, 42) <= input(10);
output(4, 43) <= input(11);
output(4, 44) <= input(12);
output(4, 45) <= input(13);
output(4, 46) <= input(14);
output(4, 47) <= input(15);
output(4, 48) <= input(0);
output(4, 49) <= input(1);
output(4, 50) <= input(2);
output(4, 51) <= input(3);
output(4, 52) <= input(4);
output(4, 53) <= input(5);
output(4, 54) <= input(6);
output(4, 55) <= input(7);
output(4, 56) <= input(8);
output(4, 57) <= input(9);
output(4, 58) <= input(10);
output(4, 59) <= input(11);
output(4, 60) <= input(12);
output(4, 61) <= input(13);
output(4, 62) <= input(14);
output(4, 63) <= input(15);
output(4, 64) <= input(0);
output(4, 65) <= input(1);
output(4, 66) <= input(2);
output(4, 67) <= input(3);
output(4, 68) <= input(4);
output(4, 69) <= input(5);
output(4, 70) <= input(6);
output(4, 71) <= input(7);
output(4, 72) <= input(8);
output(4, 73) <= input(9);
output(4, 74) <= input(10);
output(4, 75) <= input(11);
output(4, 76) <= input(12);
output(4, 77) <= input(13);
output(4, 78) <= input(14);
output(4, 79) <= input(15);
output(4, 80) <= input(0);
output(4, 81) <= input(1);
output(4, 82) <= input(2);
output(4, 83) <= input(3);
output(4, 84) <= input(4);
output(4, 85) <= input(5);
output(4, 86) <= input(6);
output(4, 87) <= input(7);
output(4, 88) <= input(8);
output(4, 89) <= input(9);
output(4, 90) <= input(10);
output(4, 91) <= input(11);
output(4, 92) <= input(12);
output(4, 93) <= input(13);
output(4, 94) <= input(14);
output(4, 95) <= input(15);
output(4, 96) <= input(0);
output(4, 97) <= input(1);
output(4, 98) <= input(2);
output(4, 99) <= input(3);
output(4, 100) <= input(4);
output(4, 101) <= input(5);
output(4, 102) <= input(6);
output(4, 103) <= input(7);
output(4, 104) <= input(8);
output(4, 105) <= input(9);
output(4, 106) <= input(10);
output(4, 107) <= input(11);
output(4, 108) <= input(12);
output(4, 109) <= input(13);
output(4, 110) <= input(14);
output(4, 111) <= input(15);
output(4, 112) <= input(0);
output(4, 113) <= input(1);
output(4, 114) <= input(2);
output(4, 115) <= input(3);
output(4, 116) <= input(4);
output(4, 117) <= input(5);
output(4, 118) <= input(6);
output(4, 119) <= input(7);
output(4, 120) <= input(8);
output(4, 121) <= input(9);
output(4, 122) <= input(10);
output(4, 123) <= input(11);
output(4, 124) <= input(12);
output(4, 125) <= input(13);
output(4, 126) <= input(14);
output(4, 127) <= input(15);
output(4, 128) <= input(0);
output(4, 129) <= input(1);
output(4, 130) <= input(2);
output(4, 131) <= input(3);
output(4, 132) <= input(4);
output(4, 133) <= input(5);
output(4, 134) <= input(6);
output(4, 135) <= input(7);
output(4, 136) <= input(8);
output(4, 137) <= input(9);
output(4, 138) <= input(10);
output(4, 139) <= input(11);
output(4, 140) <= input(12);
output(4, 141) <= input(13);
output(4, 142) <= input(14);
output(4, 143) <= input(15);
output(4, 144) <= input(0);
output(4, 145) <= input(1);
output(4, 146) <= input(2);
output(4, 147) <= input(3);
output(4, 148) <= input(4);
output(4, 149) <= input(5);
output(4, 150) <= input(6);
output(4, 151) <= input(7);
output(4, 152) <= input(8);
output(4, 153) <= input(9);
output(4, 154) <= input(10);
output(4, 155) <= input(11);
output(4, 156) <= input(12);
output(4, 157) <= input(13);
output(4, 158) <= input(14);
output(4, 159) <= input(15);
output(4, 160) <= input(0);
output(4, 161) <= input(1);
output(4, 162) <= input(2);
output(4, 163) <= input(3);
output(4, 164) <= input(4);
output(4, 165) <= input(5);
output(4, 166) <= input(6);
output(4, 167) <= input(7);
output(4, 168) <= input(8);
output(4, 169) <= input(9);
output(4, 170) <= input(10);
output(4, 171) <= input(11);
output(4, 172) <= input(12);
output(4, 173) <= input(13);
output(4, 174) <= input(14);
output(4, 175) <= input(15);
output(4, 176) <= input(0);
output(4, 177) <= input(1);
output(4, 178) <= input(2);
output(4, 179) <= input(3);
output(4, 180) <= input(4);
output(4, 181) <= input(5);
output(4, 182) <= input(6);
output(4, 183) <= input(7);
output(4, 184) <= input(8);
output(4, 185) <= input(9);
output(4, 186) <= input(10);
output(4, 187) <= input(11);
output(4, 188) <= input(12);
output(4, 189) <= input(13);
output(4, 190) <= input(14);
output(4, 191) <= input(15);
output(4, 192) <= input(0);
output(4, 193) <= input(1);
output(4, 194) <= input(2);
output(4, 195) <= input(3);
output(4, 196) <= input(4);
output(4, 197) <= input(5);
output(4, 198) <= input(6);
output(4, 199) <= input(7);
output(4, 200) <= input(8);
output(4, 201) <= input(9);
output(4, 202) <= input(10);
output(4, 203) <= input(11);
output(4, 204) <= input(12);
output(4, 205) <= input(13);
output(4, 206) <= input(14);
output(4, 207) <= input(15);
output(4, 208) <= input(0);
output(4, 209) <= input(1);
output(4, 210) <= input(2);
output(4, 211) <= input(3);
output(4, 212) <= input(4);
output(4, 213) <= input(5);
output(4, 214) <= input(6);
output(4, 215) <= input(7);
output(4, 216) <= input(8);
output(4, 217) <= input(9);
output(4, 218) <= input(10);
output(4, 219) <= input(11);
output(4, 220) <= input(12);
output(4, 221) <= input(13);
output(4, 222) <= input(14);
output(4, 223) <= input(15);
output(4, 224) <= input(0);
output(4, 225) <= input(1);
output(4, 226) <= input(2);
output(4, 227) <= input(3);
output(4, 228) <= input(4);
output(4, 229) <= input(5);
output(4, 230) <= input(6);
output(4, 231) <= input(7);
output(4, 232) <= input(8);
output(4, 233) <= input(9);
output(4, 234) <= input(10);
output(4, 235) <= input(11);
output(4, 236) <= input(12);
output(4, 237) <= input(13);
output(4, 238) <= input(14);
output(4, 239) <= input(15);
output(4, 240) <= input(0);
output(4, 241) <= input(1);
output(4, 242) <= input(2);
output(4, 243) <= input(3);
output(4, 244) <= input(4);
output(4, 245) <= input(5);
output(4, 246) <= input(6);
output(4, 247) <= input(7);
output(4, 248) <= input(8);
output(4, 249) <= input(9);
output(4, 250) <= input(10);
output(4, 251) <= input(11);
output(4, 252) <= input(12);
output(4, 253) <= input(13);
output(4, 254) <= input(14);
output(4, 255) <= input(15);
output(5, 0) <= input(35);
output(5, 1) <= input(16);
output(5, 2) <= input(17);
output(5, 3) <= input(18);
output(5, 4) <= input(19);
output(5, 5) <= input(20);
output(5, 6) <= input(21);
output(5, 7) <= input(22);
output(5, 8) <= input(23);
output(5, 9) <= input(24);
output(5, 10) <= input(25);
output(5, 11) <= input(26);
output(5, 12) <= input(27);
output(5, 13) <= input(28);
output(5, 14) <= input(29);
output(5, 15) <= input(30);
output(5, 16) <= input(35);
output(5, 17) <= input(16);
output(5, 18) <= input(17);
output(5, 19) <= input(18);
output(5, 20) <= input(19);
output(5, 21) <= input(20);
output(5, 22) <= input(21);
output(5, 23) <= input(22);
output(5, 24) <= input(23);
output(5, 25) <= input(24);
output(5, 26) <= input(25);
output(5, 27) <= input(26);
output(5, 28) <= input(27);
output(5, 29) <= input(28);
output(5, 30) <= input(29);
output(5, 31) <= input(30);
output(5, 32) <= input(35);
output(5, 33) <= input(16);
output(5, 34) <= input(17);
output(5, 35) <= input(18);
output(5, 36) <= input(19);
output(5, 37) <= input(20);
output(5, 38) <= input(21);
output(5, 39) <= input(22);
output(5, 40) <= input(23);
output(5, 41) <= input(24);
output(5, 42) <= input(25);
output(5, 43) <= input(26);
output(5, 44) <= input(27);
output(5, 45) <= input(28);
output(5, 46) <= input(29);
output(5, 47) <= input(30);
output(5, 48) <= input(35);
output(5, 49) <= input(16);
output(5, 50) <= input(17);
output(5, 51) <= input(18);
output(5, 52) <= input(19);
output(5, 53) <= input(20);
output(5, 54) <= input(21);
output(5, 55) <= input(22);
output(5, 56) <= input(23);
output(5, 57) <= input(24);
output(5, 58) <= input(25);
output(5, 59) <= input(26);
output(5, 60) <= input(27);
output(5, 61) <= input(28);
output(5, 62) <= input(29);
output(5, 63) <= input(30);
output(5, 64) <= input(35);
output(5, 65) <= input(16);
output(5, 66) <= input(17);
output(5, 67) <= input(18);
output(5, 68) <= input(19);
output(5, 69) <= input(20);
output(5, 70) <= input(21);
output(5, 71) <= input(22);
output(5, 72) <= input(23);
output(5, 73) <= input(24);
output(5, 74) <= input(25);
output(5, 75) <= input(26);
output(5, 76) <= input(27);
output(5, 77) <= input(28);
output(5, 78) <= input(29);
output(5, 79) <= input(30);
output(5, 80) <= input(35);
output(5, 81) <= input(16);
output(5, 82) <= input(17);
output(5, 83) <= input(18);
output(5, 84) <= input(19);
output(5, 85) <= input(20);
output(5, 86) <= input(21);
output(5, 87) <= input(22);
output(5, 88) <= input(23);
output(5, 89) <= input(24);
output(5, 90) <= input(25);
output(5, 91) <= input(26);
output(5, 92) <= input(27);
output(5, 93) <= input(28);
output(5, 94) <= input(29);
output(5, 95) <= input(30);
output(5, 96) <= input(35);
output(5, 97) <= input(16);
output(5, 98) <= input(17);
output(5, 99) <= input(18);
output(5, 100) <= input(19);
output(5, 101) <= input(20);
output(5, 102) <= input(21);
output(5, 103) <= input(22);
output(5, 104) <= input(23);
output(5, 105) <= input(24);
output(5, 106) <= input(25);
output(5, 107) <= input(26);
output(5, 108) <= input(27);
output(5, 109) <= input(28);
output(5, 110) <= input(29);
output(5, 111) <= input(30);
output(5, 112) <= input(35);
output(5, 113) <= input(16);
output(5, 114) <= input(17);
output(5, 115) <= input(18);
output(5, 116) <= input(19);
output(5, 117) <= input(20);
output(5, 118) <= input(21);
output(5, 119) <= input(22);
output(5, 120) <= input(23);
output(5, 121) <= input(24);
output(5, 122) <= input(25);
output(5, 123) <= input(26);
output(5, 124) <= input(27);
output(5, 125) <= input(28);
output(5, 126) <= input(29);
output(5, 127) <= input(30);
output(5, 128) <= input(35);
output(5, 129) <= input(16);
output(5, 130) <= input(17);
output(5, 131) <= input(18);
output(5, 132) <= input(19);
output(5, 133) <= input(20);
output(5, 134) <= input(21);
output(5, 135) <= input(22);
output(5, 136) <= input(23);
output(5, 137) <= input(24);
output(5, 138) <= input(25);
output(5, 139) <= input(26);
output(5, 140) <= input(27);
output(5, 141) <= input(28);
output(5, 142) <= input(29);
output(5, 143) <= input(30);
output(5, 144) <= input(35);
output(5, 145) <= input(16);
output(5, 146) <= input(17);
output(5, 147) <= input(18);
output(5, 148) <= input(19);
output(5, 149) <= input(20);
output(5, 150) <= input(21);
output(5, 151) <= input(22);
output(5, 152) <= input(23);
output(5, 153) <= input(24);
output(5, 154) <= input(25);
output(5, 155) <= input(26);
output(5, 156) <= input(27);
output(5, 157) <= input(28);
output(5, 158) <= input(29);
output(5, 159) <= input(30);
output(5, 160) <= input(35);
output(5, 161) <= input(16);
output(5, 162) <= input(17);
output(5, 163) <= input(18);
output(5, 164) <= input(19);
output(5, 165) <= input(20);
output(5, 166) <= input(21);
output(5, 167) <= input(22);
output(5, 168) <= input(23);
output(5, 169) <= input(24);
output(5, 170) <= input(25);
output(5, 171) <= input(26);
output(5, 172) <= input(27);
output(5, 173) <= input(28);
output(5, 174) <= input(29);
output(5, 175) <= input(30);
output(5, 176) <= input(35);
output(5, 177) <= input(16);
output(5, 178) <= input(17);
output(5, 179) <= input(18);
output(5, 180) <= input(19);
output(5, 181) <= input(20);
output(5, 182) <= input(21);
output(5, 183) <= input(22);
output(5, 184) <= input(23);
output(5, 185) <= input(24);
output(5, 186) <= input(25);
output(5, 187) <= input(26);
output(5, 188) <= input(27);
output(5, 189) <= input(28);
output(5, 190) <= input(29);
output(5, 191) <= input(30);
output(5, 192) <= input(35);
output(5, 193) <= input(16);
output(5, 194) <= input(17);
output(5, 195) <= input(18);
output(5, 196) <= input(19);
output(5, 197) <= input(20);
output(5, 198) <= input(21);
output(5, 199) <= input(22);
output(5, 200) <= input(23);
output(5, 201) <= input(24);
output(5, 202) <= input(25);
output(5, 203) <= input(26);
output(5, 204) <= input(27);
output(5, 205) <= input(28);
output(5, 206) <= input(29);
output(5, 207) <= input(30);
output(5, 208) <= input(35);
output(5, 209) <= input(16);
output(5, 210) <= input(17);
output(5, 211) <= input(18);
output(5, 212) <= input(19);
output(5, 213) <= input(20);
output(5, 214) <= input(21);
output(5, 215) <= input(22);
output(5, 216) <= input(23);
output(5, 217) <= input(24);
output(5, 218) <= input(25);
output(5, 219) <= input(26);
output(5, 220) <= input(27);
output(5, 221) <= input(28);
output(5, 222) <= input(29);
output(5, 223) <= input(30);
output(5, 224) <= input(35);
output(5, 225) <= input(16);
output(5, 226) <= input(17);
output(5, 227) <= input(18);
output(5, 228) <= input(19);
output(5, 229) <= input(20);
output(5, 230) <= input(21);
output(5, 231) <= input(22);
output(5, 232) <= input(23);
output(5, 233) <= input(24);
output(5, 234) <= input(25);
output(5, 235) <= input(26);
output(5, 236) <= input(27);
output(5, 237) <= input(28);
output(5, 238) <= input(29);
output(5, 239) <= input(30);
output(5, 240) <= input(35);
output(5, 241) <= input(16);
output(5, 242) <= input(17);
output(5, 243) <= input(18);
output(5, 244) <= input(19);
output(5, 245) <= input(20);
output(5, 246) <= input(21);
output(5, 247) <= input(22);
output(5, 248) <= input(23);
output(5, 249) <= input(24);
output(5, 250) <= input(25);
output(5, 251) <= input(26);
output(5, 252) <= input(27);
output(5, 253) <= input(28);
output(5, 254) <= input(29);
output(5, 255) <= input(30);
output(6, 0) <= input(35);
output(6, 1) <= input(16);
output(6, 2) <= input(17);
output(6, 3) <= input(18);
output(6, 4) <= input(19);
output(6, 5) <= input(20);
output(6, 6) <= input(21);
output(6, 7) <= input(22);
output(6, 8) <= input(23);
output(6, 9) <= input(24);
output(6, 10) <= input(25);
output(6, 11) <= input(26);
output(6, 12) <= input(27);
output(6, 13) <= input(28);
output(6, 14) <= input(29);
output(6, 15) <= input(30);
output(6, 16) <= input(35);
output(6, 17) <= input(16);
output(6, 18) <= input(17);
output(6, 19) <= input(18);
output(6, 20) <= input(19);
output(6, 21) <= input(20);
output(6, 22) <= input(21);
output(6, 23) <= input(22);
output(6, 24) <= input(23);
output(6, 25) <= input(24);
output(6, 26) <= input(25);
output(6, 27) <= input(26);
output(6, 28) <= input(27);
output(6, 29) <= input(28);
output(6, 30) <= input(29);
output(6, 31) <= input(30);
output(6, 32) <= input(35);
output(6, 33) <= input(16);
output(6, 34) <= input(17);
output(6, 35) <= input(18);
output(6, 36) <= input(19);
output(6, 37) <= input(20);
output(6, 38) <= input(21);
output(6, 39) <= input(22);
output(6, 40) <= input(23);
output(6, 41) <= input(24);
output(6, 42) <= input(25);
output(6, 43) <= input(26);
output(6, 44) <= input(27);
output(6, 45) <= input(28);
output(6, 46) <= input(29);
output(6, 47) <= input(30);
output(6, 48) <= input(35);
output(6, 49) <= input(16);
output(6, 50) <= input(17);
output(6, 51) <= input(18);
output(6, 52) <= input(19);
output(6, 53) <= input(20);
output(6, 54) <= input(21);
output(6, 55) <= input(22);
output(6, 56) <= input(23);
output(6, 57) <= input(24);
output(6, 58) <= input(25);
output(6, 59) <= input(26);
output(6, 60) <= input(27);
output(6, 61) <= input(28);
output(6, 62) <= input(29);
output(6, 63) <= input(30);
output(6, 64) <= input(35);
output(6, 65) <= input(16);
output(6, 66) <= input(17);
output(6, 67) <= input(18);
output(6, 68) <= input(19);
output(6, 69) <= input(20);
output(6, 70) <= input(21);
output(6, 71) <= input(22);
output(6, 72) <= input(23);
output(6, 73) <= input(24);
output(6, 74) <= input(25);
output(6, 75) <= input(26);
output(6, 76) <= input(27);
output(6, 77) <= input(28);
output(6, 78) <= input(29);
output(6, 79) <= input(30);
output(6, 80) <= input(35);
output(6, 81) <= input(16);
output(6, 82) <= input(17);
output(6, 83) <= input(18);
output(6, 84) <= input(19);
output(6, 85) <= input(20);
output(6, 86) <= input(21);
output(6, 87) <= input(22);
output(6, 88) <= input(23);
output(6, 89) <= input(24);
output(6, 90) <= input(25);
output(6, 91) <= input(26);
output(6, 92) <= input(27);
output(6, 93) <= input(28);
output(6, 94) <= input(29);
output(6, 95) <= input(30);
output(6, 96) <= input(35);
output(6, 97) <= input(16);
output(6, 98) <= input(17);
output(6, 99) <= input(18);
output(6, 100) <= input(19);
output(6, 101) <= input(20);
output(6, 102) <= input(21);
output(6, 103) <= input(22);
output(6, 104) <= input(23);
output(6, 105) <= input(24);
output(6, 106) <= input(25);
output(6, 107) <= input(26);
output(6, 108) <= input(27);
output(6, 109) <= input(28);
output(6, 110) <= input(29);
output(6, 111) <= input(30);
output(6, 112) <= input(35);
output(6, 113) <= input(16);
output(6, 114) <= input(17);
output(6, 115) <= input(18);
output(6, 116) <= input(19);
output(6, 117) <= input(20);
output(6, 118) <= input(21);
output(6, 119) <= input(22);
output(6, 120) <= input(23);
output(6, 121) <= input(24);
output(6, 122) <= input(25);
output(6, 123) <= input(26);
output(6, 124) <= input(27);
output(6, 125) <= input(28);
output(6, 126) <= input(29);
output(6, 127) <= input(30);
output(6, 128) <= input(36);
output(6, 129) <= input(0);
output(6, 130) <= input(1);
output(6, 131) <= input(2);
output(6, 132) <= input(3);
output(6, 133) <= input(4);
output(6, 134) <= input(5);
output(6, 135) <= input(6);
output(6, 136) <= input(7);
output(6, 137) <= input(8);
output(6, 138) <= input(9);
output(6, 139) <= input(10);
output(6, 140) <= input(11);
output(6, 141) <= input(12);
output(6, 142) <= input(13);
output(6, 143) <= input(14);
output(6, 144) <= input(36);
output(6, 145) <= input(0);
output(6, 146) <= input(1);
output(6, 147) <= input(2);
output(6, 148) <= input(3);
output(6, 149) <= input(4);
output(6, 150) <= input(5);
output(6, 151) <= input(6);
output(6, 152) <= input(7);
output(6, 153) <= input(8);
output(6, 154) <= input(9);
output(6, 155) <= input(10);
output(6, 156) <= input(11);
output(6, 157) <= input(12);
output(6, 158) <= input(13);
output(6, 159) <= input(14);
output(6, 160) <= input(36);
output(6, 161) <= input(0);
output(6, 162) <= input(1);
output(6, 163) <= input(2);
output(6, 164) <= input(3);
output(6, 165) <= input(4);
output(6, 166) <= input(5);
output(6, 167) <= input(6);
output(6, 168) <= input(7);
output(6, 169) <= input(8);
output(6, 170) <= input(9);
output(6, 171) <= input(10);
output(6, 172) <= input(11);
output(6, 173) <= input(12);
output(6, 174) <= input(13);
output(6, 175) <= input(14);
output(6, 176) <= input(36);
output(6, 177) <= input(0);
output(6, 178) <= input(1);
output(6, 179) <= input(2);
output(6, 180) <= input(3);
output(6, 181) <= input(4);
output(6, 182) <= input(5);
output(6, 183) <= input(6);
output(6, 184) <= input(7);
output(6, 185) <= input(8);
output(6, 186) <= input(9);
output(6, 187) <= input(10);
output(6, 188) <= input(11);
output(6, 189) <= input(12);
output(6, 190) <= input(13);
output(6, 191) <= input(14);
output(6, 192) <= input(36);
output(6, 193) <= input(0);
output(6, 194) <= input(1);
output(6, 195) <= input(2);
output(6, 196) <= input(3);
output(6, 197) <= input(4);
output(6, 198) <= input(5);
output(6, 199) <= input(6);
output(6, 200) <= input(7);
output(6, 201) <= input(8);
output(6, 202) <= input(9);
output(6, 203) <= input(10);
output(6, 204) <= input(11);
output(6, 205) <= input(12);
output(6, 206) <= input(13);
output(6, 207) <= input(14);
output(6, 208) <= input(36);
output(6, 209) <= input(0);
output(6, 210) <= input(1);
output(6, 211) <= input(2);
output(6, 212) <= input(3);
output(6, 213) <= input(4);
output(6, 214) <= input(5);
output(6, 215) <= input(6);
output(6, 216) <= input(7);
output(6, 217) <= input(8);
output(6, 218) <= input(9);
output(6, 219) <= input(10);
output(6, 220) <= input(11);
output(6, 221) <= input(12);
output(6, 222) <= input(13);
output(6, 223) <= input(14);
output(6, 224) <= input(36);
output(6, 225) <= input(0);
output(6, 226) <= input(1);
output(6, 227) <= input(2);
output(6, 228) <= input(3);
output(6, 229) <= input(4);
output(6, 230) <= input(5);
output(6, 231) <= input(6);
output(6, 232) <= input(7);
output(6, 233) <= input(8);
output(6, 234) <= input(9);
output(6, 235) <= input(10);
output(6, 236) <= input(11);
output(6, 237) <= input(12);
output(6, 238) <= input(13);
output(6, 239) <= input(14);
output(6, 240) <= input(36);
output(6, 241) <= input(0);
output(6, 242) <= input(1);
output(6, 243) <= input(2);
output(6, 244) <= input(3);
output(6, 245) <= input(4);
output(6, 246) <= input(5);
output(6, 247) <= input(6);
output(6, 248) <= input(7);
output(6, 249) <= input(8);
output(6, 250) <= input(9);
output(6, 251) <= input(10);
output(6, 252) <= input(11);
output(6, 253) <= input(12);
output(6, 254) <= input(13);
output(6, 255) <= input(14);
output(7, 0) <= input(35);
output(7, 1) <= input(16);
output(7, 2) <= input(17);
output(7, 3) <= input(18);
output(7, 4) <= input(19);
output(7, 5) <= input(20);
output(7, 6) <= input(21);
output(7, 7) <= input(22);
output(7, 8) <= input(23);
output(7, 9) <= input(24);
output(7, 10) <= input(25);
output(7, 11) <= input(26);
output(7, 12) <= input(27);
output(7, 13) <= input(28);
output(7, 14) <= input(29);
output(7, 15) <= input(30);
output(7, 16) <= input(35);
output(7, 17) <= input(16);
output(7, 18) <= input(17);
output(7, 19) <= input(18);
output(7, 20) <= input(19);
output(7, 21) <= input(20);
output(7, 22) <= input(21);
output(7, 23) <= input(22);
output(7, 24) <= input(23);
output(7, 25) <= input(24);
output(7, 26) <= input(25);
output(7, 27) <= input(26);
output(7, 28) <= input(27);
output(7, 29) <= input(28);
output(7, 30) <= input(29);
output(7, 31) <= input(30);
output(7, 32) <= input(35);
output(7, 33) <= input(16);
output(7, 34) <= input(17);
output(7, 35) <= input(18);
output(7, 36) <= input(19);
output(7, 37) <= input(20);
output(7, 38) <= input(21);
output(7, 39) <= input(22);
output(7, 40) <= input(23);
output(7, 41) <= input(24);
output(7, 42) <= input(25);
output(7, 43) <= input(26);
output(7, 44) <= input(27);
output(7, 45) <= input(28);
output(7, 46) <= input(29);
output(7, 47) <= input(30);
output(7, 48) <= input(35);
output(7, 49) <= input(16);
output(7, 50) <= input(17);
output(7, 51) <= input(18);
output(7, 52) <= input(19);
output(7, 53) <= input(20);
output(7, 54) <= input(21);
output(7, 55) <= input(22);
output(7, 56) <= input(23);
output(7, 57) <= input(24);
output(7, 58) <= input(25);
output(7, 59) <= input(26);
output(7, 60) <= input(27);
output(7, 61) <= input(28);
output(7, 62) <= input(29);
output(7, 63) <= input(30);
output(7, 64) <= input(35);
output(7, 65) <= input(16);
output(7, 66) <= input(17);
output(7, 67) <= input(18);
output(7, 68) <= input(19);
output(7, 69) <= input(20);
output(7, 70) <= input(21);
output(7, 71) <= input(22);
output(7, 72) <= input(23);
output(7, 73) <= input(24);
output(7, 74) <= input(25);
output(7, 75) <= input(26);
output(7, 76) <= input(27);
output(7, 77) <= input(28);
output(7, 78) <= input(29);
output(7, 79) <= input(30);
output(7, 80) <= input(36);
output(7, 81) <= input(0);
output(7, 82) <= input(1);
output(7, 83) <= input(2);
output(7, 84) <= input(3);
output(7, 85) <= input(4);
output(7, 86) <= input(5);
output(7, 87) <= input(6);
output(7, 88) <= input(7);
output(7, 89) <= input(8);
output(7, 90) <= input(9);
output(7, 91) <= input(10);
output(7, 92) <= input(11);
output(7, 93) <= input(12);
output(7, 94) <= input(13);
output(7, 95) <= input(14);
output(7, 96) <= input(36);
output(7, 97) <= input(0);
output(7, 98) <= input(1);
output(7, 99) <= input(2);
output(7, 100) <= input(3);
output(7, 101) <= input(4);
output(7, 102) <= input(5);
output(7, 103) <= input(6);
output(7, 104) <= input(7);
output(7, 105) <= input(8);
output(7, 106) <= input(9);
output(7, 107) <= input(10);
output(7, 108) <= input(11);
output(7, 109) <= input(12);
output(7, 110) <= input(13);
output(7, 111) <= input(14);
output(7, 112) <= input(36);
output(7, 113) <= input(0);
output(7, 114) <= input(1);
output(7, 115) <= input(2);
output(7, 116) <= input(3);
output(7, 117) <= input(4);
output(7, 118) <= input(5);
output(7, 119) <= input(6);
output(7, 120) <= input(7);
output(7, 121) <= input(8);
output(7, 122) <= input(9);
output(7, 123) <= input(10);
output(7, 124) <= input(11);
output(7, 125) <= input(12);
output(7, 126) <= input(13);
output(7, 127) <= input(14);
output(7, 128) <= input(36);
output(7, 129) <= input(0);
output(7, 130) <= input(1);
output(7, 131) <= input(2);
output(7, 132) <= input(3);
output(7, 133) <= input(4);
output(7, 134) <= input(5);
output(7, 135) <= input(6);
output(7, 136) <= input(7);
output(7, 137) <= input(8);
output(7, 138) <= input(9);
output(7, 139) <= input(10);
output(7, 140) <= input(11);
output(7, 141) <= input(12);
output(7, 142) <= input(13);
output(7, 143) <= input(14);
output(7, 144) <= input(36);
output(7, 145) <= input(0);
output(7, 146) <= input(1);
output(7, 147) <= input(2);
output(7, 148) <= input(3);
output(7, 149) <= input(4);
output(7, 150) <= input(5);
output(7, 151) <= input(6);
output(7, 152) <= input(7);
output(7, 153) <= input(8);
output(7, 154) <= input(9);
output(7, 155) <= input(10);
output(7, 156) <= input(11);
output(7, 157) <= input(12);
output(7, 158) <= input(13);
output(7, 159) <= input(14);
output(7, 160) <= input(37);
output(7, 161) <= input(35);
output(7, 162) <= input(16);
output(7, 163) <= input(17);
output(7, 164) <= input(18);
output(7, 165) <= input(19);
output(7, 166) <= input(20);
output(7, 167) <= input(21);
output(7, 168) <= input(22);
output(7, 169) <= input(23);
output(7, 170) <= input(24);
output(7, 171) <= input(25);
output(7, 172) <= input(26);
output(7, 173) <= input(27);
output(7, 174) <= input(28);
output(7, 175) <= input(29);
output(7, 176) <= input(37);
output(7, 177) <= input(35);
output(7, 178) <= input(16);
output(7, 179) <= input(17);
output(7, 180) <= input(18);
output(7, 181) <= input(19);
output(7, 182) <= input(20);
output(7, 183) <= input(21);
output(7, 184) <= input(22);
output(7, 185) <= input(23);
output(7, 186) <= input(24);
output(7, 187) <= input(25);
output(7, 188) <= input(26);
output(7, 189) <= input(27);
output(7, 190) <= input(28);
output(7, 191) <= input(29);
output(7, 192) <= input(37);
output(7, 193) <= input(35);
output(7, 194) <= input(16);
output(7, 195) <= input(17);
output(7, 196) <= input(18);
output(7, 197) <= input(19);
output(7, 198) <= input(20);
output(7, 199) <= input(21);
output(7, 200) <= input(22);
output(7, 201) <= input(23);
output(7, 202) <= input(24);
output(7, 203) <= input(25);
output(7, 204) <= input(26);
output(7, 205) <= input(27);
output(7, 206) <= input(28);
output(7, 207) <= input(29);
output(7, 208) <= input(37);
output(7, 209) <= input(35);
output(7, 210) <= input(16);
output(7, 211) <= input(17);
output(7, 212) <= input(18);
output(7, 213) <= input(19);
output(7, 214) <= input(20);
output(7, 215) <= input(21);
output(7, 216) <= input(22);
output(7, 217) <= input(23);
output(7, 218) <= input(24);
output(7, 219) <= input(25);
output(7, 220) <= input(26);
output(7, 221) <= input(27);
output(7, 222) <= input(28);
output(7, 223) <= input(29);
output(7, 224) <= input(37);
output(7, 225) <= input(35);
output(7, 226) <= input(16);
output(7, 227) <= input(17);
output(7, 228) <= input(18);
output(7, 229) <= input(19);
output(7, 230) <= input(20);
output(7, 231) <= input(21);
output(7, 232) <= input(22);
output(7, 233) <= input(23);
output(7, 234) <= input(24);
output(7, 235) <= input(25);
output(7, 236) <= input(26);
output(7, 237) <= input(27);
output(7, 238) <= input(28);
output(7, 239) <= input(29);
output(7, 240) <= input(37);
output(7, 241) <= input(35);
output(7, 242) <= input(16);
output(7, 243) <= input(17);
output(7, 244) <= input(18);
output(7, 245) <= input(19);
output(7, 246) <= input(20);
output(7, 247) <= input(21);
output(7, 248) <= input(22);
output(7, 249) <= input(23);
output(7, 250) <= input(24);
output(7, 251) <= input(25);
output(7, 252) <= input(26);
output(7, 253) <= input(27);
output(7, 254) <= input(28);
output(7, 255) <= input(29);
when "0011" =>
output(0, 0) <= input(0);
output(0, 1) <= input(1);
output(0, 2) <= input(2);
output(0, 3) <= input(3);
output(0, 4) <= input(4);
output(0, 5) <= input(5);
output(0, 6) <= input(6);
output(0, 7) <= input(7);
output(0, 8) <= input(8);
output(0, 9) <= input(9);
output(0, 10) <= input(10);
output(0, 11) <= input(11);
output(0, 12) <= input(12);
output(0, 13) <= input(13);
output(0, 14) <= input(14);
output(0, 15) <= input(15);
output(0, 16) <= input(0);
output(0, 17) <= input(1);
output(0, 18) <= input(2);
output(0, 19) <= input(3);
output(0, 20) <= input(4);
output(0, 21) <= input(5);
output(0, 22) <= input(6);
output(0, 23) <= input(7);
output(0, 24) <= input(8);
output(0, 25) <= input(9);
output(0, 26) <= input(10);
output(0, 27) <= input(11);
output(0, 28) <= input(12);
output(0, 29) <= input(13);
output(0, 30) <= input(14);
output(0, 31) <= input(15);
output(0, 32) <= input(0);
output(0, 33) <= input(1);
output(0, 34) <= input(2);
output(0, 35) <= input(3);
output(0, 36) <= input(4);
output(0, 37) <= input(5);
output(0, 38) <= input(6);
output(0, 39) <= input(7);
output(0, 40) <= input(8);
output(0, 41) <= input(9);
output(0, 42) <= input(10);
output(0, 43) <= input(11);
output(0, 44) <= input(12);
output(0, 45) <= input(13);
output(0, 46) <= input(14);
output(0, 47) <= input(15);
output(0, 48) <= input(0);
output(0, 49) <= input(1);
output(0, 50) <= input(2);
output(0, 51) <= input(3);
output(0, 52) <= input(4);
output(0, 53) <= input(5);
output(0, 54) <= input(6);
output(0, 55) <= input(7);
output(0, 56) <= input(8);
output(0, 57) <= input(9);
output(0, 58) <= input(10);
output(0, 59) <= input(11);
output(0, 60) <= input(12);
output(0, 61) <= input(13);
output(0, 62) <= input(14);
output(0, 63) <= input(15);
output(0, 64) <= input(16);
output(0, 65) <= input(17);
output(0, 66) <= input(18);
output(0, 67) <= input(19);
output(0, 68) <= input(20);
output(0, 69) <= input(21);
output(0, 70) <= input(22);
output(0, 71) <= input(23);
output(0, 72) <= input(24);
output(0, 73) <= input(25);
output(0, 74) <= input(26);
output(0, 75) <= input(27);
output(0, 76) <= input(28);
output(0, 77) <= input(29);
output(0, 78) <= input(30);
output(0, 79) <= input(31);
output(0, 80) <= input(16);
output(0, 81) <= input(17);
output(0, 82) <= input(18);
output(0, 83) <= input(19);
output(0, 84) <= input(20);
output(0, 85) <= input(21);
output(0, 86) <= input(22);
output(0, 87) <= input(23);
output(0, 88) <= input(24);
output(0, 89) <= input(25);
output(0, 90) <= input(26);
output(0, 91) <= input(27);
output(0, 92) <= input(28);
output(0, 93) <= input(29);
output(0, 94) <= input(30);
output(0, 95) <= input(31);
output(0, 96) <= input(16);
output(0, 97) <= input(17);
output(0, 98) <= input(18);
output(0, 99) <= input(19);
output(0, 100) <= input(20);
output(0, 101) <= input(21);
output(0, 102) <= input(22);
output(0, 103) <= input(23);
output(0, 104) <= input(24);
output(0, 105) <= input(25);
output(0, 106) <= input(26);
output(0, 107) <= input(27);
output(0, 108) <= input(28);
output(0, 109) <= input(29);
output(0, 110) <= input(30);
output(0, 111) <= input(31);
output(0, 112) <= input(16);
output(0, 113) <= input(17);
output(0, 114) <= input(18);
output(0, 115) <= input(19);
output(0, 116) <= input(20);
output(0, 117) <= input(21);
output(0, 118) <= input(22);
output(0, 119) <= input(23);
output(0, 120) <= input(24);
output(0, 121) <= input(25);
output(0, 122) <= input(26);
output(0, 123) <= input(27);
output(0, 124) <= input(28);
output(0, 125) <= input(29);
output(0, 126) <= input(30);
output(0, 127) <= input(31);
output(0, 128) <= input(32);
output(0, 129) <= input(0);
output(0, 130) <= input(1);
output(0, 131) <= input(2);
output(0, 132) <= input(3);
output(0, 133) <= input(4);
output(0, 134) <= input(5);
output(0, 135) <= input(6);
output(0, 136) <= input(7);
output(0, 137) <= input(8);
output(0, 138) <= input(9);
output(0, 139) <= input(10);
output(0, 140) <= input(11);
output(0, 141) <= input(12);
output(0, 142) <= input(13);
output(0, 143) <= input(14);
output(0, 144) <= input(32);
output(0, 145) <= input(0);
output(0, 146) <= input(1);
output(0, 147) <= input(2);
output(0, 148) <= input(3);
output(0, 149) <= input(4);
output(0, 150) <= input(5);
output(0, 151) <= input(6);
output(0, 152) <= input(7);
output(0, 153) <= input(8);
output(0, 154) <= input(9);
output(0, 155) <= input(10);
output(0, 156) <= input(11);
output(0, 157) <= input(12);
output(0, 158) <= input(13);
output(0, 159) <= input(14);
output(0, 160) <= input(32);
output(0, 161) <= input(0);
output(0, 162) <= input(1);
output(0, 163) <= input(2);
output(0, 164) <= input(3);
output(0, 165) <= input(4);
output(0, 166) <= input(5);
output(0, 167) <= input(6);
output(0, 168) <= input(7);
output(0, 169) <= input(8);
output(0, 170) <= input(9);
output(0, 171) <= input(10);
output(0, 172) <= input(11);
output(0, 173) <= input(12);
output(0, 174) <= input(13);
output(0, 175) <= input(14);
output(0, 176) <= input(32);
output(0, 177) <= input(0);
output(0, 178) <= input(1);
output(0, 179) <= input(2);
output(0, 180) <= input(3);
output(0, 181) <= input(4);
output(0, 182) <= input(5);
output(0, 183) <= input(6);
output(0, 184) <= input(7);
output(0, 185) <= input(8);
output(0, 186) <= input(9);
output(0, 187) <= input(10);
output(0, 188) <= input(11);
output(0, 189) <= input(12);
output(0, 190) <= input(13);
output(0, 191) <= input(14);
output(0, 192) <= input(33);
output(0, 193) <= input(16);
output(0, 194) <= input(17);
output(0, 195) <= input(18);
output(0, 196) <= input(19);
output(0, 197) <= input(20);
output(0, 198) <= input(21);
output(0, 199) <= input(22);
output(0, 200) <= input(23);
output(0, 201) <= input(24);
output(0, 202) <= input(25);
output(0, 203) <= input(26);
output(0, 204) <= input(27);
output(0, 205) <= input(28);
output(0, 206) <= input(29);
output(0, 207) <= input(30);
output(0, 208) <= input(33);
output(0, 209) <= input(16);
output(0, 210) <= input(17);
output(0, 211) <= input(18);
output(0, 212) <= input(19);
output(0, 213) <= input(20);
output(0, 214) <= input(21);
output(0, 215) <= input(22);
output(0, 216) <= input(23);
output(0, 217) <= input(24);
output(0, 218) <= input(25);
output(0, 219) <= input(26);
output(0, 220) <= input(27);
output(0, 221) <= input(28);
output(0, 222) <= input(29);
output(0, 223) <= input(30);
output(0, 224) <= input(33);
output(0, 225) <= input(16);
output(0, 226) <= input(17);
output(0, 227) <= input(18);
output(0, 228) <= input(19);
output(0, 229) <= input(20);
output(0, 230) <= input(21);
output(0, 231) <= input(22);
output(0, 232) <= input(23);
output(0, 233) <= input(24);
output(0, 234) <= input(25);
output(0, 235) <= input(26);
output(0, 236) <= input(27);
output(0, 237) <= input(28);
output(0, 238) <= input(29);
output(0, 239) <= input(30);
output(0, 240) <= input(33);
output(0, 241) <= input(16);
output(0, 242) <= input(17);
output(0, 243) <= input(18);
output(0, 244) <= input(19);
output(0, 245) <= input(20);
output(0, 246) <= input(21);
output(0, 247) <= input(22);
output(0, 248) <= input(23);
output(0, 249) <= input(24);
output(0, 250) <= input(25);
output(0, 251) <= input(26);
output(0, 252) <= input(27);
output(0, 253) <= input(28);
output(0, 254) <= input(29);
output(0, 255) <= input(30);
output(1, 0) <= input(0);
output(1, 1) <= input(1);
output(1, 2) <= input(2);
output(1, 3) <= input(3);
output(1, 4) <= input(4);
output(1, 5) <= input(5);
output(1, 6) <= input(6);
output(1, 7) <= input(7);
output(1, 8) <= input(8);
output(1, 9) <= input(9);
output(1, 10) <= input(10);
output(1, 11) <= input(11);
output(1, 12) <= input(12);
output(1, 13) <= input(13);
output(1, 14) <= input(14);
output(1, 15) <= input(15);
output(1, 16) <= input(0);
output(1, 17) <= input(1);
output(1, 18) <= input(2);
output(1, 19) <= input(3);
output(1, 20) <= input(4);
output(1, 21) <= input(5);
output(1, 22) <= input(6);
output(1, 23) <= input(7);
output(1, 24) <= input(8);
output(1, 25) <= input(9);
output(1, 26) <= input(10);
output(1, 27) <= input(11);
output(1, 28) <= input(12);
output(1, 29) <= input(13);
output(1, 30) <= input(14);
output(1, 31) <= input(15);
output(1, 32) <= input(16);
output(1, 33) <= input(17);
output(1, 34) <= input(18);
output(1, 35) <= input(19);
output(1, 36) <= input(20);
output(1, 37) <= input(21);
output(1, 38) <= input(22);
output(1, 39) <= input(23);
output(1, 40) <= input(24);
output(1, 41) <= input(25);
output(1, 42) <= input(26);
output(1, 43) <= input(27);
output(1, 44) <= input(28);
output(1, 45) <= input(29);
output(1, 46) <= input(30);
output(1, 47) <= input(31);
output(1, 48) <= input(16);
output(1, 49) <= input(17);
output(1, 50) <= input(18);
output(1, 51) <= input(19);
output(1, 52) <= input(20);
output(1, 53) <= input(21);
output(1, 54) <= input(22);
output(1, 55) <= input(23);
output(1, 56) <= input(24);
output(1, 57) <= input(25);
output(1, 58) <= input(26);
output(1, 59) <= input(27);
output(1, 60) <= input(28);
output(1, 61) <= input(29);
output(1, 62) <= input(30);
output(1, 63) <= input(31);
output(1, 64) <= input(16);
output(1, 65) <= input(17);
output(1, 66) <= input(18);
output(1, 67) <= input(19);
output(1, 68) <= input(20);
output(1, 69) <= input(21);
output(1, 70) <= input(22);
output(1, 71) <= input(23);
output(1, 72) <= input(24);
output(1, 73) <= input(25);
output(1, 74) <= input(26);
output(1, 75) <= input(27);
output(1, 76) <= input(28);
output(1, 77) <= input(29);
output(1, 78) <= input(30);
output(1, 79) <= input(31);
output(1, 80) <= input(32);
output(1, 81) <= input(0);
output(1, 82) <= input(1);
output(1, 83) <= input(2);
output(1, 84) <= input(3);
output(1, 85) <= input(4);
output(1, 86) <= input(5);
output(1, 87) <= input(6);
output(1, 88) <= input(7);
output(1, 89) <= input(8);
output(1, 90) <= input(9);
output(1, 91) <= input(10);
output(1, 92) <= input(11);
output(1, 93) <= input(12);
output(1, 94) <= input(13);
output(1, 95) <= input(14);
output(1, 96) <= input(32);
output(1, 97) <= input(0);
output(1, 98) <= input(1);
output(1, 99) <= input(2);
output(1, 100) <= input(3);
output(1, 101) <= input(4);
output(1, 102) <= input(5);
output(1, 103) <= input(6);
output(1, 104) <= input(7);
output(1, 105) <= input(8);
output(1, 106) <= input(9);
output(1, 107) <= input(10);
output(1, 108) <= input(11);
output(1, 109) <= input(12);
output(1, 110) <= input(13);
output(1, 111) <= input(14);
output(1, 112) <= input(32);
output(1, 113) <= input(0);
output(1, 114) <= input(1);
output(1, 115) <= input(2);
output(1, 116) <= input(3);
output(1, 117) <= input(4);
output(1, 118) <= input(5);
output(1, 119) <= input(6);
output(1, 120) <= input(7);
output(1, 121) <= input(8);
output(1, 122) <= input(9);
output(1, 123) <= input(10);
output(1, 124) <= input(11);
output(1, 125) <= input(12);
output(1, 126) <= input(13);
output(1, 127) <= input(14);
output(1, 128) <= input(33);
output(1, 129) <= input(16);
output(1, 130) <= input(17);
output(1, 131) <= input(18);
output(1, 132) <= input(19);
output(1, 133) <= input(20);
output(1, 134) <= input(21);
output(1, 135) <= input(22);
output(1, 136) <= input(23);
output(1, 137) <= input(24);
output(1, 138) <= input(25);
output(1, 139) <= input(26);
output(1, 140) <= input(27);
output(1, 141) <= input(28);
output(1, 142) <= input(29);
output(1, 143) <= input(30);
output(1, 144) <= input(33);
output(1, 145) <= input(16);
output(1, 146) <= input(17);
output(1, 147) <= input(18);
output(1, 148) <= input(19);
output(1, 149) <= input(20);
output(1, 150) <= input(21);
output(1, 151) <= input(22);
output(1, 152) <= input(23);
output(1, 153) <= input(24);
output(1, 154) <= input(25);
output(1, 155) <= input(26);
output(1, 156) <= input(27);
output(1, 157) <= input(28);
output(1, 158) <= input(29);
output(1, 159) <= input(30);
output(1, 160) <= input(34);
output(1, 161) <= input(32);
output(1, 162) <= input(0);
output(1, 163) <= input(1);
output(1, 164) <= input(2);
output(1, 165) <= input(3);
output(1, 166) <= input(4);
output(1, 167) <= input(5);
output(1, 168) <= input(6);
output(1, 169) <= input(7);
output(1, 170) <= input(8);
output(1, 171) <= input(9);
output(1, 172) <= input(10);
output(1, 173) <= input(11);
output(1, 174) <= input(12);
output(1, 175) <= input(13);
output(1, 176) <= input(34);
output(1, 177) <= input(32);
output(1, 178) <= input(0);
output(1, 179) <= input(1);
output(1, 180) <= input(2);
output(1, 181) <= input(3);
output(1, 182) <= input(4);
output(1, 183) <= input(5);
output(1, 184) <= input(6);
output(1, 185) <= input(7);
output(1, 186) <= input(8);
output(1, 187) <= input(9);
output(1, 188) <= input(10);
output(1, 189) <= input(11);
output(1, 190) <= input(12);
output(1, 191) <= input(13);
output(1, 192) <= input(34);
output(1, 193) <= input(32);
output(1, 194) <= input(0);
output(1, 195) <= input(1);
output(1, 196) <= input(2);
output(1, 197) <= input(3);
output(1, 198) <= input(4);
output(1, 199) <= input(5);
output(1, 200) <= input(6);
output(1, 201) <= input(7);
output(1, 202) <= input(8);
output(1, 203) <= input(9);
output(1, 204) <= input(10);
output(1, 205) <= input(11);
output(1, 206) <= input(12);
output(1, 207) <= input(13);
output(1, 208) <= input(35);
output(1, 209) <= input(33);
output(1, 210) <= input(16);
output(1, 211) <= input(17);
output(1, 212) <= input(18);
output(1, 213) <= input(19);
output(1, 214) <= input(20);
output(1, 215) <= input(21);
output(1, 216) <= input(22);
output(1, 217) <= input(23);
output(1, 218) <= input(24);
output(1, 219) <= input(25);
output(1, 220) <= input(26);
output(1, 221) <= input(27);
output(1, 222) <= input(28);
output(1, 223) <= input(29);
output(1, 224) <= input(35);
output(1, 225) <= input(33);
output(1, 226) <= input(16);
output(1, 227) <= input(17);
output(1, 228) <= input(18);
output(1, 229) <= input(19);
output(1, 230) <= input(20);
output(1, 231) <= input(21);
output(1, 232) <= input(22);
output(1, 233) <= input(23);
output(1, 234) <= input(24);
output(1, 235) <= input(25);
output(1, 236) <= input(26);
output(1, 237) <= input(27);
output(1, 238) <= input(28);
output(1, 239) <= input(29);
output(1, 240) <= input(35);
output(1, 241) <= input(33);
output(1, 242) <= input(16);
output(1, 243) <= input(17);
output(1, 244) <= input(18);
output(1, 245) <= input(19);
output(1, 246) <= input(20);
output(1, 247) <= input(21);
output(1, 248) <= input(22);
output(1, 249) <= input(23);
output(1, 250) <= input(24);
output(1, 251) <= input(25);
output(1, 252) <= input(26);
output(1, 253) <= input(27);
output(1, 254) <= input(28);
output(1, 255) <= input(29);
output(2, 0) <= input(0);
output(2, 1) <= input(1);
output(2, 2) <= input(2);
output(2, 3) <= input(3);
output(2, 4) <= input(4);
output(2, 5) <= input(5);
output(2, 6) <= input(6);
output(2, 7) <= input(7);
output(2, 8) <= input(8);
output(2, 9) <= input(9);
output(2, 10) <= input(10);
output(2, 11) <= input(11);
output(2, 12) <= input(12);
output(2, 13) <= input(13);
output(2, 14) <= input(14);
output(2, 15) <= input(15);
output(2, 16) <= input(0);
output(2, 17) <= input(1);
output(2, 18) <= input(2);
output(2, 19) <= input(3);
output(2, 20) <= input(4);
output(2, 21) <= input(5);
output(2, 22) <= input(6);
output(2, 23) <= input(7);
output(2, 24) <= input(8);
output(2, 25) <= input(9);
output(2, 26) <= input(10);
output(2, 27) <= input(11);
output(2, 28) <= input(12);
output(2, 29) <= input(13);
output(2, 30) <= input(14);
output(2, 31) <= input(15);
output(2, 32) <= input(16);
output(2, 33) <= input(17);
output(2, 34) <= input(18);
output(2, 35) <= input(19);
output(2, 36) <= input(20);
output(2, 37) <= input(21);
output(2, 38) <= input(22);
output(2, 39) <= input(23);
output(2, 40) <= input(24);
output(2, 41) <= input(25);
output(2, 42) <= input(26);
output(2, 43) <= input(27);
output(2, 44) <= input(28);
output(2, 45) <= input(29);
output(2, 46) <= input(30);
output(2, 47) <= input(31);
output(2, 48) <= input(16);
output(2, 49) <= input(17);
output(2, 50) <= input(18);
output(2, 51) <= input(19);
output(2, 52) <= input(20);
output(2, 53) <= input(21);
output(2, 54) <= input(22);
output(2, 55) <= input(23);
output(2, 56) <= input(24);
output(2, 57) <= input(25);
output(2, 58) <= input(26);
output(2, 59) <= input(27);
output(2, 60) <= input(28);
output(2, 61) <= input(29);
output(2, 62) <= input(30);
output(2, 63) <= input(31);
output(2, 64) <= input(32);
output(2, 65) <= input(0);
output(2, 66) <= input(1);
output(2, 67) <= input(2);
output(2, 68) <= input(3);
output(2, 69) <= input(4);
output(2, 70) <= input(5);
output(2, 71) <= input(6);
output(2, 72) <= input(7);
output(2, 73) <= input(8);
output(2, 74) <= input(9);
output(2, 75) <= input(10);
output(2, 76) <= input(11);
output(2, 77) <= input(12);
output(2, 78) <= input(13);
output(2, 79) <= input(14);
output(2, 80) <= input(32);
output(2, 81) <= input(0);
output(2, 82) <= input(1);
output(2, 83) <= input(2);
output(2, 84) <= input(3);
output(2, 85) <= input(4);
output(2, 86) <= input(5);
output(2, 87) <= input(6);
output(2, 88) <= input(7);
output(2, 89) <= input(8);
output(2, 90) <= input(9);
output(2, 91) <= input(10);
output(2, 92) <= input(11);
output(2, 93) <= input(12);
output(2, 94) <= input(13);
output(2, 95) <= input(14);
output(2, 96) <= input(33);
output(2, 97) <= input(16);
output(2, 98) <= input(17);
output(2, 99) <= input(18);
output(2, 100) <= input(19);
output(2, 101) <= input(20);
output(2, 102) <= input(21);
output(2, 103) <= input(22);
output(2, 104) <= input(23);
output(2, 105) <= input(24);
output(2, 106) <= input(25);
output(2, 107) <= input(26);
output(2, 108) <= input(27);
output(2, 109) <= input(28);
output(2, 110) <= input(29);
output(2, 111) <= input(30);
output(2, 112) <= input(33);
output(2, 113) <= input(16);
output(2, 114) <= input(17);
output(2, 115) <= input(18);
output(2, 116) <= input(19);
output(2, 117) <= input(20);
output(2, 118) <= input(21);
output(2, 119) <= input(22);
output(2, 120) <= input(23);
output(2, 121) <= input(24);
output(2, 122) <= input(25);
output(2, 123) <= input(26);
output(2, 124) <= input(27);
output(2, 125) <= input(28);
output(2, 126) <= input(29);
output(2, 127) <= input(30);
output(2, 128) <= input(34);
output(2, 129) <= input(32);
output(2, 130) <= input(0);
output(2, 131) <= input(1);
output(2, 132) <= input(2);
output(2, 133) <= input(3);
output(2, 134) <= input(4);
output(2, 135) <= input(5);
output(2, 136) <= input(6);
output(2, 137) <= input(7);
output(2, 138) <= input(8);
output(2, 139) <= input(9);
output(2, 140) <= input(10);
output(2, 141) <= input(11);
output(2, 142) <= input(12);
output(2, 143) <= input(13);
output(2, 144) <= input(34);
output(2, 145) <= input(32);
output(2, 146) <= input(0);
output(2, 147) <= input(1);
output(2, 148) <= input(2);
output(2, 149) <= input(3);
output(2, 150) <= input(4);
output(2, 151) <= input(5);
output(2, 152) <= input(6);
output(2, 153) <= input(7);
output(2, 154) <= input(8);
output(2, 155) <= input(9);
output(2, 156) <= input(10);
output(2, 157) <= input(11);
output(2, 158) <= input(12);
output(2, 159) <= input(13);
output(2, 160) <= input(35);
output(2, 161) <= input(33);
output(2, 162) <= input(16);
output(2, 163) <= input(17);
output(2, 164) <= input(18);
output(2, 165) <= input(19);
output(2, 166) <= input(20);
output(2, 167) <= input(21);
output(2, 168) <= input(22);
output(2, 169) <= input(23);
output(2, 170) <= input(24);
output(2, 171) <= input(25);
output(2, 172) <= input(26);
output(2, 173) <= input(27);
output(2, 174) <= input(28);
output(2, 175) <= input(29);
output(2, 176) <= input(35);
output(2, 177) <= input(33);
output(2, 178) <= input(16);
output(2, 179) <= input(17);
output(2, 180) <= input(18);
output(2, 181) <= input(19);
output(2, 182) <= input(20);
output(2, 183) <= input(21);
output(2, 184) <= input(22);
output(2, 185) <= input(23);
output(2, 186) <= input(24);
output(2, 187) <= input(25);
output(2, 188) <= input(26);
output(2, 189) <= input(27);
output(2, 190) <= input(28);
output(2, 191) <= input(29);
output(2, 192) <= input(36);
output(2, 193) <= input(34);
output(2, 194) <= input(32);
output(2, 195) <= input(0);
output(2, 196) <= input(1);
output(2, 197) <= input(2);
output(2, 198) <= input(3);
output(2, 199) <= input(4);
output(2, 200) <= input(5);
output(2, 201) <= input(6);
output(2, 202) <= input(7);
output(2, 203) <= input(8);
output(2, 204) <= input(9);
output(2, 205) <= input(10);
output(2, 206) <= input(11);
output(2, 207) <= input(12);
output(2, 208) <= input(36);
output(2, 209) <= input(34);
output(2, 210) <= input(32);
output(2, 211) <= input(0);
output(2, 212) <= input(1);
output(2, 213) <= input(2);
output(2, 214) <= input(3);
output(2, 215) <= input(4);
output(2, 216) <= input(5);
output(2, 217) <= input(6);
output(2, 218) <= input(7);
output(2, 219) <= input(8);
output(2, 220) <= input(9);
output(2, 221) <= input(10);
output(2, 222) <= input(11);
output(2, 223) <= input(12);
output(2, 224) <= input(37);
output(2, 225) <= input(35);
output(2, 226) <= input(33);
output(2, 227) <= input(16);
output(2, 228) <= input(17);
output(2, 229) <= input(18);
output(2, 230) <= input(19);
output(2, 231) <= input(20);
output(2, 232) <= input(21);
output(2, 233) <= input(22);
output(2, 234) <= input(23);
output(2, 235) <= input(24);
output(2, 236) <= input(25);
output(2, 237) <= input(26);
output(2, 238) <= input(27);
output(2, 239) <= input(28);
output(2, 240) <= input(37);
output(2, 241) <= input(35);
output(2, 242) <= input(33);
output(2, 243) <= input(16);
output(2, 244) <= input(17);
output(2, 245) <= input(18);
output(2, 246) <= input(19);
output(2, 247) <= input(20);
output(2, 248) <= input(21);
output(2, 249) <= input(22);
output(2, 250) <= input(23);
output(2, 251) <= input(24);
output(2, 252) <= input(25);
output(2, 253) <= input(26);
output(2, 254) <= input(27);
output(2, 255) <= input(28);
when "0100" =>
output(0, 0) <= input(0);
output(0, 1) <= input(1);
output(0, 2) <= input(2);
output(0, 3) <= input(3);
output(0, 4) <= input(4);
output(0, 5) <= input(5);
output(0, 6) <= input(6);
output(0, 7) <= input(7);
output(0, 8) <= input(8);
output(0, 9) <= input(9);
output(0, 10) <= input(10);
output(0, 11) <= input(11);
output(0, 12) <= input(12);
output(0, 13) <= input(13);
output(0, 14) <= input(14);
output(0, 15) <= input(15);
output(0, 16) <= input(16);
output(0, 17) <= input(17);
output(0, 18) <= input(18);
output(0, 19) <= input(19);
output(0, 20) <= input(20);
output(0, 21) <= input(21);
output(0, 22) <= input(22);
output(0, 23) <= input(23);
output(0, 24) <= input(24);
output(0, 25) <= input(25);
output(0, 26) <= input(26);
output(0, 27) <= input(27);
output(0, 28) <= input(28);
output(0, 29) <= input(29);
output(0, 30) <= input(30);
output(0, 31) <= input(31);
output(0, 32) <= input(16);
output(0, 33) <= input(17);
output(0, 34) <= input(18);
output(0, 35) <= input(19);
output(0, 36) <= input(20);
output(0, 37) <= input(21);
output(0, 38) <= input(22);
output(0, 39) <= input(23);
output(0, 40) <= input(24);
output(0, 41) <= input(25);
output(0, 42) <= input(26);
output(0, 43) <= input(27);
output(0, 44) <= input(28);
output(0, 45) <= input(29);
output(0, 46) <= input(30);
output(0, 47) <= input(31);
output(0, 48) <= input(32);
output(0, 49) <= input(0);
output(0, 50) <= input(1);
output(0, 51) <= input(2);
output(0, 52) <= input(3);
output(0, 53) <= input(4);
output(0, 54) <= input(5);
output(0, 55) <= input(6);
output(0, 56) <= input(7);
output(0, 57) <= input(8);
output(0, 58) <= input(9);
output(0, 59) <= input(10);
output(0, 60) <= input(11);
output(0, 61) <= input(12);
output(0, 62) <= input(13);
output(0, 63) <= input(14);
output(0, 64) <= input(33);
output(0, 65) <= input(16);
output(0, 66) <= input(17);
output(0, 67) <= input(18);
output(0, 68) <= input(19);
output(0, 69) <= input(20);
output(0, 70) <= input(21);
output(0, 71) <= input(22);
output(0, 72) <= input(23);
output(0, 73) <= input(24);
output(0, 74) <= input(25);
output(0, 75) <= input(26);
output(0, 76) <= input(27);
output(0, 77) <= input(28);
output(0, 78) <= input(29);
output(0, 79) <= input(30);
output(0, 80) <= input(33);
output(0, 81) <= input(16);
output(0, 82) <= input(17);
output(0, 83) <= input(18);
output(0, 84) <= input(19);
output(0, 85) <= input(20);
output(0, 86) <= input(21);
output(0, 87) <= input(22);
output(0, 88) <= input(23);
output(0, 89) <= input(24);
output(0, 90) <= input(25);
output(0, 91) <= input(26);
output(0, 92) <= input(27);
output(0, 93) <= input(28);
output(0, 94) <= input(29);
output(0, 95) <= input(30);
output(0, 96) <= input(34);
output(0, 97) <= input(32);
output(0, 98) <= input(0);
output(0, 99) <= input(1);
output(0, 100) <= input(2);
output(0, 101) <= input(3);
output(0, 102) <= input(4);
output(0, 103) <= input(5);
output(0, 104) <= input(6);
output(0, 105) <= input(7);
output(0, 106) <= input(8);
output(0, 107) <= input(9);
output(0, 108) <= input(10);
output(0, 109) <= input(11);
output(0, 110) <= input(12);
output(0, 111) <= input(13);
output(0, 112) <= input(34);
output(0, 113) <= input(32);
output(0, 114) <= input(0);
output(0, 115) <= input(1);
output(0, 116) <= input(2);
output(0, 117) <= input(3);
output(0, 118) <= input(4);
output(0, 119) <= input(5);
output(0, 120) <= input(6);
output(0, 121) <= input(7);
output(0, 122) <= input(8);
output(0, 123) <= input(9);
output(0, 124) <= input(10);
output(0, 125) <= input(11);
output(0, 126) <= input(12);
output(0, 127) <= input(13);
output(0, 128) <= input(35);
output(0, 129) <= input(33);
output(0, 130) <= input(16);
output(0, 131) <= input(17);
output(0, 132) <= input(18);
output(0, 133) <= input(19);
output(0, 134) <= input(20);
output(0, 135) <= input(21);
output(0, 136) <= input(22);
output(0, 137) <= input(23);
output(0, 138) <= input(24);
output(0, 139) <= input(25);
output(0, 140) <= input(26);
output(0, 141) <= input(27);
output(0, 142) <= input(28);
output(0, 143) <= input(29);
output(0, 144) <= input(36);
output(0, 145) <= input(34);
output(0, 146) <= input(32);
output(0, 147) <= input(0);
output(0, 148) <= input(1);
output(0, 149) <= input(2);
output(0, 150) <= input(3);
output(0, 151) <= input(4);
output(0, 152) <= input(5);
output(0, 153) <= input(6);
output(0, 154) <= input(7);
output(0, 155) <= input(8);
output(0, 156) <= input(9);
output(0, 157) <= input(10);
output(0, 158) <= input(11);
output(0, 159) <= input(12);
output(0, 160) <= input(36);
output(0, 161) <= input(34);
output(0, 162) <= input(32);
output(0, 163) <= input(0);
output(0, 164) <= input(1);
output(0, 165) <= input(2);
output(0, 166) <= input(3);
output(0, 167) <= input(4);
output(0, 168) <= input(5);
output(0, 169) <= input(6);
output(0, 170) <= input(7);
output(0, 171) <= input(8);
output(0, 172) <= input(9);
output(0, 173) <= input(10);
output(0, 174) <= input(11);
output(0, 175) <= input(12);
output(0, 176) <= input(37);
output(0, 177) <= input(35);
output(0, 178) <= input(33);
output(0, 179) <= input(16);
output(0, 180) <= input(17);
output(0, 181) <= input(18);
output(0, 182) <= input(19);
output(0, 183) <= input(20);
output(0, 184) <= input(21);
output(0, 185) <= input(22);
output(0, 186) <= input(23);
output(0, 187) <= input(24);
output(0, 188) <= input(25);
output(0, 189) <= input(26);
output(0, 190) <= input(27);
output(0, 191) <= input(28);
output(0, 192) <= input(38);
output(0, 193) <= input(36);
output(0, 194) <= input(34);
output(0, 195) <= input(32);
output(0, 196) <= input(0);
output(0, 197) <= input(1);
output(0, 198) <= input(2);
output(0, 199) <= input(3);
output(0, 200) <= input(4);
output(0, 201) <= input(5);
output(0, 202) <= input(6);
output(0, 203) <= input(7);
output(0, 204) <= input(8);
output(0, 205) <= input(9);
output(0, 206) <= input(10);
output(0, 207) <= input(11);
output(0, 208) <= input(38);
output(0, 209) <= input(36);
output(0, 210) <= input(34);
output(0, 211) <= input(32);
output(0, 212) <= input(0);
output(0, 213) <= input(1);
output(0, 214) <= input(2);
output(0, 215) <= input(3);
output(0, 216) <= input(4);
output(0, 217) <= input(5);
output(0, 218) <= input(6);
output(0, 219) <= input(7);
output(0, 220) <= input(8);
output(0, 221) <= input(9);
output(0, 222) <= input(10);
output(0, 223) <= input(11);
output(0, 224) <= input(39);
output(0, 225) <= input(37);
output(0, 226) <= input(35);
output(0, 227) <= input(33);
output(0, 228) <= input(16);
output(0, 229) <= input(17);
output(0, 230) <= input(18);
output(0, 231) <= input(19);
output(0, 232) <= input(20);
output(0, 233) <= input(21);
output(0, 234) <= input(22);
output(0, 235) <= input(23);
output(0, 236) <= input(24);
output(0, 237) <= input(25);
output(0, 238) <= input(26);
output(0, 239) <= input(27);
output(0, 240) <= input(39);
output(0, 241) <= input(37);
output(0, 242) <= input(35);
output(0, 243) <= input(33);
output(0, 244) <= input(16);
output(0, 245) <= input(17);
output(0, 246) <= input(18);
output(0, 247) <= input(19);
output(0, 248) <= input(20);
output(0, 249) <= input(21);
output(0, 250) <= input(22);
output(0, 251) <= input(23);
output(0, 252) <= input(24);
output(0, 253) <= input(25);
output(0, 254) <= input(26);
output(0, 255) <= input(27);
output(1, 0) <= input(0);
output(1, 1) <= input(1);
output(1, 2) <= input(2);
output(1, 3) <= input(3);
output(1, 4) <= input(4);
output(1, 5) <= input(5);
output(1, 6) <= input(6);
output(1, 7) <= input(7);
output(1, 8) <= input(8);
output(1, 9) <= input(9);
output(1, 10) <= input(10);
output(1, 11) <= input(11);
output(1, 12) <= input(12);
output(1, 13) <= input(13);
output(1, 14) <= input(14);
output(1, 15) <= input(15);
output(1, 16) <= input(16);
output(1, 17) <= input(17);
output(1, 18) <= input(18);
output(1, 19) <= input(19);
output(1, 20) <= input(20);
output(1, 21) <= input(21);
output(1, 22) <= input(22);
output(1, 23) <= input(23);
output(1, 24) <= input(24);
output(1, 25) <= input(25);
output(1, 26) <= input(26);
output(1, 27) <= input(27);
output(1, 28) <= input(28);
output(1, 29) <= input(29);
output(1, 30) <= input(30);
output(1, 31) <= input(31);
output(1, 32) <= input(32);
output(1, 33) <= input(0);
output(1, 34) <= input(1);
output(1, 35) <= input(2);
output(1, 36) <= input(3);
output(1, 37) <= input(4);
output(1, 38) <= input(5);
output(1, 39) <= input(6);
output(1, 40) <= input(7);
output(1, 41) <= input(8);
output(1, 42) <= input(9);
output(1, 43) <= input(10);
output(1, 44) <= input(11);
output(1, 45) <= input(12);
output(1, 46) <= input(13);
output(1, 47) <= input(14);
output(1, 48) <= input(32);
output(1, 49) <= input(0);
output(1, 50) <= input(1);
output(1, 51) <= input(2);
output(1, 52) <= input(3);
output(1, 53) <= input(4);
output(1, 54) <= input(5);
output(1, 55) <= input(6);
output(1, 56) <= input(7);
output(1, 57) <= input(8);
output(1, 58) <= input(9);
output(1, 59) <= input(10);
output(1, 60) <= input(11);
output(1, 61) <= input(12);
output(1, 62) <= input(13);
output(1, 63) <= input(14);
output(1, 64) <= input(33);
output(1, 65) <= input(16);
output(1, 66) <= input(17);
output(1, 67) <= input(18);
output(1, 68) <= input(19);
output(1, 69) <= input(20);
output(1, 70) <= input(21);
output(1, 71) <= input(22);
output(1, 72) <= input(23);
output(1, 73) <= input(24);
output(1, 74) <= input(25);
output(1, 75) <= input(26);
output(1, 76) <= input(27);
output(1, 77) <= input(28);
output(1, 78) <= input(29);
output(1, 79) <= input(30);
output(1, 80) <= input(34);
output(1, 81) <= input(32);
output(1, 82) <= input(0);
output(1, 83) <= input(1);
output(1, 84) <= input(2);
output(1, 85) <= input(3);
output(1, 86) <= input(4);
output(1, 87) <= input(5);
output(1, 88) <= input(6);
output(1, 89) <= input(7);
output(1, 90) <= input(8);
output(1, 91) <= input(9);
output(1, 92) <= input(10);
output(1, 93) <= input(11);
output(1, 94) <= input(12);
output(1, 95) <= input(13);
output(1, 96) <= input(35);
output(1, 97) <= input(33);
output(1, 98) <= input(16);
output(1, 99) <= input(17);
output(1, 100) <= input(18);
output(1, 101) <= input(19);
output(1, 102) <= input(20);
output(1, 103) <= input(21);
output(1, 104) <= input(22);
output(1, 105) <= input(23);
output(1, 106) <= input(24);
output(1, 107) <= input(25);
output(1, 108) <= input(26);
output(1, 109) <= input(27);
output(1, 110) <= input(28);
output(1, 111) <= input(29);
output(1, 112) <= input(35);
output(1, 113) <= input(33);
output(1, 114) <= input(16);
output(1, 115) <= input(17);
output(1, 116) <= input(18);
output(1, 117) <= input(19);
output(1, 118) <= input(20);
output(1, 119) <= input(21);
output(1, 120) <= input(22);
output(1, 121) <= input(23);
output(1, 122) <= input(24);
output(1, 123) <= input(25);
output(1, 124) <= input(26);
output(1, 125) <= input(27);
output(1, 126) <= input(28);
output(1, 127) <= input(29);
output(1, 128) <= input(36);
output(1, 129) <= input(34);
output(1, 130) <= input(32);
output(1, 131) <= input(0);
output(1, 132) <= input(1);
output(1, 133) <= input(2);
output(1, 134) <= input(3);
output(1, 135) <= input(4);
output(1, 136) <= input(5);
output(1, 137) <= input(6);
output(1, 138) <= input(7);
output(1, 139) <= input(8);
output(1, 140) <= input(9);
output(1, 141) <= input(10);
output(1, 142) <= input(11);
output(1, 143) <= input(12);
output(1, 144) <= input(37);
output(1, 145) <= input(35);
output(1, 146) <= input(33);
output(1, 147) <= input(16);
output(1, 148) <= input(17);
output(1, 149) <= input(18);
output(1, 150) <= input(19);
output(1, 151) <= input(20);
output(1, 152) <= input(21);
output(1, 153) <= input(22);
output(1, 154) <= input(23);
output(1, 155) <= input(24);
output(1, 156) <= input(25);
output(1, 157) <= input(26);
output(1, 158) <= input(27);
output(1, 159) <= input(28);
output(1, 160) <= input(38);
output(1, 161) <= input(36);
output(1, 162) <= input(34);
output(1, 163) <= input(32);
output(1, 164) <= input(0);
output(1, 165) <= input(1);
output(1, 166) <= input(2);
output(1, 167) <= input(3);
output(1, 168) <= input(4);
output(1, 169) <= input(5);
output(1, 170) <= input(6);
output(1, 171) <= input(7);
output(1, 172) <= input(8);
output(1, 173) <= input(9);
output(1, 174) <= input(10);
output(1, 175) <= input(11);
output(1, 176) <= input(38);
output(1, 177) <= input(36);
output(1, 178) <= input(34);
output(1, 179) <= input(32);
output(1, 180) <= input(0);
output(1, 181) <= input(1);
output(1, 182) <= input(2);
output(1, 183) <= input(3);
output(1, 184) <= input(4);
output(1, 185) <= input(5);
output(1, 186) <= input(6);
output(1, 187) <= input(7);
output(1, 188) <= input(8);
output(1, 189) <= input(9);
output(1, 190) <= input(10);
output(1, 191) <= input(11);
output(1, 192) <= input(39);
output(1, 193) <= input(37);
output(1, 194) <= input(35);
output(1, 195) <= input(33);
output(1, 196) <= input(16);
output(1, 197) <= input(17);
output(1, 198) <= input(18);
output(1, 199) <= input(19);
output(1, 200) <= input(20);
output(1, 201) <= input(21);
output(1, 202) <= input(22);
output(1, 203) <= input(23);
output(1, 204) <= input(24);
output(1, 205) <= input(25);
output(1, 206) <= input(26);
output(1, 207) <= input(27);
output(1, 208) <= input(40);
output(1, 209) <= input(38);
output(1, 210) <= input(36);
output(1, 211) <= input(34);
output(1, 212) <= input(32);
output(1, 213) <= input(0);
output(1, 214) <= input(1);
output(1, 215) <= input(2);
output(1, 216) <= input(3);
output(1, 217) <= input(4);
output(1, 218) <= input(5);
output(1, 219) <= input(6);
output(1, 220) <= input(7);
output(1, 221) <= input(8);
output(1, 222) <= input(9);
output(1, 223) <= input(10);
output(1, 224) <= input(41);
output(1, 225) <= input(39);
output(1, 226) <= input(37);
output(1, 227) <= input(35);
output(1, 228) <= input(33);
output(1, 229) <= input(16);
output(1, 230) <= input(17);
output(1, 231) <= input(18);
output(1, 232) <= input(19);
output(1, 233) <= input(20);
output(1, 234) <= input(21);
output(1, 235) <= input(22);
output(1, 236) <= input(23);
output(1, 237) <= input(24);
output(1, 238) <= input(25);
output(1, 239) <= input(26);
output(1, 240) <= input(41);
output(1, 241) <= input(39);
output(1, 242) <= input(37);
output(1, 243) <= input(35);
output(1, 244) <= input(33);
output(1, 245) <= input(16);
output(1, 246) <= input(17);
output(1, 247) <= input(18);
output(1, 248) <= input(19);
output(1, 249) <= input(20);
output(1, 250) <= input(21);
output(1, 251) <= input(22);
output(1, 252) <= input(23);
output(1, 253) <= input(24);
output(1, 254) <= input(25);
output(1, 255) <= input(26);
output(2, 0) <= input(0);
output(2, 1) <= input(1);
output(2, 2) <= input(2);
output(2, 3) <= input(3);
output(2, 4) <= input(4);
output(2, 5) <= input(5);
output(2, 6) <= input(6);
output(2, 7) <= input(7);
output(2, 8) <= input(8);
output(2, 9) <= input(9);
output(2, 10) <= input(10);
output(2, 11) <= input(11);
output(2, 12) <= input(12);
output(2, 13) <= input(13);
output(2, 14) <= input(14);
output(2, 15) <= input(15);
output(2, 16) <= input(16);
output(2, 17) <= input(17);
output(2, 18) <= input(18);
output(2, 19) <= input(19);
output(2, 20) <= input(20);
output(2, 21) <= input(21);
output(2, 22) <= input(22);
output(2, 23) <= input(23);
output(2, 24) <= input(24);
output(2, 25) <= input(25);
output(2, 26) <= input(26);
output(2, 27) <= input(27);
output(2, 28) <= input(28);
output(2, 29) <= input(29);
output(2, 30) <= input(30);
output(2, 31) <= input(31);
output(2, 32) <= input(32);
output(2, 33) <= input(0);
output(2, 34) <= input(1);
output(2, 35) <= input(2);
output(2, 36) <= input(3);
output(2, 37) <= input(4);
output(2, 38) <= input(5);
output(2, 39) <= input(6);
output(2, 40) <= input(7);
output(2, 41) <= input(8);
output(2, 42) <= input(9);
output(2, 43) <= input(10);
output(2, 44) <= input(11);
output(2, 45) <= input(12);
output(2, 46) <= input(13);
output(2, 47) <= input(14);
output(2, 48) <= input(33);
output(2, 49) <= input(16);
output(2, 50) <= input(17);
output(2, 51) <= input(18);
output(2, 52) <= input(19);
output(2, 53) <= input(20);
output(2, 54) <= input(21);
output(2, 55) <= input(22);
output(2, 56) <= input(23);
output(2, 57) <= input(24);
output(2, 58) <= input(25);
output(2, 59) <= input(26);
output(2, 60) <= input(27);
output(2, 61) <= input(28);
output(2, 62) <= input(29);
output(2, 63) <= input(30);
output(2, 64) <= input(34);
output(2, 65) <= input(32);
output(2, 66) <= input(0);
output(2, 67) <= input(1);
output(2, 68) <= input(2);
output(2, 69) <= input(3);
output(2, 70) <= input(4);
output(2, 71) <= input(5);
output(2, 72) <= input(6);
output(2, 73) <= input(7);
output(2, 74) <= input(8);
output(2, 75) <= input(9);
output(2, 76) <= input(10);
output(2, 77) <= input(11);
output(2, 78) <= input(12);
output(2, 79) <= input(13);
output(2, 80) <= input(35);
output(2, 81) <= input(33);
output(2, 82) <= input(16);
output(2, 83) <= input(17);
output(2, 84) <= input(18);
output(2, 85) <= input(19);
output(2, 86) <= input(20);
output(2, 87) <= input(21);
output(2, 88) <= input(22);
output(2, 89) <= input(23);
output(2, 90) <= input(24);
output(2, 91) <= input(25);
output(2, 92) <= input(26);
output(2, 93) <= input(27);
output(2, 94) <= input(28);
output(2, 95) <= input(29);
output(2, 96) <= input(36);
output(2, 97) <= input(34);
output(2, 98) <= input(32);
output(2, 99) <= input(0);
output(2, 100) <= input(1);
output(2, 101) <= input(2);
output(2, 102) <= input(3);
output(2, 103) <= input(4);
output(2, 104) <= input(5);
output(2, 105) <= input(6);
output(2, 106) <= input(7);
output(2, 107) <= input(8);
output(2, 108) <= input(9);
output(2, 109) <= input(10);
output(2, 110) <= input(11);
output(2, 111) <= input(12);
output(2, 112) <= input(36);
output(2, 113) <= input(34);
output(2, 114) <= input(32);
output(2, 115) <= input(0);
output(2, 116) <= input(1);
output(2, 117) <= input(2);
output(2, 118) <= input(3);
output(2, 119) <= input(4);
output(2, 120) <= input(5);
output(2, 121) <= input(6);
output(2, 122) <= input(7);
output(2, 123) <= input(8);
output(2, 124) <= input(9);
output(2, 125) <= input(10);
output(2, 126) <= input(11);
output(2, 127) <= input(12);
output(2, 128) <= input(37);
output(2, 129) <= input(35);
output(2, 130) <= input(33);
output(2, 131) <= input(16);
output(2, 132) <= input(17);
output(2, 133) <= input(18);
output(2, 134) <= input(19);
output(2, 135) <= input(20);
output(2, 136) <= input(21);
output(2, 137) <= input(22);
output(2, 138) <= input(23);
output(2, 139) <= input(24);
output(2, 140) <= input(25);
output(2, 141) <= input(26);
output(2, 142) <= input(27);
output(2, 143) <= input(28);
output(2, 144) <= input(38);
output(2, 145) <= input(36);
output(2, 146) <= input(34);
output(2, 147) <= input(32);
output(2, 148) <= input(0);
output(2, 149) <= input(1);
output(2, 150) <= input(2);
output(2, 151) <= input(3);
output(2, 152) <= input(4);
output(2, 153) <= input(5);
output(2, 154) <= input(6);
output(2, 155) <= input(7);
output(2, 156) <= input(8);
output(2, 157) <= input(9);
output(2, 158) <= input(10);
output(2, 159) <= input(11);
output(2, 160) <= input(39);
output(2, 161) <= input(37);
output(2, 162) <= input(35);
output(2, 163) <= input(33);
output(2, 164) <= input(16);
output(2, 165) <= input(17);
output(2, 166) <= input(18);
output(2, 167) <= input(19);
output(2, 168) <= input(20);
output(2, 169) <= input(21);
output(2, 170) <= input(22);
output(2, 171) <= input(23);
output(2, 172) <= input(24);
output(2, 173) <= input(25);
output(2, 174) <= input(26);
output(2, 175) <= input(27);
output(2, 176) <= input(40);
output(2, 177) <= input(38);
output(2, 178) <= input(36);
output(2, 179) <= input(34);
output(2, 180) <= input(32);
output(2, 181) <= input(0);
output(2, 182) <= input(1);
output(2, 183) <= input(2);
output(2, 184) <= input(3);
output(2, 185) <= input(4);
output(2, 186) <= input(5);
output(2, 187) <= input(6);
output(2, 188) <= input(7);
output(2, 189) <= input(8);
output(2, 190) <= input(9);
output(2, 191) <= input(10);
output(2, 192) <= input(41);
output(2, 193) <= input(39);
output(2, 194) <= input(37);
output(2, 195) <= input(35);
output(2, 196) <= input(33);
output(2, 197) <= input(16);
output(2, 198) <= input(17);
output(2, 199) <= input(18);
output(2, 200) <= input(19);
output(2, 201) <= input(20);
output(2, 202) <= input(21);
output(2, 203) <= input(22);
output(2, 204) <= input(23);
output(2, 205) <= input(24);
output(2, 206) <= input(25);
output(2, 207) <= input(26);
output(2, 208) <= input(42);
output(2, 209) <= input(40);
output(2, 210) <= input(38);
output(2, 211) <= input(36);
output(2, 212) <= input(34);
output(2, 213) <= input(32);
output(2, 214) <= input(0);
output(2, 215) <= input(1);
output(2, 216) <= input(2);
output(2, 217) <= input(3);
output(2, 218) <= input(4);
output(2, 219) <= input(5);
output(2, 220) <= input(6);
output(2, 221) <= input(7);
output(2, 222) <= input(8);
output(2, 223) <= input(9);
output(2, 224) <= input(43);
output(2, 225) <= input(41);
output(2, 226) <= input(39);
output(2, 227) <= input(37);
output(2, 228) <= input(35);
output(2, 229) <= input(33);
output(2, 230) <= input(16);
output(2, 231) <= input(17);
output(2, 232) <= input(18);
output(2, 233) <= input(19);
output(2, 234) <= input(20);
output(2, 235) <= input(21);
output(2, 236) <= input(22);
output(2, 237) <= input(23);
output(2, 238) <= input(24);
output(2, 239) <= input(25);
output(2, 240) <= input(43);
output(2, 241) <= input(41);
output(2, 242) <= input(39);
output(2, 243) <= input(37);
output(2, 244) <= input(35);
output(2, 245) <= input(33);
output(2, 246) <= input(16);
output(2, 247) <= input(17);
output(2, 248) <= input(18);
output(2, 249) <= input(19);
output(2, 250) <= input(20);
output(2, 251) <= input(21);
output(2, 252) <= input(22);
output(2, 253) <= input(23);
output(2, 254) <= input(24);
output(2, 255) <= input(25);
when "0101" =>
output(0, 0) <= input(0);
output(0, 1) <= input(1);
output(0, 2) <= input(2);
output(0, 3) <= input(3);
output(0, 4) <= input(4);
output(0, 5) <= input(5);
output(0, 6) <= input(6);
output(0, 7) <= input(7);
output(0, 8) <= input(8);
output(0, 9) <= input(9);
output(0, 10) <= input(10);
output(0, 11) <= input(11);
output(0, 12) <= input(12);
output(0, 13) <= input(13);
output(0, 14) <= input(14);
output(0, 15) <= input(15);
output(0, 16) <= input(16);
output(0, 17) <= input(17);
output(0, 18) <= input(18);
output(0, 19) <= input(19);
output(0, 20) <= input(20);
output(0, 21) <= input(21);
output(0, 22) <= input(22);
output(0, 23) <= input(23);
output(0, 24) <= input(24);
output(0, 25) <= input(25);
output(0, 26) <= input(26);
output(0, 27) <= input(27);
output(0, 28) <= input(28);
output(0, 29) <= input(29);
output(0, 30) <= input(30);
output(0, 31) <= input(31);
output(0, 32) <= input(32);
output(0, 33) <= input(0);
output(0, 34) <= input(1);
output(0, 35) <= input(2);
output(0, 36) <= input(3);
output(0, 37) <= input(4);
output(0, 38) <= input(5);
output(0, 39) <= input(6);
output(0, 40) <= input(7);
output(0, 41) <= input(8);
output(0, 42) <= input(9);
output(0, 43) <= input(10);
output(0, 44) <= input(11);
output(0, 45) <= input(12);
output(0, 46) <= input(13);
output(0, 47) <= input(14);
output(0, 48) <= input(33);
output(0, 49) <= input(16);
output(0, 50) <= input(17);
output(0, 51) <= input(18);
output(0, 52) <= input(19);
output(0, 53) <= input(20);
output(0, 54) <= input(21);
output(0, 55) <= input(22);
output(0, 56) <= input(23);
output(0, 57) <= input(24);
output(0, 58) <= input(25);
output(0, 59) <= input(26);
output(0, 60) <= input(27);
output(0, 61) <= input(28);
output(0, 62) <= input(29);
output(0, 63) <= input(30);
output(0, 64) <= input(34);
output(0, 65) <= input(32);
output(0, 66) <= input(0);
output(0, 67) <= input(1);
output(0, 68) <= input(2);
output(0, 69) <= input(3);
output(0, 70) <= input(4);
output(0, 71) <= input(5);
output(0, 72) <= input(6);
output(0, 73) <= input(7);
output(0, 74) <= input(8);
output(0, 75) <= input(9);
output(0, 76) <= input(10);
output(0, 77) <= input(11);
output(0, 78) <= input(12);
output(0, 79) <= input(13);
output(0, 80) <= input(35);
output(0, 81) <= input(33);
output(0, 82) <= input(16);
output(0, 83) <= input(17);
output(0, 84) <= input(18);
output(0, 85) <= input(19);
output(0, 86) <= input(20);
output(0, 87) <= input(21);
output(0, 88) <= input(22);
output(0, 89) <= input(23);
output(0, 90) <= input(24);
output(0, 91) <= input(25);
output(0, 92) <= input(26);
output(0, 93) <= input(27);
output(0, 94) <= input(28);
output(0, 95) <= input(29);
output(0, 96) <= input(36);
output(0, 97) <= input(34);
output(0, 98) <= input(32);
output(0, 99) <= input(0);
output(0, 100) <= input(1);
output(0, 101) <= input(2);
output(0, 102) <= input(3);
output(0, 103) <= input(4);
output(0, 104) <= input(5);
output(0, 105) <= input(6);
output(0, 106) <= input(7);
output(0, 107) <= input(8);
output(0, 108) <= input(9);
output(0, 109) <= input(10);
output(0, 110) <= input(11);
output(0, 111) <= input(12);
output(0, 112) <= input(37);
output(0, 113) <= input(35);
output(0, 114) <= input(33);
output(0, 115) <= input(16);
output(0, 116) <= input(17);
output(0, 117) <= input(18);
output(0, 118) <= input(19);
output(0, 119) <= input(20);
output(0, 120) <= input(21);
output(0, 121) <= input(22);
output(0, 122) <= input(23);
output(0, 123) <= input(24);
output(0, 124) <= input(25);
output(0, 125) <= input(26);
output(0, 126) <= input(27);
output(0, 127) <= input(28);
output(0, 128) <= input(38);
output(0, 129) <= input(36);
output(0, 130) <= input(34);
output(0, 131) <= input(32);
output(0, 132) <= input(0);
output(0, 133) <= input(1);
output(0, 134) <= input(2);
output(0, 135) <= input(3);
output(0, 136) <= input(4);
output(0, 137) <= input(5);
output(0, 138) <= input(6);
output(0, 139) <= input(7);
output(0, 140) <= input(8);
output(0, 141) <= input(9);
output(0, 142) <= input(10);
output(0, 143) <= input(11);
output(0, 144) <= input(39);
output(0, 145) <= input(37);
output(0, 146) <= input(35);
output(0, 147) <= input(33);
output(0, 148) <= input(16);
output(0, 149) <= input(17);
output(0, 150) <= input(18);
output(0, 151) <= input(19);
output(0, 152) <= input(20);
output(0, 153) <= input(21);
output(0, 154) <= input(22);
output(0, 155) <= input(23);
output(0, 156) <= input(24);
output(0, 157) <= input(25);
output(0, 158) <= input(26);
output(0, 159) <= input(27);
output(0, 160) <= input(40);
output(0, 161) <= input(38);
output(0, 162) <= input(36);
output(0, 163) <= input(34);
output(0, 164) <= input(32);
output(0, 165) <= input(0);
output(0, 166) <= input(1);
output(0, 167) <= input(2);
output(0, 168) <= input(3);
output(0, 169) <= input(4);
output(0, 170) <= input(5);
output(0, 171) <= input(6);
output(0, 172) <= input(7);
output(0, 173) <= input(8);
output(0, 174) <= input(9);
output(0, 175) <= input(10);
output(0, 176) <= input(41);
output(0, 177) <= input(39);
output(0, 178) <= input(37);
output(0, 179) <= input(35);
output(0, 180) <= input(33);
output(0, 181) <= input(16);
output(0, 182) <= input(17);
output(0, 183) <= input(18);
output(0, 184) <= input(19);
output(0, 185) <= input(20);
output(0, 186) <= input(21);
output(0, 187) <= input(22);
output(0, 188) <= input(23);
output(0, 189) <= input(24);
output(0, 190) <= input(25);
output(0, 191) <= input(26);
output(0, 192) <= input(42);
output(0, 193) <= input(40);
output(0, 194) <= input(38);
output(0, 195) <= input(36);
output(0, 196) <= input(34);
output(0, 197) <= input(32);
output(0, 198) <= input(0);
output(0, 199) <= input(1);
output(0, 200) <= input(2);
output(0, 201) <= input(3);
output(0, 202) <= input(4);
output(0, 203) <= input(5);
output(0, 204) <= input(6);
output(0, 205) <= input(7);
output(0, 206) <= input(8);
output(0, 207) <= input(9);
output(0, 208) <= input(43);
output(0, 209) <= input(41);
output(0, 210) <= input(39);
output(0, 211) <= input(37);
output(0, 212) <= input(35);
output(0, 213) <= input(33);
output(0, 214) <= input(16);
output(0, 215) <= input(17);
output(0, 216) <= input(18);
output(0, 217) <= input(19);
output(0, 218) <= input(20);
output(0, 219) <= input(21);
output(0, 220) <= input(22);
output(0, 221) <= input(23);
output(0, 222) <= input(24);
output(0, 223) <= input(25);
output(0, 224) <= input(44);
output(0, 225) <= input(42);
output(0, 226) <= input(40);
output(0, 227) <= input(38);
output(0, 228) <= input(36);
output(0, 229) <= input(34);
output(0, 230) <= input(32);
output(0, 231) <= input(0);
output(0, 232) <= input(1);
output(0, 233) <= input(2);
output(0, 234) <= input(3);
output(0, 235) <= input(4);
output(0, 236) <= input(5);
output(0, 237) <= input(6);
output(0, 238) <= input(7);
output(0, 239) <= input(8);
output(0, 240) <= input(45);
output(0, 241) <= input(43);
output(0, 242) <= input(41);
output(0, 243) <= input(39);
output(0, 244) <= input(37);
output(0, 245) <= input(35);
output(0, 246) <= input(33);
output(0, 247) <= input(16);
output(0, 248) <= input(17);
output(0, 249) <= input(18);
output(0, 250) <= input(19);
output(0, 251) <= input(20);
output(0, 252) <= input(21);
output(0, 253) <= input(22);
output(0, 254) <= input(23);
output(0, 255) <= input(24);
output(1, 0) <= input(16);
output(1, 1) <= input(17);
output(1, 2) <= input(18);
output(1, 3) <= input(19);
output(1, 4) <= input(20);
output(1, 5) <= input(21);
output(1, 6) <= input(22);
output(1, 7) <= input(23);
output(1, 8) <= input(24);
output(1, 9) <= input(25);
output(1, 10) <= input(26);
output(1, 11) <= input(27);
output(1, 12) <= input(28);
output(1, 13) <= input(29);
output(1, 14) <= input(30);
output(1, 15) <= input(31);
output(1, 16) <= input(32);
output(1, 17) <= input(0);
output(1, 18) <= input(1);
output(1, 19) <= input(2);
output(1, 20) <= input(3);
output(1, 21) <= input(4);
output(1, 22) <= input(5);
output(1, 23) <= input(6);
output(1, 24) <= input(7);
output(1, 25) <= input(8);
output(1, 26) <= input(9);
output(1, 27) <= input(10);
output(1, 28) <= input(11);
output(1, 29) <= input(12);
output(1, 30) <= input(13);
output(1, 31) <= input(14);
output(1, 32) <= input(33);
output(1, 33) <= input(16);
output(1, 34) <= input(17);
output(1, 35) <= input(18);
output(1, 36) <= input(19);
output(1, 37) <= input(20);
output(1, 38) <= input(21);
output(1, 39) <= input(22);
output(1, 40) <= input(23);
output(1, 41) <= input(24);
output(1, 42) <= input(25);
output(1, 43) <= input(26);
output(1, 44) <= input(27);
output(1, 45) <= input(28);
output(1, 46) <= input(29);
output(1, 47) <= input(30);
output(1, 48) <= input(34);
output(1, 49) <= input(32);
output(1, 50) <= input(0);
output(1, 51) <= input(1);
output(1, 52) <= input(2);
output(1, 53) <= input(3);
output(1, 54) <= input(4);
output(1, 55) <= input(5);
output(1, 56) <= input(6);
output(1, 57) <= input(7);
output(1, 58) <= input(8);
output(1, 59) <= input(9);
output(1, 60) <= input(10);
output(1, 61) <= input(11);
output(1, 62) <= input(12);
output(1, 63) <= input(13);
output(1, 64) <= input(35);
output(1, 65) <= input(33);
output(1, 66) <= input(16);
output(1, 67) <= input(17);
output(1, 68) <= input(18);
output(1, 69) <= input(19);
output(1, 70) <= input(20);
output(1, 71) <= input(21);
output(1, 72) <= input(22);
output(1, 73) <= input(23);
output(1, 74) <= input(24);
output(1, 75) <= input(25);
output(1, 76) <= input(26);
output(1, 77) <= input(27);
output(1, 78) <= input(28);
output(1, 79) <= input(29);
output(1, 80) <= input(36);
output(1, 81) <= input(34);
output(1, 82) <= input(32);
output(1, 83) <= input(0);
output(1, 84) <= input(1);
output(1, 85) <= input(2);
output(1, 86) <= input(3);
output(1, 87) <= input(4);
output(1, 88) <= input(5);
output(1, 89) <= input(6);
output(1, 90) <= input(7);
output(1, 91) <= input(8);
output(1, 92) <= input(9);
output(1, 93) <= input(10);
output(1, 94) <= input(11);
output(1, 95) <= input(12);
output(1, 96) <= input(37);
output(1, 97) <= input(35);
output(1, 98) <= input(33);
output(1, 99) <= input(16);
output(1, 100) <= input(17);
output(1, 101) <= input(18);
output(1, 102) <= input(19);
output(1, 103) <= input(20);
output(1, 104) <= input(21);
output(1, 105) <= input(22);
output(1, 106) <= input(23);
output(1, 107) <= input(24);
output(1, 108) <= input(25);
output(1, 109) <= input(26);
output(1, 110) <= input(27);
output(1, 111) <= input(28);
output(1, 112) <= input(38);
output(1, 113) <= input(36);
output(1, 114) <= input(34);
output(1, 115) <= input(32);
output(1, 116) <= input(0);
output(1, 117) <= input(1);
output(1, 118) <= input(2);
output(1, 119) <= input(3);
output(1, 120) <= input(4);
output(1, 121) <= input(5);
output(1, 122) <= input(6);
output(1, 123) <= input(7);
output(1, 124) <= input(8);
output(1, 125) <= input(9);
output(1, 126) <= input(10);
output(1, 127) <= input(11);
output(1, 128) <= input(40);
output(1, 129) <= input(38);
output(1, 130) <= input(36);
output(1, 131) <= input(34);
output(1, 132) <= input(32);
output(1, 133) <= input(0);
output(1, 134) <= input(1);
output(1, 135) <= input(2);
output(1, 136) <= input(3);
output(1, 137) <= input(4);
output(1, 138) <= input(5);
output(1, 139) <= input(6);
output(1, 140) <= input(7);
output(1, 141) <= input(8);
output(1, 142) <= input(9);
output(1, 143) <= input(10);
output(1, 144) <= input(41);
output(1, 145) <= input(39);
output(1, 146) <= input(37);
output(1, 147) <= input(35);
output(1, 148) <= input(33);
output(1, 149) <= input(16);
output(1, 150) <= input(17);
output(1, 151) <= input(18);
output(1, 152) <= input(19);
output(1, 153) <= input(20);
output(1, 154) <= input(21);
output(1, 155) <= input(22);
output(1, 156) <= input(23);
output(1, 157) <= input(24);
output(1, 158) <= input(25);
output(1, 159) <= input(26);
output(1, 160) <= input(42);
output(1, 161) <= input(40);
output(1, 162) <= input(38);
output(1, 163) <= input(36);
output(1, 164) <= input(34);
output(1, 165) <= input(32);
output(1, 166) <= input(0);
output(1, 167) <= input(1);
output(1, 168) <= input(2);
output(1, 169) <= input(3);
output(1, 170) <= input(4);
output(1, 171) <= input(5);
output(1, 172) <= input(6);
output(1, 173) <= input(7);
output(1, 174) <= input(8);
output(1, 175) <= input(9);
output(1, 176) <= input(43);
output(1, 177) <= input(41);
output(1, 178) <= input(39);
output(1, 179) <= input(37);
output(1, 180) <= input(35);
output(1, 181) <= input(33);
output(1, 182) <= input(16);
output(1, 183) <= input(17);
output(1, 184) <= input(18);
output(1, 185) <= input(19);
output(1, 186) <= input(20);
output(1, 187) <= input(21);
output(1, 188) <= input(22);
output(1, 189) <= input(23);
output(1, 190) <= input(24);
output(1, 191) <= input(25);
output(1, 192) <= input(44);
output(1, 193) <= input(42);
output(1, 194) <= input(40);
output(1, 195) <= input(38);
output(1, 196) <= input(36);
output(1, 197) <= input(34);
output(1, 198) <= input(32);
output(1, 199) <= input(0);
output(1, 200) <= input(1);
output(1, 201) <= input(2);
output(1, 202) <= input(3);
output(1, 203) <= input(4);
output(1, 204) <= input(5);
output(1, 205) <= input(6);
output(1, 206) <= input(7);
output(1, 207) <= input(8);
output(1, 208) <= input(45);
output(1, 209) <= input(43);
output(1, 210) <= input(41);
output(1, 211) <= input(39);
output(1, 212) <= input(37);
output(1, 213) <= input(35);
output(1, 214) <= input(33);
output(1, 215) <= input(16);
output(1, 216) <= input(17);
output(1, 217) <= input(18);
output(1, 218) <= input(19);
output(1, 219) <= input(20);
output(1, 220) <= input(21);
output(1, 221) <= input(22);
output(1, 222) <= input(23);
output(1, 223) <= input(24);
output(1, 224) <= input(46);
output(1, 225) <= input(44);
output(1, 226) <= input(42);
output(1, 227) <= input(40);
output(1, 228) <= input(38);
output(1, 229) <= input(36);
output(1, 230) <= input(34);
output(1, 231) <= input(32);
output(1, 232) <= input(0);
output(1, 233) <= input(1);
output(1, 234) <= input(2);
output(1, 235) <= input(3);
output(1, 236) <= input(4);
output(1, 237) <= input(5);
output(1, 238) <= input(6);
output(1, 239) <= input(7);
output(1, 240) <= input(47);
output(1, 241) <= input(45);
output(1, 242) <= input(43);
output(1, 243) <= input(41);
output(1, 244) <= input(39);
output(1, 245) <= input(37);
output(1, 246) <= input(35);
output(1, 247) <= input(33);
output(1, 248) <= input(16);
output(1, 249) <= input(17);
output(1, 250) <= input(18);
output(1, 251) <= input(19);
output(1, 252) <= input(20);
output(1, 253) <= input(21);
output(1, 254) <= input(22);
output(1, 255) <= input(23);
when "0110" =>
output(0, 0) <= input(0);
output(0, 1) <= input(1);
output(0, 2) <= input(2);
output(0, 3) <= input(3);
output(0, 4) <= input(4);
output(0, 5) <= input(5);
output(0, 6) <= input(6);
output(0, 7) <= input(7);
output(0, 8) <= input(8);
output(0, 9) <= input(9);
output(0, 10) <= input(10);
output(0, 11) <= input(11);
output(0, 12) <= input(12);
output(0, 13) <= input(13);
output(0, 14) <= input(14);
output(0, 15) <= input(15);
output(0, 16) <= input(16);
output(0, 17) <= input(17);
output(0, 18) <= input(18);
output(0, 19) <= input(19);
output(0, 20) <= input(20);
output(0, 21) <= input(21);
output(0, 22) <= input(22);
output(0, 23) <= input(23);
output(0, 24) <= input(24);
output(0, 25) <= input(25);
output(0, 26) <= input(26);
output(0, 27) <= input(27);
output(0, 28) <= input(28);
output(0, 29) <= input(29);
output(0, 30) <= input(30);
output(0, 31) <= input(31);
output(0, 32) <= input(32);
output(0, 33) <= input(0);
output(0, 34) <= input(1);
output(0, 35) <= input(2);
output(0, 36) <= input(3);
output(0, 37) <= input(4);
output(0, 38) <= input(5);
output(0, 39) <= input(6);
output(0, 40) <= input(7);
output(0, 41) <= input(8);
output(0, 42) <= input(9);
output(0, 43) <= input(10);
output(0, 44) <= input(11);
output(0, 45) <= input(12);
output(0, 46) <= input(13);
output(0, 47) <= input(14);
output(0, 48) <= input(33);
output(0, 49) <= input(16);
output(0, 50) <= input(17);
output(0, 51) <= input(18);
output(0, 52) <= input(19);
output(0, 53) <= input(20);
output(0, 54) <= input(21);
output(0, 55) <= input(22);
output(0, 56) <= input(23);
output(0, 57) <= input(24);
output(0, 58) <= input(25);
output(0, 59) <= input(26);
output(0, 60) <= input(27);
output(0, 61) <= input(28);
output(0, 62) <= input(29);
output(0, 63) <= input(30);
output(0, 64) <= input(34);
output(0, 65) <= input(33);
output(0, 66) <= input(16);
output(0, 67) <= input(17);
output(0, 68) <= input(18);
output(0, 69) <= input(19);
output(0, 70) <= input(20);
output(0, 71) <= input(21);
output(0, 72) <= input(22);
output(0, 73) <= input(23);
output(0, 74) <= input(24);
output(0, 75) <= input(25);
output(0, 76) <= input(26);
output(0, 77) <= input(27);
output(0, 78) <= input(28);
output(0, 79) <= input(29);
output(0, 80) <= input(35);
output(0, 81) <= input(36);
output(0, 82) <= input(32);
output(0, 83) <= input(0);
output(0, 84) <= input(1);
output(0, 85) <= input(2);
output(0, 86) <= input(3);
output(0, 87) <= input(4);
output(0, 88) <= input(5);
output(0, 89) <= input(6);
output(0, 90) <= input(7);
output(0, 91) <= input(8);
output(0, 92) <= input(9);
output(0, 93) <= input(10);
output(0, 94) <= input(11);
output(0, 95) <= input(12);
output(0, 96) <= input(37);
output(0, 97) <= input(34);
output(0, 98) <= input(33);
output(0, 99) <= input(16);
output(0, 100) <= input(17);
output(0, 101) <= input(18);
output(0, 102) <= input(19);
output(0, 103) <= input(20);
output(0, 104) <= input(21);
output(0, 105) <= input(22);
output(0, 106) <= input(23);
output(0, 107) <= input(24);
output(0, 108) <= input(25);
output(0, 109) <= input(26);
output(0, 110) <= input(27);
output(0, 111) <= input(28);
output(0, 112) <= input(38);
output(0, 113) <= input(35);
output(0, 114) <= input(36);
output(0, 115) <= input(32);
output(0, 116) <= input(0);
output(0, 117) <= input(1);
output(0, 118) <= input(2);
output(0, 119) <= input(3);
output(0, 120) <= input(4);
output(0, 121) <= input(5);
output(0, 122) <= input(6);
output(0, 123) <= input(7);
output(0, 124) <= input(8);
output(0, 125) <= input(9);
output(0, 126) <= input(10);
output(0, 127) <= input(11);
output(0, 128) <= input(39);
output(0, 129) <= input(38);
output(0, 130) <= input(35);
output(0, 131) <= input(36);
output(0, 132) <= input(32);
output(0, 133) <= input(0);
output(0, 134) <= input(1);
output(0, 135) <= input(2);
output(0, 136) <= input(3);
output(0, 137) <= input(4);
output(0, 138) <= input(5);
output(0, 139) <= input(6);
output(0, 140) <= input(7);
output(0, 141) <= input(8);
output(0, 142) <= input(9);
output(0, 143) <= input(10);
output(0, 144) <= input(40);
output(0, 145) <= input(41);
output(0, 146) <= input(37);
output(0, 147) <= input(34);
output(0, 148) <= input(33);
output(0, 149) <= input(16);
output(0, 150) <= input(17);
output(0, 151) <= input(18);
output(0, 152) <= input(19);
output(0, 153) <= input(20);
output(0, 154) <= input(21);
output(0, 155) <= input(22);
output(0, 156) <= input(23);
output(0, 157) <= input(24);
output(0, 158) <= input(25);
output(0, 159) <= input(26);
output(0, 160) <= input(42);
output(0, 161) <= input(39);
output(0, 162) <= input(38);
output(0, 163) <= input(35);
output(0, 164) <= input(36);
output(0, 165) <= input(32);
output(0, 166) <= input(0);
output(0, 167) <= input(1);
output(0, 168) <= input(2);
output(0, 169) <= input(3);
output(0, 170) <= input(4);
output(0, 171) <= input(5);
output(0, 172) <= input(6);
output(0, 173) <= input(7);
output(0, 174) <= input(8);
output(0, 175) <= input(9);
output(0, 176) <= input(43);
output(0, 177) <= input(40);
output(0, 178) <= input(41);
output(0, 179) <= input(37);
output(0, 180) <= input(34);
output(0, 181) <= input(33);
output(0, 182) <= input(16);
output(0, 183) <= input(17);
output(0, 184) <= input(18);
output(0, 185) <= input(19);
output(0, 186) <= input(20);
output(0, 187) <= input(21);
output(0, 188) <= input(22);
output(0, 189) <= input(23);
output(0, 190) <= input(24);
output(0, 191) <= input(25);
output(0, 192) <= input(44);
output(0, 193) <= input(43);
output(0, 194) <= input(40);
output(0, 195) <= input(41);
output(0, 196) <= input(37);
output(0, 197) <= input(34);
output(0, 198) <= input(33);
output(0, 199) <= input(16);
output(0, 200) <= input(17);
output(0, 201) <= input(18);
output(0, 202) <= input(19);
output(0, 203) <= input(20);
output(0, 204) <= input(21);
output(0, 205) <= input(22);
output(0, 206) <= input(23);
output(0, 207) <= input(24);
output(0, 208) <= input(45);
output(0, 209) <= input(46);
output(0, 210) <= input(42);
output(0, 211) <= input(39);
output(0, 212) <= input(38);
output(0, 213) <= input(35);
output(0, 214) <= input(36);
output(0, 215) <= input(32);
output(0, 216) <= input(0);
output(0, 217) <= input(1);
output(0, 218) <= input(2);
output(0, 219) <= input(3);
output(0, 220) <= input(4);
output(0, 221) <= input(5);
output(0, 222) <= input(6);
output(0, 223) <= input(7);
output(0, 224) <= input(47);
output(0, 225) <= input(44);
output(0, 226) <= input(43);
output(0, 227) <= input(40);
output(0, 228) <= input(41);
output(0, 229) <= input(37);
output(0, 230) <= input(34);
output(0, 231) <= input(33);
output(0, 232) <= input(16);
output(0, 233) <= input(17);
output(0, 234) <= input(18);
output(0, 235) <= input(19);
output(0, 236) <= input(20);
output(0, 237) <= input(21);
output(0, 238) <= input(22);
output(0, 239) <= input(23);
output(0, 240) <= input(48);
output(0, 241) <= input(45);
output(0, 242) <= input(46);
output(0, 243) <= input(42);
output(0, 244) <= input(39);
output(0, 245) <= input(38);
output(0, 246) <= input(35);
output(0, 247) <= input(36);
output(0, 248) <= input(32);
output(0, 249) <= input(0);
output(0, 250) <= input(1);
output(0, 251) <= input(2);
output(0, 252) <= input(3);
output(0, 253) <= input(4);
output(0, 254) <= input(5);
output(0, 255) <= input(6);
output(1, 0) <= input(0);
output(1, 1) <= input(1);
output(1, 2) <= input(2);
output(1, 3) <= input(3);
output(1, 4) <= input(4);
output(1, 5) <= input(5);
output(1, 6) <= input(6);
output(1, 7) <= input(7);
output(1, 8) <= input(8);
output(1, 9) <= input(9);
output(1, 10) <= input(10);
output(1, 11) <= input(11);
output(1, 12) <= input(12);
output(1, 13) <= input(13);
output(1, 14) <= input(14);
output(1, 15) <= input(15);
output(1, 16) <= input(16);
output(1, 17) <= input(17);
output(1, 18) <= input(18);
output(1, 19) <= input(19);
output(1, 20) <= input(20);
output(1, 21) <= input(21);
output(1, 22) <= input(22);
output(1, 23) <= input(23);
output(1, 24) <= input(24);
output(1, 25) <= input(25);
output(1, 26) <= input(26);
output(1, 27) <= input(27);
output(1, 28) <= input(28);
output(1, 29) <= input(29);
output(1, 30) <= input(30);
output(1, 31) <= input(31);
output(1, 32) <= input(33);
output(1, 33) <= input(16);
output(1, 34) <= input(17);
output(1, 35) <= input(18);
output(1, 36) <= input(19);
output(1, 37) <= input(20);
output(1, 38) <= input(21);
output(1, 39) <= input(22);
output(1, 40) <= input(23);
output(1, 41) <= input(24);
output(1, 42) <= input(25);
output(1, 43) <= input(26);
output(1, 44) <= input(27);
output(1, 45) <= input(28);
output(1, 46) <= input(29);
output(1, 47) <= input(30);
output(1, 48) <= input(36);
output(1, 49) <= input(32);
output(1, 50) <= input(0);
output(1, 51) <= input(1);
output(1, 52) <= input(2);
output(1, 53) <= input(3);
output(1, 54) <= input(4);
output(1, 55) <= input(5);
output(1, 56) <= input(6);
output(1, 57) <= input(7);
output(1, 58) <= input(8);
output(1, 59) <= input(9);
output(1, 60) <= input(10);
output(1, 61) <= input(11);
output(1, 62) <= input(12);
output(1, 63) <= input(13);
output(1, 64) <= input(35);
output(1, 65) <= input(36);
output(1, 66) <= input(32);
output(1, 67) <= input(0);
output(1, 68) <= input(1);
output(1, 69) <= input(2);
output(1, 70) <= input(3);
output(1, 71) <= input(4);
output(1, 72) <= input(5);
output(1, 73) <= input(6);
output(1, 74) <= input(7);
output(1, 75) <= input(8);
output(1, 76) <= input(9);
output(1, 77) <= input(10);
output(1, 78) <= input(11);
output(1, 79) <= input(12);
output(1, 80) <= input(37);
output(1, 81) <= input(34);
output(1, 82) <= input(33);
output(1, 83) <= input(16);
output(1, 84) <= input(17);
output(1, 85) <= input(18);
output(1, 86) <= input(19);
output(1, 87) <= input(20);
output(1, 88) <= input(21);
output(1, 89) <= input(22);
output(1, 90) <= input(23);
output(1, 91) <= input(24);
output(1, 92) <= input(25);
output(1, 93) <= input(26);
output(1, 94) <= input(27);
output(1, 95) <= input(28);
output(1, 96) <= input(41);
output(1, 97) <= input(37);
output(1, 98) <= input(34);
output(1, 99) <= input(33);
output(1, 100) <= input(16);
output(1, 101) <= input(17);
output(1, 102) <= input(18);
output(1, 103) <= input(19);
output(1, 104) <= input(20);
output(1, 105) <= input(21);
output(1, 106) <= input(22);
output(1, 107) <= input(23);
output(1, 108) <= input(24);
output(1, 109) <= input(25);
output(1, 110) <= input(26);
output(1, 111) <= input(27);
output(1, 112) <= input(39);
output(1, 113) <= input(38);
output(1, 114) <= input(35);
output(1, 115) <= input(36);
output(1, 116) <= input(32);
output(1, 117) <= input(0);
output(1, 118) <= input(1);
output(1, 119) <= input(2);
output(1, 120) <= input(3);
output(1, 121) <= input(4);
output(1, 122) <= input(5);
output(1, 123) <= input(6);
output(1, 124) <= input(7);
output(1, 125) <= input(8);
output(1, 126) <= input(9);
output(1, 127) <= input(10);
output(1, 128) <= input(40);
output(1, 129) <= input(41);
output(1, 130) <= input(37);
output(1, 131) <= input(34);
output(1, 132) <= input(33);
output(1, 133) <= input(16);
output(1, 134) <= input(17);
output(1, 135) <= input(18);
output(1, 136) <= input(19);
output(1, 137) <= input(20);
output(1, 138) <= input(21);
output(1, 139) <= input(22);
output(1, 140) <= input(23);
output(1, 141) <= input(24);
output(1, 142) <= input(25);
output(1, 143) <= input(26);
output(1, 144) <= input(43);
output(1, 145) <= input(40);
output(1, 146) <= input(41);
output(1, 147) <= input(37);
output(1, 148) <= input(34);
output(1, 149) <= input(33);
output(1, 150) <= input(16);
output(1, 151) <= input(17);
output(1, 152) <= input(18);
output(1, 153) <= input(19);
output(1, 154) <= input(20);
output(1, 155) <= input(21);
output(1, 156) <= input(22);
output(1, 157) <= input(23);
output(1, 158) <= input(24);
output(1, 159) <= input(25);
output(1, 160) <= input(46);
output(1, 161) <= input(42);
output(1, 162) <= input(39);
output(1, 163) <= input(38);
output(1, 164) <= input(35);
output(1, 165) <= input(36);
output(1, 166) <= input(32);
output(1, 167) <= input(0);
output(1, 168) <= input(1);
output(1, 169) <= input(2);
output(1, 170) <= input(3);
output(1, 171) <= input(4);
output(1, 172) <= input(5);
output(1, 173) <= input(6);
output(1, 174) <= input(7);
output(1, 175) <= input(8);
output(1, 176) <= input(45);
output(1, 177) <= input(46);
output(1, 178) <= input(42);
output(1, 179) <= input(39);
output(1, 180) <= input(38);
output(1, 181) <= input(35);
output(1, 182) <= input(36);
output(1, 183) <= input(32);
output(1, 184) <= input(0);
output(1, 185) <= input(1);
output(1, 186) <= input(2);
output(1, 187) <= input(3);
output(1, 188) <= input(4);
output(1, 189) <= input(5);
output(1, 190) <= input(6);
output(1, 191) <= input(7);
output(1, 192) <= input(47);
output(1, 193) <= input(44);
output(1, 194) <= input(43);
output(1, 195) <= input(40);
output(1, 196) <= input(41);
output(1, 197) <= input(37);
output(1, 198) <= input(34);
output(1, 199) <= input(33);
output(1, 200) <= input(16);
output(1, 201) <= input(17);
output(1, 202) <= input(18);
output(1, 203) <= input(19);
output(1, 204) <= input(20);
output(1, 205) <= input(21);
output(1, 206) <= input(22);
output(1, 207) <= input(23);
output(1, 208) <= input(49);
output(1, 209) <= input(47);
output(1, 210) <= input(44);
output(1, 211) <= input(43);
output(1, 212) <= input(40);
output(1, 213) <= input(41);
output(1, 214) <= input(37);
output(1, 215) <= input(34);
output(1, 216) <= input(33);
output(1, 217) <= input(16);
output(1, 218) <= input(17);
output(1, 219) <= input(18);
output(1, 220) <= input(19);
output(1, 221) <= input(20);
output(1, 222) <= input(21);
output(1, 223) <= input(22);
output(1, 224) <= input(50);
output(1, 225) <= input(48);
output(1, 226) <= input(45);
output(1, 227) <= input(46);
output(1, 228) <= input(42);
output(1, 229) <= input(39);
output(1, 230) <= input(38);
output(1, 231) <= input(35);
output(1, 232) <= input(36);
output(1, 233) <= input(32);
output(1, 234) <= input(0);
output(1, 235) <= input(1);
output(1, 236) <= input(2);
output(1, 237) <= input(3);
output(1, 238) <= input(4);
output(1, 239) <= input(5);
output(1, 240) <= input(51);
output(1, 241) <= input(49);
output(1, 242) <= input(47);
output(1, 243) <= input(44);
output(1, 244) <= input(43);
output(1, 245) <= input(40);
output(1, 246) <= input(41);
output(1, 247) <= input(37);
output(1, 248) <= input(34);
output(1, 249) <= input(33);
output(1, 250) <= input(16);
output(1, 251) <= input(17);
output(1, 252) <= input(18);
output(1, 253) <= input(19);
output(1, 254) <= input(20);
output(1, 255) <= input(21);
output(2, 0) <= input(0);
output(2, 1) <= input(1);
output(2, 2) <= input(2);
output(2, 3) <= input(3);
output(2, 4) <= input(4);
output(2, 5) <= input(5);
output(2, 6) <= input(6);
output(2, 7) <= input(7);
output(2, 8) <= input(8);
output(2, 9) <= input(9);
output(2, 10) <= input(10);
output(2, 11) <= input(11);
output(2, 12) <= input(12);
output(2, 13) <= input(13);
output(2, 14) <= input(14);
output(2, 15) <= input(15);
output(2, 16) <= input(32);
output(2, 17) <= input(0);
output(2, 18) <= input(1);
output(2, 19) <= input(2);
output(2, 20) <= input(3);
output(2, 21) <= input(4);
output(2, 22) <= input(5);
output(2, 23) <= input(6);
output(2, 24) <= input(7);
output(2, 25) <= input(8);
output(2, 26) <= input(9);
output(2, 27) <= input(10);
output(2, 28) <= input(11);
output(2, 29) <= input(12);
output(2, 30) <= input(13);
output(2, 31) <= input(14);
output(2, 32) <= input(33);
output(2, 33) <= input(16);
output(2, 34) <= input(17);
output(2, 35) <= input(18);
output(2, 36) <= input(19);
output(2, 37) <= input(20);
output(2, 38) <= input(21);
output(2, 39) <= input(22);
output(2, 40) <= input(23);
output(2, 41) <= input(24);
output(2, 42) <= input(25);
output(2, 43) <= input(26);
output(2, 44) <= input(27);
output(2, 45) <= input(28);
output(2, 46) <= input(29);
output(2, 47) <= input(30);
output(2, 48) <= input(34);
output(2, 49) <= input(33);
output(2, 50) <= input(16);
output(2, 51) <= input(17);
output(2, 52) <= input(18);
output(2, 53) <= input(19);
output(2, 54) <= input(20);
output(2, 55) <= input(21);
output(2, 56) <= input(22);
output(2, 57) <= input(23);
output(2, 58) <= input(24);
output(2, 59) <= input(25);
output(2, 60) <= input(26);
output(2, 61) <= input(27);
output(2, 62) <= input(28);
output(2, 63) <= input(29);
output(2, 64) <= input(37);
output(2, 65) <= input(34);
output(2, 66) <= input(33);
output(2, 67) <= input(16);
output(2, 68) <= input(17);
output(2, 69) <= input(18);
output(2, 70) <= input(19);
output(2, 71) <= input(20);
output(2, 72) <= input(21);
output(2, 73) <= input(22);
output(2, 74) <= input(23);
output(2, 75) <= input(24);
output(2, 76) <= input(25);
output(2, 77) <= input(26);
output(2, 78) <= input(27);
output(2, 79) <= input(28);
output(2, 80) <= input(38);
output(2, 81) <= input(35);
output(2, 82) <= input(36);
output(2, 83) <= input(32);
output(2, 84) <= input(0);
output(2, 85) <= input(1);
output(2, 86) <= input(2);
output(2, 87) <= input(3);
output(2, 88) <= input(4);
output(2, 89) <= input(5);
output(2, 90) <= input(6);
output(2, 91) <= input(7);
output(2, 92) <= input(8);
output(2, 93) <= input(9);
output(2, 94) <= input(10);
output(2, 95) <= input(11);
output(2, 96) <= input(39);
output(2, 97) <= input(38);
output(2, 98) <= input(35);
output(2, 99) <= input(36);
output(2, 100) <= input(32);
output(2, 101) <= input(0);
output(2, 102) <= input(1);
output(2, 103) <= input(2);
output(2, 104) <= input(3);
output(2, 105) <= input(4);
output(2, 106) <= input(5);
output(2, 107) <= input(6);
output(2, 108) <= input(7);
output(2, 109) <= input(8);
output(2, 110) <= input(9);
output(2, 111) <= input(10);
output(2, 112) <= input(40);
output(2, 113) <= input(41);
output(2, 114) <= input(37);
output(2, 115) <= input(34);
output(2, 116) <= input(33);
output(2, 117) <= input(16);
output(2, 118) <= input(17);
output(2, 119) <= input(18);
output(2, 120) <= input(19);
output(2, 121) <= input(20);
output(2, 122) <= input(21);
output(2, 123) <= input(22);
output(2, 124) <= input(23);
output(2, 125) <= input(24);
output(2, 126) <= input(25);
output(2, 127) <= input(26);
output(2, 128) <= input(43);
output(2, 129) <= input(40);
output(2, 130) <= input(41);
output(2, 131) <= input(37);
output(2, 132) <= input(34);
output(2, 133) <= input(33);
output(2, 134) <= input(16);
output(2, 135) <= input(17);
output(2, 136) <= input(18);
output(2, 137) <= input(19);
output(2, 138) <= input(20);
output(2, 139) <= input(21);
output(2, 140) <= input(22);
output(2, 141) <= input(23);
output(2, 142) <= input(24);
output(2, 143) <= input(25);
output(2, 144) <= input(44);
output(2, 145) <= input(43);
output(2, 146) <= input(40);
output(2, 147) <= input(41);
output(2, 148) <= input(37);
output(2, 149) <= input(34);
output(2, 150) <= input(33);
output(2, 151) <= input(16);
output(2, 152) <= input(17);
output(2, 153) <= input(18);
output(2, 154) <= input(19);
output(2, 155) <= input(20);
output(2, 156) <= input(21);
output(2, 157) <= input(22);
output(2, 158) <= input(23);
output(2, 159) <= input(24);
output(2, 160) <= input(45);
output(2, 161) <= input(46);
output(2, 162) <= input(42);
output(2, 163) <= input(39);
output(2, 164) <= input(38);
output(2, 165) <= input(35);
output(2, 166) <= input(36);
output(2, 167) <= input(32);
output(2, 168) <= input(0);
output(2, 169) <= input(1);
output(2, 170) <= input(2);
output(2, 171) <= input(3);
output(2, 172) <= input(4);
output(2, 173) <= input(5);
output(2, 174) <= input(6);
output(2, 175) <= input(7);
output(2, 176) <= input(48);
output(2, 177) <= input(45);
output(2, 178) <= input(46);
output(2, 179) <= input(42);
output(2, 180) <= input(39);
output(2, 181) <= input(38);
output(2, 182) <= input(35);
output(2, 183) <= input(36);
output(2, 184) <= input(32);
output(2, 185) <= input(0);
output(2, 186) <= input(1);
output(2, 187) <= input(2);
output(2, 188) <= input(3);
output(2, 189) <= input(4);
output(2, 190) <= input(5);
output(2, 191) <= input(6);
output(2, 192) <= input(50);
output(2, 193) <= input(48);
output(2, 194) <= input(45);
output(2, 195) <= input(46);
output(2, 196) <= input(42);
output(2, 197) <= input(39);
output(2, 198) <= input(38);
output(2, 199) <= input(35);
output(2, 200) <= input(36);
output(2, 201) <= input(32);
output(2, 202) <= input(0);
output(2, 203) <= input(1);
output(2, 204) <= input(2);
output(2, 205) <= input(3);
output(2, 206) <= input(4);
output(2, 207) <= input(5);
output(2, 208) <= input(51);
output(2, 209) <= input(49);
output(2, 210) <= input(47);
output(2, 211) <= input(44);
output(2, 212) <= input(43);
output(2, 213) <= input(40);
output(2, 214) <= input(41);
output(2, 215) <= input(37);
output(2, 216) <= input(34);
output(2, 217) <= input(33);
output(2, 218) <= input(16);
output(2, 219) <= input(17);
output(2, 220) <= input(18);
output(2, 221) <= input(19);
output(2, 222) <= input(20);
output(2, 223) <= input(21);
output(2, 224) <= input(52);
output(2, 225) <= input(51);
output(2, 226) <= input(49);
output(2, 227) <= input(47);
output(2, 228) <= input(44);
output(2, 229) <= input(43);
output(2, 230) <= input(40);
output(2, 231) <= input(41);
output(2, 232) <= input(37);
output(2, 233) <= input(34);
output(2, 234) <= input(33);
output(2, 235) <= input(16);
output(2, 236) <= input(17);
output(2, 237) <= input(18);
output(2, 238) <= input(19);
output(2, 239) <= input(20);
output(2, 240) <= input(53);
output(2, 241) <= input(54);
output(2, 242) <= input(50);
output(2, 243) <= input(48);
output(2, 244) <= input(45);
output(2, 245) <= input(46);
output(2, 246) <= input(42);
output(2, 247) <= input(39);
output(2, 248) <= input(38);
output(2, 249) <= input(35);
output(2, 250) <= input(36);
output(2, 251) <= input(32);
output(2, 252) <= input(0);
output(2, 253) <= input(1);
output(2, 254) <= input(2);
output(2, 255) <= input(3);
when "0111" =>
output(0, 0) <= input(0);
output(0, 1) <= input(1);
output(0, 2) <= input(2);
output(0, 3) <= input(3);
output(0, 4) <= input(4);
output(0, 5) <= input(5);
output(0, 6) <= input(6);
output(0, 7) <= input(7);
output(0, 8) <= input(8);
output(0, 9) <= input(9);
output(0, 10) <= input(10);
output(0, 11) <= input(11);
output(0, 12) <= input(12);
output(0, 13) <= input(13);
output(0, 14) <= input(14);
output(0, 15) <= input(15);
output(0, 16) <= input(16);
output(0, 17) <= input(0);
output(0, 18) <= input(1);
output(0, 19) <= input(2);
output(0, 20) <= input(3);
output(0, 21) <= input(4);
output(0, 22) <= input(5);
output(0, 23) <= input(6);
output(0, 24) <= input(7);
output(0, 25) <= input(8);
output(0, 26) <= input(9);
output(0, 27) <= input(10);
output(0, 28) <= input(11);
output(0, 29) <= input(12);
output(0, 30) <= input(13);
output(0, 31) <= input(14);
output(0, 32) <= input(17);
output(0, 33) <= input(16);
output(0, 34) <= input(0);
output(0, 35) <= input(1);
output(0, 36) <= input(2);
output(0, 37) <= input(3);
output(0, 38) <= input(4);
output(0, 39) <= input(5);
output(0, 40) <= input(6);
output(0, 41) <= input(7);
output(0, 42) <= input(8);
output(0, 43) <= input(9);
output(0, 44) <= input(10);
output(0, 45) <= input(11);
output(0, 46) <= input(12);
output(0, 47) <= input(13);
output(0, 48) <= input(18);
output(0, 49) <= input(17);
output(0, 50) <= input(16);
output(0, 51) <= input(0);
output(0, 52) <= input(1);
output(0, 53) <= input(2);
output(0, 54) <= input(3);
output(0, 55) <= input(4);
output(0, 56) <= input(5);
output(0, 57) <= input(6);
output(0, 58) <= input(7);
output(0, 59) <= input(8);
output(0, 60) <= input(9);
output(0, 61) <= input(10);
output(0, 62) <= input(11);
output(0, 63) <= input(12);
output(0, 64) <= input(19);
output(0, 65) <= input(18);
output(0, 66) <= input(17);
output(0, 67) <= input(16);
output(0, 68) <= input(0);
output(0, 69) <= input(1);
output(0, 70) <= input(2);
output(0, 71) <= input(3);
output(0, 72) <= input(4);
output(0, 73) <= input(5);
output(0, 74) <= input(6);
output(0, 75) <= input(7);
output(0, 76) <= input(8);
output(0, 77) <= input(9);
output(0, 78) <= input(10);
output(0, 79) <= input(11);
output(0, 80) <= input(20);
output(0, 81) <= input(21);
output(0, 82) <= input(22);
output(0, 83) <= input(23);
output(0, 84) <= input(24);
output(0, 85) <= input(25);
output(0, 86) <= input(26);
output(0, 87) <= input(27);
output(0, 88) <= input(28);
output(0, 89) <= input(29);
output(0, 90) <= input(30);
output(0, 91) <= input(31);
output(0, 92) <= input(32);
output(0, 93) <= input(33);
output(0, 94) <= input(34);
output(0, 95) <= input(35);
output(0, 96) <= input(36);
output(0, 97) <= input(20);
output(0, 98) <= input(21);
output(0, 99) <= input(22);
output(0, 100) <= input(23);
output(0, 101) <= input(24);
output(0, 102) <= input(25);
output(0, 103) <= input(26);
output(0, 104) <= input(27);
output(0, 105) <= input(28);
output(0, 106) <= input(29);
output(0, 107) <= input(30);
output(0, 108) <= input(31);
output(0, 109) <= input(32);
output(0, 110) <= input(33);
output(0, 111) <= input(34);
output(0, 112) <= input(37);
output(0, 113) <= input(36);
output(0, 114) <= input(20);
output(0, 115) <= input(21);
output(0, 116) <= input(22);
output(0, 117) <= input(23);
output(0, 118) <= input(24);
output(0, 119) <= input(25);
output(0, 120) <= input(26);
output(0, 121) <= input(27);
output(0, 122) <= input(28);
output(0, 123) <= input(29);
output(0, 124) <= input(30);
output(0, 125) <= input(31);
output(0, 126) <= input(32);
output(0, 127) <= input(33);
output(0, 128) <= input(38);
output(0, 129) <= input(37);
output(0, 130) <= input(36);
output(0, 131) <= input(20);
output(0, 132) <= input(21);
output(0, 133) <= input(22);
output(0, 134) <= input(23);
output(0, 135) <= input(24);
output(0, 136) <= input(25);
output(0, 137) <= input(26);
output(0, 138) <= input(27);
output(0, 139) <= input(28);
output(0, 140) <= input(29);
output(0, 141) <= input(30);
output(0, 142) <= input(31);
output(0, 143) <= input(32);
output(0, 144) <= input(39);
output(0, 145) <= input(38);
output(0, 146) <= input(37);
output(0, 147) <= input(36);
output(0, 148) <= input(20);
output(0, 149) <= input(21);
output(0, 150) <= input(22);
output(0, 151) <= input(23);
output(0, 152) <= input(24);
output(0, 153) <= input(25);
output(0, 154) <= input(26);
output(0, 155) <= input(27);
output(0, 156) <= input(28);
output(0, 157) <= input(29);
output(0, 158) <= input(30);
output(0, 159) <= input(31);
output(0, 160) <= input(40);
output(0, 161) <= input(41);
output(0, 162) <= input(42);
output(0, 163) <= input(43);
output(0, 164) <= input(44);
output(0, 165) <= input(19);
output(0, 166) <= input(18);
output(0, 167) <= input(17);
output(0, 168) <= input(16);
output(0, 169) <= input(0);
output(0, 170) <= input(1);
output(0, 171) <= input(2);
output(0, 172) <= input(3);
output(0, 173) <= input(4);
output(0, 174) <= input(5);
output(0, 175) <= input(6);
output(0, 176) <= input(45);
output(0, 177) <= input(40);
output(0, 178) <= input(41);
output(0, 179) <= input(42);
output(0, 180) <= input(43);
output(0, 181) <= input(44);
output(0, 182) <= input(19);
output(0, 183) <= input(18);
output(0, 184) <= input(17);
output(0, 185) <= input(16);
output(0, 186) <= input(0);
output(0, 187) <= input(1);
output(0, 188) <= input(2);
output(0, 189) <= input(3);
output(0, 190) <= input(4);
output(0, 191) <= input(5);
output(0, 192) <= input(46);
output(0, 193) <= input(45);
output(0, 194) <= input(40);
output(0, 195) <= input(41);
output(0, 196) <= input(42);
output(0, 197) <= input(43);
output(0, 198) <= input(44);
output(0, 199) <= input(19);
output(0, 200) <= input(18);
output(0, 201) <= input(17);
output(0, 202) <= input(16);
output(0, 203) <= input(0);
output(0, 204) <= input(1);
output(0, 205) <= input(2);
output(0, 206) <= input(3);
output(0, 207) <= input(4);
output(0, 208) <= input(47);
output(0, 209) <= input(46);
output(0, 210) <= input(45);
output(0, 211) <= input(40);
output(0, 212) <= input(41);
output(0, 213) <= input(42);
output(0, 214) <= input(43);
output(0, 215) <= input(44);
output(0, 216) <= input(19);
output(0, 217) <= input(18);
output(0, 218) <= input(17);
output(0, 219) <= input(16);
output(0, 220) <= input(0);
output(0, 221) <= input(1);
output(0, 222) <= input(2);
output(0, 223) <= input(3);
output(0, 224) <= input(48);
output(0, 225) <= input(47);
output(0, 226) <= input(46);
output(0, 227) <= input(45);
output(0, 228) <= input(40);
output(0, 229) <= input(41);
output(0, 230) <= input(42);
output(0, 231) <= input(43);
output(0, 232) <= input(44);
output(0, 233) <= input(19);
output(0, 234) <= input(18);
output(0, 235) <= input(17);
output(0, 236) <= input(16);
output(0, 237) <= input(0);
output(0, 238) <= input(1);
output(0, 239) <= input(2);
output(0, 240) <= input(49);
output(0, 241) <= input(50);
output(0, 242) <= input(51);
output(0, 243) <= input(52);
output(0, 244) <= input(53);
output(0, 245) <= input(39);
output(0, 246) <= input(38);
output(0, 247) <= input(37);
output(0, 248) <= input(36);
output(0, 249) <= input(20);
output(0, 250) <= input(21);
output(0, 251) <= input(22);
output(0, 252) <= input(23);
output(0, 253) <= input(24);
output(0, 254) <= input(25);
output(0, 255) <= input(26);
output(1, 0) <= input(54);
output(1, 1) <= input(55);
output(1, 2) <= input(56);
output(1, 3) <= input(57);
output(1, 4) <= input(58);
output(1, 5) <= input(59);
output(1, 6) <= input(60);
output(1, 7) <= input(61);
output(1, 8) <= input(62);
output(1, 9) <= input(63);
output(1, 10) <= input(64);
output(1, 11) <= input(65);
output(1, 12) <= input(66);
output(1, 13) <= input(67);
output(1, 14) <= input(68);
output(1, 15) <= input(69);
output(1, 16) <= input(70);
output(1, 17) <= input(54);
output(1, 18) <= input(55);
output(1, 19) <= input(56);
output(1, 20) <= input(57);
output(1, 21) <= input(58);
output(1, 22) <= input(59);
output(1, 23) <= input(60);
output(1, 24) <= input(61);
output(1, 25) <= input(62);
output(1, 26) <= input(63);
output(1, 27) <= input(64);
output(1, 28) <= input(65);
output(1, 29) <= input(66);
output(1, 30) <= input(67);
output(1, 31) <= input(68);
output(1, 32) <= input(71);
output(1, 33) <= input(70);
output(1, 34) <= input(54);
output(1, 35) <= input(55);
output(1, 36) <= input(56);
output(1, 37) <= input(57);
output(1, 38) <= input(58);
output(1, 39) <= input(59);
output(1, 40) <= input(60);
output(1, 41) <= input(61);
output(1, 42) <= input(62);
output(1, 43) <= input(63);
output(1, 44) <= input(64);
output(1, 45) <= input(65);
output(1, 46) <= input(66);
output(1, 47) <= input(67);
output(1, 48) <= input(72);
output(1, 49) <= input(71);
output(1, 50) <= input(70);
output(1, 51) <= input(54);
output(1, 52) <= input(55);
output(1, 53) <= input(56);
output(1, 54) <= input(57);
output(1, 55) <= input(58);
output(1, 56) <= input(59);
output(1, 57) <= input(60);
output(1, 58) <= input(61);
output(1, 59) <= input(62);
output(1, 60) <= input(63);
output(1, 61) <= input(64);
output(1, 62) <= input(65);
output(1, 63) <= input(66);
output(1, 64) <= input(73);
output(1, 65) <= input(72);
output(1, 66) <= input(71);
output(1, 67) <= input(70);
output(1, 68) <= input(54);
output(1, 69) <= input(55);
output(1, 70) <= input(56);
output(1, 71) <= input(57);
output(1, 72) <= input(58);
output(1, 73) <= input(59);
output(1, 74) <= input(60);
output(1, 75) <= input(61);
output(1, 76) <= input(62);
output(1, 77) <= input(63);
output(1, 78) <= input(64);
output(1, 79) <= input(65);
output(1, 80) <= input(74);
output(1, 81) <= input(73);
output(1, 82) <= input(72);
output(1, 83) <= input(71);
output(1, 84) <= input(70);
output(1, 85) <= input(54);
output(1, 86) <= input(55);
output(1, 87) <= input(56);
output(1, 88) <= input(57);
output(1, 89) <= input(58);
output(1, 90) <= input(59);
output(1, 91) <= input(60);
output(1, 92) <= input(61);
output(1, 93) <= input(62);
output(1, 94) <= input(63);
output(1, 95) <= input(64);
output(1, 96) <= input(75);
output(1, 97) <= input(74);
output(1, 98) <= input(73);
output(1, 99) <= input(72);
output(1, 100) <= input(71);
output(1, 101) <= input(70);
output(1, 102) <= input(54);
output(1, 103) <= input(55);
output(1, 104) <= input(56);
output(1, 105) <= input(57);
output(1, 106) <= input(58);
output(1, 107) <= input(59);
output(1, 108) <= input(60);
output(1, 109) <= input(61);
output(1, 110) <= input(62);
output(1, 111) <= input(63);
output(1, 112) <= input(76);
output(1, 113) <= input(75);
output(1, 114) <= input(74);
output(1, 115) <= input(73);
output(1, 116) <= input(72);
output(1, 117) <= input(71);
output(1, 118) <= input(70);
output(1, 119) <= input(54);
output(1, 120) <= input(55);
output(1, 121) <= input(56);
output(1, 122) <= input(57);
output(1, 123) <= input(58);
output(1, 124) <= input(59);
output(1, 125) <= input(60);
output(1, 126) <= input(61);
output(1, 127) <= input(62);
output(1, 128) <= input(77);
output(1, 129) <= input(76);
output(1, 130) <= input(75);
output(1, 131) <= input(74);
output(1, 132) <= input(73);
output(1, 133) <= input(72);
output(1, 134) <= input(71);
output(1, 135) <= input(70);
output(1, 136) <= input(54);
output(1, 137) <= input(55);
output(1, 138) <= input(56);
output(1, 139) <= input(57);
output(1, 140) <= input(58);
output(1, 141) <= input(59);
output(1, 142) <= input(60);
output(1, 143) <= input(61);
output(1, 144) <= input(78);
output(1, 145) <= input(77);
output(1, 146) <= input(76);
output(1, 147) <= input(75);
output(1, 148) <= input(74);
output(1, 149) <= input(73);
output(1, 150) <= input(72);
output(1, 151) <= input(71);
output(1, 152) <= input(70);
output(1, 153) <= input(54);
output(1, 154) <= input(55);
output(1, 155) <= input(56);
output(1, 156) <= input(57);
output(1, 157) <= input(58);
output(1, 158) <= input(59);
output(1, 159) <= input(60);
output(1, 160) <= input(79);
output(1, 161) <= input(78);
output(1, 162) <= input(77);
output(1, 163) <= input(76);
output(1, 164) <= input(75);
output(1, 165) <= input(74);
output(1, 166) <= input(73);
output(1, 167) <= input(72);
output(1, 168) <= input(71);
output(1, 169) <= input(70);
output(1, 170) <= input(54);
output(1, 171) <= input(55);
output(1, 172) <= input(56);
output(1, 173) <= input(57);
output(1, 174) <= input(58);
output(1, 175) <= input(59);
output(1, 176) <= input(80);
output(1, 177) <= input(79);
output(1, 178) <= input(78);
output(1, 179) <= input(77);
output(1, 180) <= input(76);
output(1, 181) <= input(75);
output(1, 182) <= input(74);
output(1, 183) <= input(73);
output(1, 184) <= input(72);
output(1, 185) <= input(71);
output(1, 186) <= input(70);
output(1, 187) <= input(54);
output(1, 188) <= input(55);
output(1, 189) <= input(56);
output(1, 190) <= input(57);
output(1, 191) <= input(58);
output(1, 192) <= input(81);
output(1, 193) <= input(80);
output(1, 194) <= input(79);
output(1, 195) <= input(78);
output(1, 196) <= input(77);
output(1, 197) <= input(76);
output(1, 198) <= input(75);
output(1, 199) <= input(74);
output(1, 200) <= input(73);
output(1, 201) <= input(72);
output(1, 202) <= input(71);
output(1, 203) <= input(70);
output(1, 204) <= input(54);
output(1, 205) <= input(55);
output(1, 206) <= input(56);
output(1, 207) <= input(57);
output(1, 208) <= input(82);
output(1, 209) <= input(81);
output(1, 210) <= input(80);
output(1, 211) <= input(79);
output(1, 212) <= input(78);
output(1, 213) <= input(77);
output(1, 214) <= input(76);
output(1, 215) <= input(75);
output(1, 216) <= input(74);
output(1, 217) <= input(73);
output(1, 218) <= input(72);
output(1, 219) <= input(71);
output(1, 220) <= input(70);
output(1, 221) <= input(54);
output(1, 222) <= input(55);
output(1, 223) <= input(56);
output(1, 224) <= input(83);
output(1, 225) <= input(82);
output(1, 226) <= input(81);
output(1, 227) <= input(80);
output(1, 228) <= input(79);
output(1, 229) <= input(78);
output(1, 230) <= input(77);
output(1, 231) <= input(76);
output(1, 232) <= input(75);
output(1, 233) <= input(74);
output(1, 234) <= input(73);
output(1, 235) <= input(72);
output(1, 236) <= input(71);
output(1, 237) <= input(70);
output(1, 238) <= input(54);
output(1, 239) <= input(55);
output(1, 240) <= input(84);
output(1, 241) <= input(83);
output(1, 242) <= input(82);
output(1, 243) <= input(81);
output(1, 244) <= input(80);
output(1, 245) <= input(79);
output(1, 246) <= input(78);
output(1, 247) <= input(77);
output(1, 248) <= input(76);
output(1, 249) <= input(75);
output(1, 250) <= input(74);
output(1, 251) <= input(73);
output(1, 252) <= input(72);
output(1, 253) <= input(71);
output(1, 254) <= input(70);
output(1, 255) <= input(54);
when "1000" =>
output(0, 0) <= input(0);
output(0, 1) <= input(1);
output(0, 2) <= input(2);
output(0, 3) <= input(3);
output(0, 4) <= input(4);
output(0, 5) <= input(5);
output(0, 6) <= input(6);
output(0, 7) <= input(7);
output(0, 8) <= input(8);
output(0, 9) <= input(9);
output(0, 10) <= input(10);
output(0, 11) <= input(11);
output(0, 12) <= input(12);
output(0, 13) <= input(13);
output(0, 14) <= input(14);
output(0, 15) <= input(15);
output(0, 16) <= input(16);
output(0, 17) <= input(0);
output(0, 18) <= input(1);
output(0, 19) <= input(2);
output(0, 20) <= input(3);
output(0, 21) <= input(4);
output(0, 22) <= input(5);
output(0, 23) <= input(6);
output(0, 24) <= input(7);
output(0, 25) <= input(8);
output(0, 26) <= input(9);
output(0, 27) <= input(10);
output(0, 28) <= input(11);
output(0, 29) <= input(12);
output(0, 30) <= input(13);
output(0, 31) <= input(14);
output(0, 32) <= input(17);
output(0, 33) <= input(16);
output(0, 34) <= input(0);
output(0, 35) <= input(1);
output(0, 36) <= input(2);
output(0, 37) <= input(3);
output(0, 38) <= input(4);
output(0, 39) <= input(5);
output(0, 40) <= input(6);
output(0, 41) <= input(7);
output(0, 42) <= input(8);
output(0, 43) <= input(9);
output(0, 44) <= input(10);
output(0, 45) <= input(11);
output(0, 46) <= input(12);
output(0, 47) <= input(13);
output(0, 48) <= input(18);
output(0, 49) <= input(17);
output(0, 50) <= input(16);
output(0, 51) <= input(0);
output(0, 52) <= input(1);
output(0, 53) <= input(2);
output(0, 54) <= input(3);
output(0, 55) <= input(4);
output(0, 56) <= input(5);
output(0, 57) <= input(6);
output(0, 58) <= input(7);
output(0, 59) <= input(8);
output(0, 60) <= input(9);
output(0, 61) <= input(10);
output(0, 62) <= input(11);
output(0, 63) <= input(12);
output(0, 64) <= input(19);
output(0, 65) <= input(18);
output(0, 66) <= input(17);
output(0, 67) <= input(16);
output(0, 68) <= input(0);
output(0, 69) <= input(1);
output(0, 70) <= input(2);
output(0, 71) <= input(3);
output(0, 72) <= input(4);
output(0, 73) <= input(5);
output(0, 74) <= input(6);
output(0, 75) <= input(7);
output(0, 76) <= input(8);
output(0, 77) <= input(9);
output(0, 78) <= input(10);
output(0, 79) <= input(11);
output(0, 80) <= input(20);
output(0, 81) <= input(21);
output(0, 82) <= input(22);
output(0, 83) <= input(23);
output(0, 84) <= input(24);
output(0, 85) <= input(25);
output(0, 86) <= input(26);
output(0, 87) <= input(27);
output(0, 88) <= input(28);
output(0, 89) <= input(29);
output(0, 90) <= input(30);
output(0, 91) <= input(31);
output(0, 92) <= input(32);
output(0, 93) <= input(33);
output(0, 94) <= input(34);
output(0, 95) <= input(35);
output(0, 96) <= input(36);
output(0, 97) <= input(20);
output(0, 98) <= input(21);
output(0, 99) <= input(22);
output(0, 100) <= input(23);
output(0, 101) <= input(24);
output(0, 102) <= input(25);
output(0, 103) <= input(26);
output(0, 104) <= input(27);
output(0, 105) <= input(28);
output(0, 106) <= input(29);
output(0, 107) <= input(30);
output(0, 108) <= input(31);
output(0, 109) <= input(32);
output(0, 110) <= input(33);
output(0, 111) <= input(34);
output(0, 112) <= input(37);
output(0, 113) <= input(36);
output(0, 114) <= input(20);
output(0, 115) <= input(21);
output(0, 116) <= input(22);
output(0, 117) <= input(23);
output(0, 118) <= input(24);
output(0, 119) <= input(25);
output(0, 120) <= input(26);
output(0, 121) <= input(27);
output(0, 122) <= input(28);
output(0, 123) <= input(29);
output(0, 124) <= input(30);
output(0, 125) <= input(31);
output(0, 126) <= input(32);
output(0, 127) <= input(33);
output(0, 128) <= input(38);
output(0, 129) <= input(37);
output(0, 130) <= input(36);
output(0, 131) <= input(20);
output(0, 132) <= input(21);
output(0, 133) <= input(22);
output(0, 134) <= input(23);
output(0, 135) <= input(24);
output(0, 136) <= input(25);
output(0, 137) <= input(26);
output(0, 138) <= input(27);
output(0, 139) <= input(28);
output(0, 140) <= input(29);
output(0, 141) <= input(30);
output(0, 142) <= input(31);
output(0, 143) <= input(32);
output(0, 144) <= input(39);
output(0, 145) <= input(38);
output(0, 146) <= input(37);
output(0, 147) <= input(36);
output(0, 148) <= input(20);
output(0, 149) <= input(21);
output(0, 150) <= input(22);
output(0, 151) <= input(23);
output(0, 152) <= input(24);
output(0, 153) <= input(25);
output(0, 154) <= input(26);
output(0, 155) <= input(27);
output(0, 156) <= input(28);
output(0, 157) <= input(29);
output(0, 158) <= input(30);
output(0, 159) <= input(31);
output(0, 160) <= input(40);
output(0, 161) <= input(41);
output(0, 162) <= input(42);
output(0, 163) <= input(43);
output(0, 164) <= input(44);
output(0, 165) <= input(19);
output(0, 166) <= input(18);
output(0, 167) <= input(17);
output(0, 168) <= input(16);
output(0, 169) <= input(0);
output(0, 170) <= input(1);
output(0, 171) <= input(2);
output(0, 172) <= input(3);
output(0, 173) <= input(4);
output(0, 174) <= input(5);
output(0, 175) <= input(6);
output(0, 176) <= input(45);
output(0, 177) <= input(40);
output(0, 178) <= input(41);
output(0, 179) <= input(42);
output(0, 180) <= input(43);
output(0, 181) <= input(44);
output(0, 182) <= input(19);
output(0, 183) <= input(18);
output(0, 184) <= input(17);
output(0, 185) <= input(16);
output(0, 186) <= input(0);
output(0, 187) <= input(1);
output(0, 188) <= input(2);
output(0, 189) <= input(3);
output(0, 190) <= input(4);
output(0, 191) <= input(5);
output(0, 192) <= input(46);
output(0, 193) <= input(45);
output(0, 194) <= input(40);
output(0, 195) <= input(41);
output(0, 196) <= input(42);
output(0, 197) <= input(43);
output(0, 198) <= input(44);
output(0, 199) <= input(19);
output(0, 200) <= input(18);
output(0, 201) <= input(17);
output(0, 202) <= input(16);
output(0, 203) <= input(0);
output(0, 204) <= input(1);
output(0, 205) <= input(2);
output(0, 206) <= input(3);
output(0, 207) <= input(4);
output(0, 208) <= input(47);
output(0, 209) <= input(46);
output(0, 210) <= input(45);
output(0, 211) <= input(40);
output(0, 212) <= input(41);
output(0, 213) <= input(42);
output(0, 214) <= input(43);
output(0, 215) <= input(44);
output(0, 216) <= input(19);
output(0, 217) <= input(18);
output(0, 218) <= input(17);
output(0, 219) <= input(16);
output(0, 220) <= input(0);
output(0, 221) <= input(1);
output(0, 222) <= input(2);
output(0, 223) <= input(3);
output(0, 224) <= input(48);
output(0, 225) <= input(47);
output(0, 226) <= input(46);
output(0, 227) <= input(45);
output(0, 228) <= input(40);
output(0, 229) <= input(41);
output(0, 230) <= input(42);
output(0, 231) <= input(43);
output(0, 232) <= input(44);
output(0, 233) <= input(19);
output(0, 234) <= input(18);
output(0, 235) <= input(17);
output(0, 236) <= input(16);
output(0, 237) <= input(0);
output(0, 238) <= input(1);
output(0, 239) <= input(2);
output(0, 240) <= input(49);
output(0, 241) <= input(50);
output(0, 242) <= input(51);
output(0, 243) <= input(52);
output(0, 244) <= input(53);
output(0, 245) <= input(39);
output(0, 246) <= input(38);
output(0, 247) <= input(37);
output(0, 248) <= input(36);
output(0, 249) <= input(20);
output(0, 250) <= input(21);
output(0, 251) <= input(22);
output(0, 252) <= input(23);
output(0, 253) <= input(24);
output(0, 254) <= input(25);
output(0, 255) <= input(26);
when "1001" =>
output(0, 0) <= input(0);
output(0, 1) <= input(1);
output(0, 2) <= input(2);
output(0, 3) <= input(3);
output(0, 4) <= input(4);
output(0, 5) <= input(5);
output(0, 6) <= input(6);
output(0, 7) <= input(7);
output(0, 8) <= input(8);
output(0, 9) <= input(9);
output(0, 10) <= input(10);
output(0, 11) <= input(11);
output(0, 12) <= input(12);
output(0, 13) <= input(13);
output(0, 14) <= input(14);
output(0, 15) <= input(15);
output(0, 16) <= input(16);
output(0, 17) <= input(0);
output(0, 18) <= input(1);
output(0, 19) <= input(2);
output(0, 20) <= input(3);
output(0, 21) <= input(4);
output(0, 22) <= input(5);
output(0, 23) <= input(6);
output(0, 24) <= input(7);
output(0, 25) <= input(8);
output(0, 26) <= input(9);
output(0, 27) <= input(10);
output(0, 28) <= input(11);
output(0, 29) <= input(12);
output(0, 30) <= input(13);
output(0, 31) <= input(14);
output(0, 32) <= input(17);
output(0, 33) <= input(18);
output(0, 34) <= input(19);
output(0, 35) <= input(20);
output(0, 36) <= input(21);
output(0, 37) <= input(22);
output(0, 38) <= input(23);
output(0, 39) <= input(24);
output(0, 40) <= input(25);
output(0, 41) <= input(26);
output(0, 42) <= input(27);
output(0, 43) <= input(28);
output(0, 44) <= input(29);
output(0, 45) <= input(30);
output(0, 46) <= input(31);
output(0, 47) <= input(32);
output(0, 48) <= input(33);
output(0, 49) <= input(17);
output(0, 50) <= input(18);
output(0, 51) <= input(19);
output(0, 52) <= input(20);
output(0, 53) <= input(21);
output(0, 54) <= input(22);
output(0, 55) <= input(23);
output(0, 56) <= input(24);
output(0, 57) <= input(25);
output(0, 58) <= input(26);
output(0, 59) <= input(27);
output(0, 60) <= input(28);
output(0, 61) <= input(29);
output(0, 62) <= input(30);
output(0, 63) <= input(31);
output(0, 64) <= input(34);
output(0, 65) <= input(33);
output(0, 66) <= input(17);
output(0, 67) <= input(18);
output(0, 68) <= input(19);
output(0, 69) <= input(20);
output(0, 70) <= input(21);
output(0, 71) <= input(22);
output(0, 72) <= input(23);
output(0, 73) <= input(24);
output(0, 74) <= input(25);
output(0, 75) <= input(26);
output(0, 76) <= input(27);
output(0, 77) <= input(28);
output(0, 78) <= input(29);
output(0, 79) <= input(30);
output(0, 80) <= input(35);
output(0, 81) <= input(36);
output(0, 82) <= input(37);
output(0, 83) <= input(16);
output(0, 84) <= input(0);
output(0, 85) <= input(1);
output(0, 86) <= input(2);
output(0, 87) <= input(3);
output(0, 88) <= input(4);
output(0, 89) <= input(5);
output(0, 90) <= input(6);
output(0, 91) <= input(7);
output(0, 92) <= input(8);
output(0, 93) <= input(9);
output(0, 94) <= input(10);
output(0, 95) <= input(11);
output(0, 96) <= input(38);
output(0, 97) <= input(35);
output(0, 98) <= input(36);
output(0, 99) <= input(37);
output(0, 100) <= input(16);
output(0, 101) <= input(0);
output(0, 102) <= input(1);
output(0, 103) <= input(2);
output(0, 104) <= input(3);
output(0, 105) <= input(4);
output(0, 106) <= input(5);
output(0, 107) <= input(6);
output(0, 108) <= input(7);
output(0, 109) <= input(8);
output(0, 110) <= input(9);
output(0, 111) <= input(10);
output(0, 112) <= input(39);
output(0, 113) <= input(40);
output(0, 114) <= input(34);
output(0, 115) <= input(33);
output(0, 116) <= input(17);
output(0, 117) <= input(18);
output(0, 118) <= input(19);
output(0, 119) <= input(20);
output(0, 120) <= input(21);
output(0, 121) <= input(22);
output(0, 122) <= input(23);
output(0, 123) <= input(24);
output(0, 124) <= input(25);
output(0, 125) <= input(26);
output(0, 126) <= input(27);
output(0, 127) <= input(28);
output(0, 128) <= input(41);
output(0, 129) <= input(39);
output(0, 130) <= input(40);
output(0, 131) <= input(34);
output(0, 132) <= input(33);
output(0, 133) <= input(17);
output(0, 134) <= input(18);
output(0, 135) <= input(19);
output(0, 136) <= input(20);
output(0, 137) <= input(21);
output(0, 138) <= input(22);
output(0, 139) <= input(23);
output(0, 140) <= input(24);
output(0, 141) <= input(25);
output(0, 142) <= input(26);
output(0, 143) <= input(27);
output(0, 144) <= input(42);
output(0, 145) <= input(41);
output(0, 146) <= input(39);
output(0, 147) <= input(40);
output(0, 148) <= input(34);
output(0, 149) <= input(33);
output(0, 150) <= input(17);
output(0, 151) <= input(18);
output(0, 152) <= input(19);
output(0, 153) <= input(20);
output(0, 154) <= input(21);
output(0, 155) <= input(22);
output(0, 156) <= input(23);
output(0, 157) <= input(24);
output(0, 158) <= input(25);
output(0, 159) <= input(26);
output(0, 160) <= input(43);
output(0, 161) <= input(44);
output(0, 162) <= input(45);
output(0, 163) <= input(38);
output(0, 164) <= input(35);
output(0, 165) <= input(36);
output(0, 166) <= input(37);
output(0, 167) <= input(16);
output(0, 168) <= input(0);
output(0, 169) <= input(1);
output(0, 170) <= input(2);
output(0, 171) <= input(3);
output(0, 172) <= input(4);
output(0, 173) <= input(5);
output(0, 174) <= input(6);
output(0, 175) <= input(7);
output(0, 176) <= input(46);
output(0, 177) <= input(43);
output(0, 178) <= input(44);
output(0, 179) <= input(45);
output(0, 180) <= input(38);
output(0, 181) <= input(35);
output(0, 182) <= input(36);
output(0, 183) <= input(37);
output(0, 184) <= input(16);
output(0, 185) <= input(0);
output(0, 186) <= input(1);
output(0, 187) <= input(2);
output(0, 188) <= input(3);
output(0, 189) <= input(4);
output(0, 190) <= input(5);
output(0, 191) <= input(6);
output(0, 192) <= input(47);
output(0, 193) <= input(46);
output(0, 194) <= input(43);
output(0, 195) <= input(44);
output(0, 196) <= input(45);
output(0, 197) <= input(38);
output(0, 198) <= input(35);
output(0, 199) <= input(36);
output(0, 200) <= input(37);
output(0, 201) <= input(16);
output(0, 202) <= input(0);
output(0, 203) <= input(1);
output(0, 204) <= input(2);
output(0, 205) <= input(3);
output(0, 206) <= input(4);
output(0, 207) <= input(5);
output(0, 208) <= input(48);
output(0, 209) <= input(49);
output(0, 210) <= input(50);
output(0, 211) <= input(42);
output(0, 212) <= input(41);
output(0, 213) <= input(39);
output(0, 214) <= input(40);
output(0, 215) <= input(34);
output(0, 216) <= input(33);
output(0, 217) <= input(17);
output(0, 218) <= input(18);
output(0, 219) <= input(19);
output(0, 220) <= input(20);
output(0, 221) <= input(21);
output(0, 222) <= input(22);
output(0, 223) <= input(23);
output(0, 224) <= input(51);
output(0, 225) <= input(48);
output(0, 226) <= input(49);
output(0, 227) <= input(50);
output(0, 228) <= input(42);
output(0, 229) <= input(41);
output(0, 230) <= input(39);
output(0, 231) <= input(40);
output(0, 232) <= input(34);
output(0, 233) <= input(33);
output(0, 234) <= input(17);
output(0, 235) <= input(18);
output(0, 236) <= input(19);
output(0, 237) <= input(20);
output(0, 238) <= input(21);
output(0, 239) <= input(22);
output(0, 240) <= input(52);
output(0, 241) <= input(53);
output(0, 242) <= input(47);
output(0, 243) <= input(46);
output(0, 244) <= input(43);
output(0, 245) <= input(44);
output(0, 246) <= input(45);
output(0, 247) <= input(38);
output(0, 248) <= input(35);
output(0, 249) <= input(36);
output(0, 250) <= input(37);
output(0, 251) <= input(16);
output(0, 252) <= input(0);
output(0, 253) <= input(1);
output(0, 254) <= input(2);
output(0, 255) <= input(3);
output(1, 0) <= input(0);
output(1, 1) <= input(1);
output(1, 2) <= input(2);
output(1, 3) <= input(3);
output(1, 4) <= input(4);
output(1, 5) <= input(5);
output(1, 6) <= input(6);
output(1, 7) <= input(7);
output(1, 8) <= input(8);
output(1, 9) <= input(9);
output(1, 10) <= input(10);
output(1, 11) <= input(11);
output(1, 12) <= input(12);
output(1, 13) <= input(13);
output(1, 14) <= input(14);
output(1, 15) <= input(15);
output(1, 16) <= input(18);
output(1, 17) <= input(19);
output(1, 18) <= input(20);
output(1, 19) <= input(21);
output(1, 20) <= input(22);
output(1, 21) <= input(23);
output(1, 22) <= input(24);
output(1, 23) <= input(25);
output(1, 24) <= input(26);
output(1, 25) <= input(27);
output(1, 26) <= input(28);
output(1, 27) <= input(29);
output(1, 28) <= input(30);
output(1, 29) <= input(31);
output(1, 30) <= input(32);
output(1, 31) <= input(54);
output(1, 32) <= input(17);
output(1, 33) <= input(18);
output(1, 34) <= input(19);
output(1, 35) <= input(20);
output(1, 36) <= input(21);
output(1, 37) <= input(22);
output(1, 38) <= input(23);
output(1, 39) <= input(24);
output(1, 40) <= input(25);
output(1, 41) <= input(26);
output(1, 42) <= input(27);
output(1, 43) <= input(28);
output(1, 44) <= input(29);
output(1, 45) <= input(30);
output(1, 46) <= input(31);
output(1, 47) <= input(32);
output(1, 48) <= input(37);
output(1, 49) <= input(16);
output(1, 50) <= input(0);
output(1, 51) <= input(1);
output(1, 52) <= input(2);
output(1, 53) <= input(3);
output(1, 54) <= input(4);
output(1, 55) <= input(5);
output(1, 56) <= input(6);
output(1, 57) <= input(7);
output(1, 58) <= input(8);
output(1, 59) <= input(9);
output(1, 60) <= input(10);
output(1, 61) <= input(11);
output(1, 62) <= input(12);
output(1, 63) <= input(13);
output(1, 64) <= input(36);
output(1, 65) <= input(37);
output(1, 66) <= input(16);
output(1, 67) <= input(0);
output(1, 68) <= input(1);
output(1, 69) <= input(2);
output(1, 70) <= input(3);
output(1, 71) <= input(4);
output(1, 72) <= input(5);
output(1, 73) <= input(6);
output(1, 74) <= input(7);
output(1, 75) <= input(8);
output(1, 76) <= input(9);
output(1, 77) <= input(10);
output(1, 78) <= input(11);
output(1, 79) <= input(12);
output(1, 80) <= input(34);
output(1, 81) <= input(33);
output(1, 82) <= input(17);
output(1, 83) <= input(18);
output(1, 84) <= input(19);
output(1, 85) <= input(20);
output(1, 86) <= input(21);
output(1, 87) <= input(22);
output(1, 88) <= input(23);
output(1, 89) <= input(24);
output(1, 90) <= input(25);
output(1, 91) <= input(26);
output(1, 92) <= input(27);
output(1, 93) <= input(28);
output(1, 94) <= input(29);
output(1, 95) <= input(30);
output(1, 96) <= input(40);
output(1, 97) <= input(34);
output(1, 98) <= input(33);
output(1, 99) <= input(17);
output(1, 100) <= input(18);
output(1, 101) <= input(19);
output(1, 102) <= input(20);
output(1, 103) <= input(21);
output(1, 104) <= input(22);
output(1, 105) <= input(23);
output(1, 106) <= input(24);
output(1, 107) <= input(25);
output(1, 108) <= input(26);
output(1, 109) <= input(27);
output(1, 110) <= input(28);
output(1, 111) <= input(29);
output(1, 112) <= input(38);
output(1, 113) <= input(35);
output(1, 114) <= input(36);
output(1, 115) <= input(37);
output(1, 116) <= input(16);
output(1, 117) <= input(0);
output(1, 118) <= input(1);
output(1, 119) <= input(2);
output(1, 120) <= input(3);
output(1, 121) <= input(4);
output(1, 122) <= input(5);
output(1, 123) <= input(6);
output(1, 124) <= input(7);
output(1, 125) <= input(8);
output(1, 126) <= input(9);
output(1, 127) <= input(10);
output(1, 128) <= input(39);
output(1, 129) <= input(40);
output(1, 130) <= input(34);
output(1, 131) <= input(33);
output(1, 132) <= input(17);
output(1, 133) <= input(18);
output(1, 134) <= input(19);
output(1, 135) <= input(20);
output(1, 136) <= input(21);
output(1, 137) <= input(22);
output(1, 138) <= input(23);
output(1, 139) <= input(24);
output(1, 140) <= input(25);
output(1, 141) <= input(26);
output(1, 142) <= input(27);
output(1, 143) <= input(28);
output(1, 144) <= input(41);
output(1, 145) <= input(39);
output(1, 146) <= input(40);
output(1, 147) <= input(34);
output(1, 148) <= input(33);
output(1, 149) <= input(17);
output(1, 150) <= input(18);
output(1, 151) <= input(19);
output(1, 152) <= input(20);
output(1, 153) <= input(21);
output(1, 154) <= input(22);
output(1, 155) <= input(23);
output(1, 156) <= input(24);
output(1, 157) <= input(25);
output(1, 158) <= input(26);
output(1, 159) <= input(27);
output(1, 160) <= input(44);
output(1, 161) <= input(45);
output(1, 162) <= input(38);
output(1, 163) <= input(35);
output(1, 164) <= input(36);
output(1, 165) <= input(37);
output(1, 166) <= input(16);
output(1, 167) <= input(0);
output(1, 168) <= input(1);
output(1, 169) <= input(2);
output(1, 170) <= input(3);
output(1, 171) <= input(4);
output(1, 172) <= input(5);
output(1, 173) <= input(6);
output(1, 174) <= input(7);
output(1, 175) <= input(8);
output(1, 176) <= input(43);
output(1, 177) <= input(44);
output(1, 178) <= input(45);
output(1, 179) <= input(38);
output(1, 180) <= input(35);
output(1, 181) <= input(36);
output(1, 182) <= input(37);
output(1, 183) <= input(16);
output(1, 184) <= input(0);
output(1, 185) <= input(1);
output(1, 186) <= input(2);
output(1, 187) <= input(3);
output(1, 188) <= input(4);
output(1, 189) <= input(5);
output(1, 190) <= input(6);
output(1, 191) <= input(7);
output(1, 192) <= input(50);
output(1, 193) <= input(42);
output(1, 194) <= input(41);
output(1, 195) <= input(39);
output(1, 196) <= input(40);
output(1, 197) <= input(34);
output(1, 198) <= input(33);
output(1, 199) <= input(17);
output(1, 200) <= input(18);
output(1, 201) <= input(19);
output(1, 202) <= input(20);
output(1, 203) <= input(21);
output(1, 204) <= input(22);
output(1, 205) <= input(23);
output(1, 206) <= input(24);
output(1, 207) <= input(25);
output(1, 208) <= input(49);
output(1, 209) <= input(50);
output(1, 210) <= input(42);
output(1, 211) <= input(41);
output(1, 212) <= input(39);
output(1, 213) <= input(40);
output(1, 214) <= input(34);
output(1, 215) <= input(33);
output(1, 216) <= input(17);
output(1, 217) <= input(18);
output(1, 218) <= input(19);
output(1, 219) <= input(20);
output(1, 220) <= input(21);
output(1, 221) <= input(22);
output(1, 222) <= input(23);
output(1, 223) <= input(24);
output(1, 224) <= input(47);
output(1, 225) <= input(46);
output(1, 226) <= input(43);
output(1, 227) <= input(44);
output(1, 228) <= input(45);
output(1, 229) <= input(38);
output(1, 230) <= input(35);
output(1, 231) <= input(36);
output(1, 232) <= input(37);
output(1, 233) <= input(16);
output(1, 234) <= input(0);
output(1, 235) <= input(1);
output(1, 236) <= input(2);
output(1, 237) <= input(3);
output(1, 238) <= input(4);
output(1, 239) <= input(5);
output(1, 240) <= input(48);
output(1, 241) <= input(49);
output(1, 242) <= input(50);
output(1, 243) <= input(42);
output(1, 244) <= input(41);
output(1, 245) <= input(39);
output(1, 246) <= input(40);
output(1, 247) <= input(34);
output(1, 248) <= input(33);
output(1, 249) <= input(17);
output(1, 250) <= input(18);
output(1, 251) <= input(19);
output(1, 252) <= input(20);
output(1, 253) <= input(21);
output(1, 254) <= input(22);
output(1, 255) <= input(23);
output(2, 0) <= input(0);
output(2, 1) <= input(1);
output(2, 2) <= input(2);
output(2, 3) <= input(3);
output(2, 4) <= input(4);
output(2, 5) <= input(5);
output(2, 6) <= input(6);
output(2, 7) <= input(7);
output(2, 8) <= input(8);
output(2, 9) <= input(9);
output(2, 10) <= input(10);
output(2, 11) <= input(11);
output(2, 12) <= input(12);
output(2, 13) <= input(13);
output(2, 14) <= input(14);
output(2, 15) <= input(15);
output(2, 16) <= input(18);
output(2, 17) <= input(19);
output(2, 18) <= input(20);
output(2, 19) <= input(21);
output(2, 20) <= input(22);
output(2, 21) <= input(23);
output(2, 22) <= input(24);
output(2, 23) <= input(25);
output(2, 24) <= input(26);
output(2, 25) <= input(27);
output(2, 26) <= input(28);
output(2, 27) <= input(29);
output(2, 28) <= input(30);
output(2, 29) <= input(31);
output(2, 30) <= input(32);
output(2, 31) <= input(54);
output(2, 32) <= input(16);
output(2, 33) <= input(0);
output(2, 34) <= input(1);
output(2, 35) <= input(2);
output(2, 36) <= input(3);
output(2, 37) <= input(4);
output(2, 38) <= input(5);
output(2, 39) <= input(6);
output(2, 40) <= input(7);
output(2, 41) <= input(8);
output(2, 42) <= input(9);
output(2, 43) <= input(10);
output(2, 44) <= input(11);
output(2, 45) <= input(12);
output(2, 46) <= input(13);
output(2, 47) <= input(14);
output(2, 48) <= input(17);
output(2, 49) <= input(18);
output(2, 50) <= input(19);
output(2, 51) <= input(20);
output(2, 52) <= input(21);
output(2, 53) <= input(22);
output(2, 54) <= input(23);
output(2, 55) <= input(24);
output(2, 56) <= input(25);
output(2, 57) <= input(26);
output(2, 58) <= input(27);
output(2, 59) <= input(28);
output(2, 60) <= input(29);
output(2, 61) <= input(30);
output(2, 62) <= input(31);
output(2, 63) <= input(32);
output(2, 64) <= input(33);
output(2, 65) <= input(17);
output(2, 66) <= input(18);
output(2, 67) <= input(19);
output(2, 68) <= input(20);
output(2, 69) <= input(21);
output(2, 70) <= input(22);
output(2, 71) <= input(23);
output(2, 72) <= input(24);
output(2, 73) <= input(25);
output(2, 74) <= input(26);
output(2, 75) <= input(27);
output(2, 76) <= input(28);
output(2, 77) <= input(29);
output(2, 78) <= input(30);
output(2, 79) <= input(31);
output(2, 80) <= input(36);
output(2, 81) <= input(37);
output(2, 82) <= input(16);
output(2, 83) <= input(0);
output(2, 84) <= input(1);
output(2, 85) <= input(2);
output(2, 86) <= input(3);
output(2, 87) <= input(4);
output(2, 88) <= input(5);
output(2, 89) <= input(6);
output(2, 90) <= input(7);
output(2, 91) <= input(8);
output(2, 92) <= input(9);
output(2, 93) <= input(10);
output(2, 94) <= input(11);
output(2, 95) <= input(12);
output(2, 96) <= input(34);
output(2, 97) <= input(33);
output(2, 98) <= input(17);
output(2, 99) <= input(18);
output(2, 100) <= input(19);
output(2, 101) <= input(20);
output(2, 102) <= input(21);
output(2, 103) <= input(22);
output(2, 104) <= input(23);
output(2, 105) <= input(24);
output(2, 106) <= input(25);
output(2, 107) <= input(26);
output(2, 108) <= input(27);
output(2, 109) <= input(28);
output(2, 110) <= input(29);
output(2, 111) <= input(30);
output(2, 112) <= input(35);
output(2, 113) <= input(36);
output(2, 114) <= input(37);
output(2, 115) <= input(16);
output(2, 116) <= input(0);
output(2, 117) <= input(1);
output(2, 118) <= input(2);
output(2, 119) <= input(3);
output(2, 120) <= input(4);
output(2, 121) <= input(5);
output(2, 122) <= input(6);
output(2, 123) <= input(7);
output(2, 124) <= input(8);
output(2, 125) <= input(9);
output(2, 126) <= input(10);
output(2, 127) <= input(11);
output(2, 128) <= input(38);
output(2, 129) <= input(35);
output(2, 130) <= input(36);
output(2, 131) <= input(37);
output(2, 132) <= input(16);
output(2, 133) <= input(0);
output(2, 134) <= input(1);
output(2, 135) <= input(2);
output(2, 136) <= input(3);
output(2, 137) <= input(4);
output(2, 138) <= input(5);
output(2, 139) <= input(6);
output(2, 140) <= input(7);
output(2, 141) <= input(8);
output(2, 142) <= input(9);
output(2, 143) <= input(10);
output(2, 144) <= input(39);
output(2, 145) <= input(40);
output(2, 146) <= input(34);
output(2, 147) <= input(33);
output(2, 148) <= input(17);
output(2, 149) <= input(18);
output(2, 150) <= input(19);
output(2, 151) <= input(20);
output(2, 152) <= input(21);
output(2, 153) <= input(22);
output(2, 154) <= input(23);
output(2, 155) <= input(24);
output(2, 156) <= input(25);
output(2, 157) <= input(26);
output(2, 158) <= input(27);
output(2, 159) <= input(28);
output(2, 160) <= input(45);
output(2, 161) <= input(38);
output(2, 162) <= input(35);
output(2, 163) <= input(36);
output(2, 164) <= input(37);
output(2, 165) <= input(16);
output(2, 166) <= input(0);
output(2, 167) <= input(1);
output(2, 168) <= input(2);
output(2, 169) <= input(3);
output(2, 170) <= input(4);
output(2, 171) <= input(5);
output(2, 172) <= input(6);
output(2, 173) <= input(7);
output(2, 174) <= input(8);
output(2, 175) <= input(9);
output(2, 176) <= input(41);
output(2, 177) <= input(39);
output(2, 178) <= input(40);
output(2, 179) <= input(34);
output(2, 180) <= input(33);
output(2, 181) <= input(17);
output(2, 182) <= input(18);
output(2, 183) <= input(19);
output(2, 184) <= input(20);
output(2, 185) <= input(21);
output(2, 186) <= input(22);
output(2, 187) <= input(23);
output(2, 188) <= input(24);
output(2, 189) <= input(25);
output(2, 190) <= input(26);
output(2, 191) <= input(27);
output(2, 192) <= input(42);
output(2, 193) <= input(41);
output(2, 194) <= input(39);
output(2, 195) <= input(40);
output(2, 196) <= input(34);
output(2, 197) <= input(33);
output(2, 198) <= input(17);
output(2, 199) <= input(18);
output(2, 200) <= input(19);
output(2, 201) <= input(20);
output(2, 202) <= input(21);
output(2, 203) <= input(22);
output(2, 204) <= input(23);
output(2, 205) <= input(24);
output(2, 206) <= input(25);
output(2, 207) <= input(26);
output(2, 208) <= input(43);
output(2, 209) <= input(44);
output(2, 210) <= input(45);
output(2, 211) <= input(38);
output(2, 212) <= input(35);
output(2, 213) <= input(36);
output(2, 214) <= input(37);
output(2, 215) <= input(16);
output(2, 216) <= input(0);
output(2, 217) <= input(1);
output(2, 218) <= input(2);
output(2, 219) <= input(3);
output(2, 220) <= input(4);
output(2, 221) <= input(5);
output(2, 222) <= input(6);
output(2, 223) <= input(7);
output(2, 224) <= input(50);
output(2, 225) <= input(42);
output(2, 226) <= input(41);
output(2, 227) <= input(39);
output(2, 228) <= input(40);
output(2, 229) <= input(34);
output(2, 230) <= input(33);
output(2, 231) <= input(17);
output(2, 232) <= input(18);
output(2, 233) <= input(19);
output(2, 234) <= input(20);
output(2, 235) <= input(21);
output(2, 236) <= input(22);
output(2, 237) <= input(23);
output(2, 238) <= input(24);
output(2, 239) <= input(25);
output(2, 240) <= input(46);
output(2, 241) <= input(43);
output(2, 242) <= input(44);
output(2, 243) <= input(45);
output(2, 244) <= input(38);
output(2, 245) <= input(35);
output(2, 246) <= input(36);
output(2, 247) <= input(37);
output(2, 248) <= input(16);
output(2, 249) <= input(0);
output(2, 250) <= input(1);
output(2, 251) <= input(2);
output(2, 252) <= input(3);
output(2, 253) <= input(4);
output(2, 254) <= input(5);
output(2, 255) <= input(6);
when "1010" =>
output(0, 0) <= input(0);
output(0, 1) <= input(1);
output(0, 2) <= input(2);
output(0, 3) <= input(3);
output(0, 4) <= input(4);
output(0, 5) <= input(5);
output(0, 6) <= input(6);
output(0, 7) <= input(7);
output(0, 8) <= input(8);
output(0, 9) <= input(9);
output(0, 10) <= input(10);
output(0, 11) <= input(11);
output(0, 12) <= input(12);
output(0, 13) <= input(13);
output(0, 14) <= input(14);
output(0, 15) <= input(15);
output(0, 16) <= input(16);
output(0, 17) <= input(17);
output(0, 18) <= input(18);
output(0, 19) <= input(19);
output(0, 20) <= input(20);
output(0, 21) <= input(21);
output(0, 22) <= input(22);
output(0, 23) <= input(23);
output(0, 24) <= input(24);
output(0, 25) <= input(25);
output(0, 26) <= input(26);
output(0, 27) <= input(27);
output(0, 28) <= input(28);
output(0, 29) <= input(29);
output(0, 30) <= input(30);
output(0, 31) <= input(31);
output(0, 32) <= input(32);
output(0, 33) <= input(0);
output(0, 34) <= input(1);
output(0, 35) <= input(2);
output(0, 36) <= input(3);
output(0, 37) <= input(4);
output(0, 38) <= input(5);
output(0, 39) <= input(6);
output(0, 40) <= input(7);
output(0, 41) <= input(8);
output(0, 42) <= input(9);
output(0, 43) <= input(10);
output(0, 44) <= input(11);
output(0, 45) <= input(12);
output(0, 46) <= input(13);
output(0, 47) <= input(14);
output(0, 48) <= input(33);
output(0, 49) <= input(16);
output(0, 50) <= input(17);
output(0, 51) <= input(18);
output(0, 52) <= input(19);
output(0, 53) <= input(20);
output(0, 54) <= input(21);
output(0, 55) <= input(22);
output(0, 56) <= input(23);
output(0, 57) <= input(24);
output(0, 58) <= input(25);
output(0, 59) <= input(26);
output(0, 60) <= input(27);
output(0, 61) <= input(28);
output(0, 62) <= input(29);
output(0, 63) <= input(30);
output(0, 64) <= input(34);
output(0, 65) <= input(32);
output(0, 66) <= input(0);
output(0, 67) <= input(1);
output(0, 68) <= input(2);
output(0, 69) <= input(3);
output(0, 70) <= input(4);
output(0, 71) <= input(5);
output(0, 72) <= input(6);
output(0, 73) <= input(7);
output(0, 74) <= input(8);
output(0, 75) <= input(9);
output(0, 76) <= input(10);
output(0, 77) <= input(11);
output(0, 78) <= input(12);
output(0, 79) <= input(13);
output(0, 80) <= input(35);
output(0, 81) <= input(33);
output(0, 82) <= input(16);
output(0, 83) <= input(17);
output(0, 84) <= input(18);
output(0, 85) <= input(19);
output(0, 86) <= input(20);
output(0, 87) <= input(21);
output(0, 88) <= input(22);
output(0, 89) <= input(23);
output(0, 90) <= input(24);
output(0, 91) <= input(25);
output(0, 92) <= input(26);
output(0, 93) <= input(27);
output(0, 94) <= input(28);
output(0, 95) <= input(29);
output(0, 96) <= input(36);
output(0, 97) <= input(34);
output(0, 98) <= input(32);
output(0, 99) <= input(0);
output(0, 100) <= input(1);
output(0, 101) <= input(2);
output(0, 102) <= input(3);
output(0, 103) <= input(4);
output(0, 104) <= input(5);
output(0, 105) <= input(6);
output(0, 106) <= input(7);
output(0, 107) <= input(8);
output(0, 108) <= input(9);
output(0, 109) <= input(10);
output(0, 110) <= input(11);
output(0, 111) <= input(12);
output(0, 112) <= input(37);
output(0, 113) <= input(35);
output(0, 114) <= input(33);
output(0, 115) <= input(16);
output(0, 116) <= input(17);
output(0, 117) <= input(18);
output(0, 118) <= input(19);
output(0, 119) <= input(20);
output(0, 120) <= input(21);
output(0, 121) <= input(22);
output(0, 122) <= input(23);
output(0, 123) <= input(24);
output(0, 124) <= input(25);
output(0, 125) <= input(26);
output(0, 126) <= input(27);
output(0, 127) <= input(28);
output(0, 128) <= input(38);
output(0, 129) <= input(37);
output(0, 130) <= input(35);
output(0, 131) <= input(33);
output(0, 132) <= input(16);
output(0, 133) <= input(17);
output(0, 134) <= input(18);
output(0, 135) <= input(19);
output(0, 136) <= input(20);
output(0, 137) <= input(21);
output(0, 138) <= input(22);
output(0, 139) <= input(23);
output(0, 140) <= input(24);
output(0, 141) <= input(25);
output(0, 142) <= input(26);
output(0, 143) <= input(27);
output(0, 144) <= input(39);
output(0, 145) <= input(40);
output(0, 146) <= input(36);
output(0, 147) <= input(34);
output(0, 148) <= input(32);
output(0, 149) <= input(0);
output(0, 150) <= input(1);
output(0, 151) <= input(2);
output(0, 152) <= input(3);
output(0, 153) <= input(4);
output(0, 154) <= input(5);
output(0, 155) <= input(6);
output(0, 156) <= input(7);
output(0, 157) <= input(8);
output(0, 158) <= input(9);
output(0, 159) <= input(10);
output(0, 160) <= input(41);
output(0, 161) <= input(38);
output(0, 162) <= input(37);
output(0, 163) <= input(35);
output(0, 164) <= input(33);
output(0, 165) <= input(16);
output(0, 166) <= input(17);
output(0, 167) <= input(18);
output(0, 168) <= input(19);
output(0, 169) <= input(20);
output(0, 170) <= input(21);
output(0, 171) <= input(22);
output(0, 172) <= input(23);
output(0, 173) <= input(24);
output(0, 174) <= input(25);
output(0, 175) <= input(26);
output(0, 176) <= input(42);
output(0, 177) <= input(39);
output(0, 178) <= input(40);
output(0, 179) <= input(36);
output(0, 180) <= input(34);
output(0, 181) <= input(32);
output(0, 182) <= input(0);
output(0, 183) <= input(1);
output(0, 184) <= input(2);
output(0, 185) <= input(3);
output(0, 186) <= input(4);
output(0, 187) <= input(5);
output(0, 188) <= input(6);
output(0, 189) <= input(7);
output(0, 190) <= input(8);
output(0, 191) <= input(9);
output(0, 192) <= input(43);
output(0, 193) <= input(41);
output(0, 194) <= input(38);
output(0, 195) <= input(37);
output(0, 196) <= input(35);
output(0, 197) <= input(33);
output(0, 198) <= input(16);
output(0, 199) <= input(17);
output(0, 200) <= input(18);
output(0, 201) <= input(19);
output(0, 202) <= input(20);
output(0, 203) <= input(21);
output(0, 204) <= input(22);
output(0, 205) <= input(23);
output(0, 206) <= input(24);
output(0, 207) <= input(25);
output(0, 208) <= input(44);
output(0, 209) <= input(42);
output(0, 210) <= input(39);
output(0, 211) <= input(40);
output(0, 212) <= input(36);
output(0, 213) <= input(34);
output(0, 214) <= input(32);
output(0, 215) <= input(0);
output(0, 216) <= input(1);
output(0, 217) <= input(2);
output(0, 218) <= input(3);
output(0, 219) <= input(4);
output(0, 220) <= input(5);
output(0, 221) <= input(6);
output(0, 222) <= input(7);
output(0, 223) <= input(8);
output(0, 224) <= input(45);
output(0, 225) <= input(43);
output(0, 226) <= input(41);
output(0, 227) <= input(38);
output(0, 228) <= input(37);
output(0, 229) <= input(35);
output(0, 230) <= input(33);
output(0, 231) <= input(16);
output(0, 232) <= input(17);
output(0, 233) <= input(18);
output(0, 234) <= input(19);
output(0, 235) <= input(20);
output(0, 236) <= input(21);
output(0, 237) <= input(22);
output(0, 238) <= input(23);
output(0, 239) <= input(24);
output(0, 240) <= input(46);
output(0, 241) <= input(44);
output(0, 242) <= input(42);
output(0, 243) <= input(39);
output(0, 244) <= input(40);
output(0, 245) <= input(36);
output(0, 246) <= input(34);
output(0, 247) <= input(32);
output(0, 248) <= input(0);
output(0, 249) <= input(1);
output(0, 250) <= input(2);
output(0, 251) <= input(3);
output(0, 252) <= input(4);
output(0, 253) <= input(5);
output(0, 254) <= input(6);
output(0, 255) <= input(7);
output(1, 0) <= input(17);
output(1, 1) <= input(18);
output(1, 2) <= input(19);
output(1, 3) <= input(20);
output(1, 4) <= input(21);
output(1, 5) <= input(22);
output(1, 6) <= input(23);
output(1, 7) <= input(24);
output(1, 8) <= input(25);
output(1, 9) <= input(26);
output(1, 10) <= input(27);
output(1, 11) <= input(28);
output(1, 12) <= input(29);
output(1, 13) <= input(30);
output(1, 14) <= input(31);
output(1, 15) <= input(47);
output(1, 16) <= input(0);
output(1, 17) <= input(1);
output(1, 18) <= input(2);
output(1, 19) <= input(3);
output(1, 20) <= input(4);
output(1, 21) <= input(5);
output(1, 22) <= input(6);
output(1, 23) <= input(7);
output(1, 24) <= input(8);
output(1, 25) <= input(9);
output(1, 26) <= input(10);
output(1, 27) <= input(11);
output(1, 28) <= input(12);
output(1, 29) <= input(13);
output(1, 30) <= input(14);
output(1, 31) <= input(15);
output(1, 32) <= input(16);
output(1, 33) <= input(17);
output(1, 34) <= input(18);
output(1, 35) <= input(19);
output(1, 36) <= input(20);
output(1, 37) <= input(21);
output(1, 38) <= input(22);
output(1, 39) <= input(23);
output(1, 40) <= input(24);
output(1, 41) <= input(25);
output(1, 42) <= input(26);
output(1, 43) <= input(27);
output(1, 44) <= input(28);
output(1, 45) <= input(29);
output(1, 46) <= input(30);
output(1, 47) <= input(31);
output(1, 48) <= input(32);
output(1, 49) <= input(0);
output(1, 50) <= input(1);
output(1, 51) <= input(2);
output(1, 52) <= input(3);
output(1, 53) <= input(4);
output(1, 54) <= input(5);
output(1, 55) <= input(6);
output(1, 56) <= input(7);
output(1, 57) <= input(8);
output(1, 58) <= input(9);
output(1, 59) <= input(10);
output(1, 60) <= input(11);
output(1, 61) <= input(12);
output(1, 62) <= input(13);
output(1, 63) <= input(14);
output(1, 64) <= input(33);
output(1, 65) <= input(16);
output(1, 66) <= input(17);
output(1, 67) <= input(18);
output(1, 68) <= input(19);
output(1, 69) <= input(20);
output(1, 70) <= input(21);
output(1, 71) <= input(22);
output(1, 72) <= input(23);
output(1, 73) <= input(24);
output(1, 74) <= input(25);
output(1, 75) <= input(26);
output(1, 76) <= input(27);
output(1, 77) <= input(28);
output(1, 78) <= input(29);
output(1, 79) <= input(30);
output(1, 80) <= input(34);
output(1, 81) <= input(32);
output(1, 82) <= input(0);
output(1, 83) <= input(1);
output(1, 84) <= input(2);
output(1, 85) <= input(3);
output(1, 86) <= input(4);
output(1, 87) <= input(5);
output(1, 88) <= input(6);
output(1, 89) <= input(7);
output(1, 90) <= input(8);
output(1, 91) <= input(9);
output(1, 92) <= input(10);
output(1, 93) <= input(11);
output(1, 94) <= input(12);
output(1, 95) <= input(13);
output(1, 96) <= input(35);
output(1, 97) <= input(33);
output(1, 98) <= input(16);
output(1, 99) <= input(17);
output(1, 100) <= input(18);
output(1, 101) <= input(19);
output(1, 102) <= input(20);
output(1, 103) <= input(21);
output(1, 104) <= input(22);
output(1, 105) <= input(23);
output(1, 106) <= input(24);
output(1, 107) <= input(25);
output(1, 108) <= input(26);
output(1, 109) <= input(27);
output(1, 110) <= input(28);
output(1, 111) <= input(29);
output(1, 112) <= input(36);
output(1, 113) <= input(34);
output(1, 114) <= input(32);
output(1, 115) <= input(0);
output(1, 116) <= input(1);
output(1, 117) <= input(2);
output(1, 118) <= input(3);
output(1, 119) <= input(4);
output(1, 120) <= input(5);
output(1, 121) <= input(6);
output(1, 122) <= input(7);
output(1, 123) <= input(8);
output(1, 124) <= input(9);
output(1, 125) <= input(10);
output(1, 126) <= input(11);
output(1, 127) <= input(12);
output(1, 128) <= input(37);
output(1, 129) <= input(35);
output(1, 130) <= input(33);
output(1, 131) <= input(16);
output(1, 132) <= input(17);
output(1, 133) <= input(18);
output(1, 134) <= input(19);
output(1, 135) <= input(20);
output(1, 136) <= input(21);
output(1, 137) <= input(22);
output(1, 138) <= input(23);
output(1, 139) <= input(24);
output(1, 140) <= input(25);
output(1, 141) <= input(26);
output(1, 142) <= input(27);
output(1, 143) <= input(28);
output(1, 144) <= input(40);
output(1, 145) <= input(36);
output(1, 146) <= input(34);
output(1, 147) <= input(32);
output(1, 148) <= input(0);
output(1, 149) <= input(1);
output(1, 150) <= input(2);
output(1, 151) <= input(3);
output(1, 152) <= input(4);
output(1, 153) <= input(5);
output(1, 154) <= input(6);
output(1, 155) <= input(7);
output(1, 156) <= input(8);
output(1, 157) <= input(9);
output(1, 158) <= input(10);
output(1, 159) <= input(11);
output(1, 160) <= input(38);
output(1, 161) <= input(37);
output(1, 162) <= input(35);
output(1, 163) <= input(33);
output(1, 164) <= input(16);
output(1, 165) <= input(17);
output(1, 166) <= input(18);
output(1, 167) <= input(19);
output(1, 168) <= input(20);
output(1, 169) <= input(21);
output(1, 170) <= input(22);
output(1, 171) <= input(23);
output(1, 172) <= input(24);
output(1, 173) <= input(25);
output(1, 174) <= input(26);
output(1, 175) <= input(27);
output(1, 176) <= input(39);
output(1, 177) <= input(40);
output(1, 178) <= input(36);
output(1, 179) <= input(34);
output(1, 180) <= input(32);
output(1, 181) <= input(0);
output(1, 182) <= input(1);
output(1, 183) <= input(2);
output(1, 184) <= input(3);
output(1, 185) <= input(4);
output(1, 186) <= input(5);
output(1, 187) <= input(6);
output(1, 188) <= input(7);
output(1, 189) <= input(8);
output(1, 190) <= input(9);
output(1, 191) <= input(10);
output(1, 192) <= input(41);
output(1, 193) <= input(38);
output(1, 194) <= input(37);
output(1, 195) <= input(35);
output(1, 196) <= input(33);
output(1, 197) <= input(16);
output(1, 198) <= input(17);
output(1, 199) <= input(18);
output(1, 200) <= input(19);
output(1, 201) <= input(20);
output(1, 202) <= input(21);
output(1, 203) <= input(22);
output(1, 204) <= input(23);
output(1, 205) <= input(24);
output(1, 206) <= input(25);
output(1, 207) <= input(26);
output(1, 208) <= input(42);
output(1, 209) <= input(39);
output(1, 210) <= input(40);
output(1, 211) <= input(36);
output(1, 212) <= input(34);
output(1, 213) <= input(32);
output(1, 214) <= input(0);
output(1, 215) <= input(1);
output(1, 216) <= input(2);
output(1, 217) <= input(3);
output(1, 218) <= input(4);
output(1, 219) <= input(5);
output(1, 220) <= input(6);
output(1, 221) <= input(7);
output(1, 222) <= input(8);
output(1, 223) <= input(9);
output(1, 224) <= input(43);
output(1, 225) <= input(41);
output(1, 226) <= input(38);
output(1, 227) <= input(37);
output(1, 228) <= input(35);
output(1, 229) <= input(33);
output(1, 230) <= input(16);
output(1, 231) <= input(17);
output(1, 232) <= input(18);
output(1, 233) <= input(19);
output(1, 234) <= input(20);
output(1, 235) <= input(21);
output(1, 236) <= input(22);
output(1, 237) <= input(23);
output(1, 238) <= input(24);
output(1, 239) <= input(25);
output(1, 240) <= input(44);
output(1, 241) <= input(42);
output(1, 242) <= input(39);
output(1, 243) <= input(40);
output(1, 244) <= input(36);
output(1, 245) <= input(34);
output(1, 246) <= input(32);
output(1, 247) <= input(0);
output(1, 248) <= input(1);
output(1, 249) <= input(2);
output(1, 250) <= input(3);
output(1, 251) <= input(4);
output(1, 252) <= input(5);
output(1, 253) <= input(6);
output(1, 254) <= input(7);
output(1, 255) <= input(8);
when "1011" =>
output(0, 0) <= input(0);
output(0, 1) <= input(1);
output(0, 2) <= input(2);
output(0, 3) <= input(3);
output(0, 4) <= input(4);
output(0, 5) <= input(5);
output(0, 6) <= input(6);
output(0, 7) <= input(7);
output(0, 8) <= input(8);
output(0, 9) <= input(9);
output(0, 10) <= input(10);
output(0, 11) <= input(11);
output(0, 12) <= input(12);
output(0, 13) <= input(13);
output(0, 14) <= input(14);
output(0, 15) <= input(15);
output(0, 16) <= input(16);
output(0, 17) <= input(17);
output(0, 18) <= input(18);
output(0, 19) <= input(19);
output(0, 20) <= input(20);
output(0, 21) <= input(21);
output(0, 22) <= input(22);
output(0, 23) <= input(23);
output(0, 24) <= input(24);
output(0, 25) <= input(25);
output(0, 26) <= input(26);
output(0, 27) <= input(27);
output(0, 28) <= input(28);
output(0, 29) <= input(29);
output(0, 30) <= input(30);
output(0, 31) <= input(31);
output(0, 32) <= input(32);
output(0, 33) <= input(0);
output(0, 34) <= input(1);
output(0, 35) <= input(2);
output(0, 36) <= input(3);
output(0, 37) <= input(4);
output(0, 38) <= input(5);
output(0, 39) <= input(6);
output(0, 40) <= input(7);
output(0, 41) <= input(8);
output(0, 42) <= input(9);
output(0, 43) <= input(10);
output(0, 44) <= input(11);
output(0, 45) <= input(12);
output(0, 46) <= input(13);
output(0, 47) <= input(14);
output(0, 48) <= input(33);
output(0, 49) <= input(16);
output(0, 50) <= input(17);
output(0, 51) <= input(18);
output(0, 52) <= input(19);
output(0, 53) <= input(20);
output(0, 54) <= input(21);
output(0, 55) <= input(22);
output(0, 56) <= input(23);
output(0, 57) <= input(24);
output(0, 58) <= input(25);
output(0, 59) <= input(26);
output(0, 60) <= input(27);
output(0, 61) <= input(28);
output(0, 62) <= input(29);
output(0, 63) <= input(30);
output(0, 64) <= input(34);
output(0, 65) <= input(32);
output(0, 66) <= input(0);
output(0, 67) <= input(1);
output(0, 68) <= input(2);
output(0, 69) <= input(3);
output(0, 70) <= input(4);
output(0, 71) <= input(5);
output(0, 72) <= input(6);
output(0, 73) <= input(7);
output(0, 74) <= input(8);
output(0, 75) <= input(9);
output(0, 76) <= input(10);
output(0, 77) <= input(11);
output(0, 78) <= input(12);
output(0, 79) <= input(13);
output(0, 80) <= input(35);
output(0, 81) <= input(33);
output(0, 82) <= input(16);
output(0, 83) <= input(17);
output(0, 84) <= input(18);
output(0, 85) <= input(19);
output(0, 86) <= input(20);
output(0, 87) <= input(21);
output(0, 88) <= input(22);
output(0, 89) <= input(23);
output(0, 90) <= input(24);
output(0, 91) <= input(25);
output(0, 92) <= input(26);
output(0, 93) <= input(27);
output(0, 94) <= input(28);
output(0, 95) <= input(29);
output(0, 96) <= input(36);
output(0, 97) <= input(34);
output(0, 98) <= input(32);
output(0, 99) <= input(0);
output(0, 100) <= input(1);
output(0, 101) <= input(2);
output(0, 102) <= input(3);
output(0, 103) <= input(4);
output(0, 104) <= input(5);
output(0, 105) <= input(6);
output(0, 106) <= input(7);
output(0, 107) <= input(8);
output(0, 108) <= input(9);
output(0, 109) <= input(10);
output(0, 110) <= input(11);
output(0, 111) <= input(12);
output(0, 112) <= input(36);
output(0, 113) <= input(34);
output(0, 114) <= input(32);
output(0, 115) <= input(0);
output(0, 116) <= input(1);
output(0, 117) <= input(2);
output(0, 118) <= input(3);
output(0, 119) <= input(4);
output(0, 120) <= input(5);
output(0, 121) <= input(6);
output(0, 122) <= input(7);
output(0, 123) <= input(8);
output(0, 124) <= input(9);
output(0, 125) <= input(10);
output(0, 126) <= input(11);
output(0, 127) <= input(12);
output(0, 128) <= input(37);
output(0, 129) <= input(35);
output(0, 130) <= input(33);
output(0, 131) <= input(16);
output(0, 132) <= input(17);
output(0, 133) <= input(18);
output(0, 134) <= input(19);
output(0, 135) <= input(20);
output(0, 136) <= input(21);
output(0, 137) <= input(22);
output(0, 138) <= input(23);
output(0, 139) <= input(24);
output(0, 140) <= input(25);
output(0, 141) <= input(26);
output(0, 142) <= input(27);
output(0, 143) <= input(28);
output(0, 144) <= input(38);
output(0, 145) <= input(36);
output(0, 146) <= input(34);
output(0, 147) <= input(32);
output(0, 148) <= input(0);
output(0, 149) <= input(1);
output(0, 150) <= input(2);
output(0, 151) <= input(3);
output(0, 152) <= input(4);
output(0, 153) <= input(5);
output(0, 154) <= input(6);
output(0, 155) <= input(7);
output(0, 156) <= input(8);
output(0, 157) <= input(9);
output(0, 158) <= input(10);
output(0, 159) <= input(11);
output(0, 160) <= input(39);
output(0, 161) <= input(37);
output(0, 162) <= input(35);
output(0, 163) <= input(33);
output(0, 164) <= input(16);
output(0, 165) <= input(17);
output(0, 166) <= input(18);
output(0, 167) <= input(19);
output(0, 168) <= input(20);
output(0, 169) <= input(21);
output(0, 170) <= input(22);
output(0, 171) <= input(23);
output(0, 172) <= input(24);
output(0, 173) <= input(25);
output(0, 174) <= input(26);
output(0, 175) <= input(27);
output(0, 176) <= input(40);
output(0, 177) <= input(38);
output(0, 178) <= input(36);
output(0, 179) <= input(34);
output(0, 180) <= input(32);
output(0, 181) <= input(0);
output(0, 182) <= input(1);
output(0, 183) <= input(2);
output(0, 184) <= input(3);
output(0, 185) <= input(4);
output(0, 186) <= input(5);
output(0, 187) <= input(6);
output(0, 188) <= input(7);
output(0, 189) <= input(8);
output(0, 190) <= input(9);
output(0, 191) <= input(10);
output(0, 192) <= input(41);
output(0, 193) <= input(39);
output(0, 194) <= input(37);
output(0, 195) <= input(35);
output(0, 196) <= input(33);
output(0, 197) <= input(16);
output(0, 198) <= input(17);
output(0, 199) <= input(18);
output(0, 200) <= input(19);
output(0, 201) <= input(20);
output(0, 202) <= input(21);
output(0, 203) <= input(22);
output(0, 204) <= input(23);
output(0, 205) <= input(24);
output(0, 206) <= input(25);
output(0, 207) <= input(26);
output(0, 208) <= input(42);
output(0, 209) <= input(40);
output(0, 210) <= input(38);
output(0, 211) <= input(36);
output(0, 212) <= input(34);
output(0, 213) <= input(32);
output(0, 214) <= input(0);
output(0, 215) <= input(1);
output(0, 216) <= input(2);
output(0, 217) <= input(3);
output(0, 218) <= input(4);
output(0, 219) <= input(5);
output(0, 220) <= input(6);
output(0, 221) <= input(7);
output(0, 222) <= input(8);
output(0, 223) <= input(9);
output(0, 224) <= input(43);
output(0, 225) <= input(41);
output(0, 226) <= input(39);
output(0, 227) <= input(37);
output(0, 228) <= input(35);
output(0, 229) <= input(33);
output(0, 230) <= input(16);
output(0, 231) <= input(17);
output(0, 232) <= input(18);
output(0, 233) <= input(19);
output(0, 234) <= input(20);
output(0, 235) <= input(21);
output(0, 236) <= input(22);
output(0, 237) <= input(23);
output(0, 238) <= input(24);
output(0, 239) <= input(25);
output(0, 240) <= input(43);
output(0, 241) <= input(41);
output(0, 242) <= input(39);
output(0, 243) <= input(37);
output(0, 244) <= input(35);
output(0, 245) <= input(33);
output(0, 246) <= input(16);
output(0, 247) <= input(17);
output(0, 248) <= input(18);
output(0, 249) <= input(19);
output(0, 250) <= input(20);
output(0, 251) <= input(21);
output(0, 252) <= input(22);
output(0, 253) <= input(23);
output(0, 254) <= input(24);
output(0, 255) <= input(25);
output(1, 0) <= input(0);
output(1, 1) <= input(1);
output(1, 2) <= input(2);
output(1, 3) <= input(3);
output(1, 4) <= input(4);
output(1, 5) <= input(5);
output(1, 6) <= input(6);
output(1, 7) <= input(7);
output(1, 8) <= input(8);
output(1, 9) <= input(9);
output(1, 10) <= input(10);
output(1, 11) <= input(11);
output(1, 12) <= input(12);
output(1, 13) <= input(13);
output(1, 14) <= input(14);
output(1, 15) <= input(15);
output(1, 16) <= input(16);
output(1, 17) <= input(17);
output(1, 18) <= input(18);
output(1, 19) <= input(19);
output(1, 20) <= input(20);
output(1, 21) <= input(21);
output(1, 22) <= input(22);
output(1, 23) <= input(23);
output(1, 24) <= input(24);
output(1, 25) <= input(25);
output(1, 26) <= input(26);
output(1, 27) <= input(27);
output(1, 28) <= input(28);
output(1, 29) <= input(29);
output(1, 30) <= input(30);
output(1, 31) <= input(31);
output(1, 32) <= input(32);
output(1, 33) <= input(0);
output(1, 34) <= input(1);
output(1, 35) <= input(2);
output(1, 36) <= input(3);
output(1, 37) <= input(4);
output(1, 38) <= input(5);
output(1, 39) <= input(6);
output(1, 40) <= input(7);
output(1, 41) <= input(8);
output(1, 42) <= input(9);
output(1, 43) <= input(10);
output(1, 44) <= input(11);
output(1, 45) <= input(12);
output(1, 46) <= input(13);
output(1, 47) <= input(14);
output(1, 48) <= input(32);
output(1, 49) <= input(0);
output(1, 50) <= input(1);
output(1, 51) <= input(2);
output(1, 52) <= input(3);
output(1, 53) <= input(4);
output(1, 54) <= input(5);
output(1, 55) <= input(6);
output(1, 56) <= input(7);
output(1, 57) <= input(8);
output(1, 58) <= input(9);
output(1, 59) <= input(10);
output(1, 60) <= input(11);
output(1, 61) <= input(12);
output(1, 62) <= input(13);
output(1, 63) <= input(14);
output(1, 64) <= input(33);
output(1, 65) <= input(16);
output(1, 66) <= input(17);
output(1, 67) <= input(18);
output(1, 68) <= input(19);
output(1, 69) <= input(20);
output(1, 70) <= input(21);
output(1, 71) <= input(22);
output(1, 72) <= input(23);
output(1, 73) <= input(24);
output(1, 74) <= input(25);
output(1, 75) <= input(26);
output(1, 76) <= input(27);
output(1, 77) <= input(28);
output(1, 78) <= input(29);
output(1, 79) <= input(30);
output(1, 80) <= input(34);
output(1, 81) <= input(32);
output(1, 82) <= input(0);
output(1, 83) <= input(1);
output(1, 84) <= input(2);
output(1, 85) <= input(3);
output(1, 86) <= input(4);
output(1, 87) <= input(5);
output(1, 88) <= input(6);
output(1, 89) <= input(7);
output(1, 90) <= input(8);
output(1, 91) <= input(9);
output(1, 92) <= input(10);
output(1, 93) <= input(11);
output(1, 94) <= input(12);
output(1, 95) <= input(13);
output(1, 96) <= input(35);
output(1, 97) <= input(33);
output(1, 98) <= input(16);
output(1, 99) <= input(17);
output(1, 100) <= input(18);
output(1, 101) <= input(19);
output(1, 102) <= input(20);
output(1, 103) <= input(21);
output(1, 104) <= input(22);
output(1, 105) <= input(23);
output(1, 106) <= input(24);
output(1, 107) <= input(25);
output(1, 108) <= input(26);
output(1, 109) <= input(27);
output(1, 110) <= input(28);
output(1, 111) <= input(29);
output(1, 112) <= input(35);
output(1, 113) <= input(33);
output(1, 114) <= input(16);
output(1, 115) <= input(17);
output(1, 116) <= input(18);
output(1, 117) <= input(19);
output(1, 118) <= input(20);
output(1, 119) <= input(21);
output(1, 120) <= input(22);
output(1, 121) <= input(23);
output(1, 122) <= input(24);
output(1, 123) <= input(25);
output(1, 124) <= input(26);
output(1, 125) <= input(27);
output(1, 126) <= input(28);
output(1, 127) <= input(29);
output(1, 128) <= input(36);
output(1, 129) <= input(34);
output(1, 130) <= input(32);
output(1, 131) <= input(0);
output(1, 132) <= input(1);
output(1, 133) <= input(2);
output(1, 134) <= input(3);
output(1, 135) <= input(4);
output(1, 136) <= input(5);
output(1, 137) <= input(6);
output(1, 138) <= input(7);
output(1, 139) <= input(8);
output(1, 140) <= input(9);
output(1, 141) <= input(10);
output(1, 142) <= input(11);
output(1, 143) <= input(12);
output(1, 144) <= input(37);
output(1, 145) <= input(35);
output(1, 146) <= input(33);
output(1, 147) <= input(16);
output(1, 148) <= input(17);
output(1, 149) <= input(18);
output(1, 150) <= input(19);
output(1, 151) <= input(20);
output(1, 152) <= input(21);
output(1, 153) <= input(22);
output(1, 154) <= input(23);
output(1, 155) <= input(24);
output(1, 156) <= input(25);
output(1, 157) <= input(26);
output(1, 158) <= input(27);
output(1, 159) <= input(28);
output(1, 160) <= input(38);
output(1, 161) <= input(36);
output(1, 162) <= input(34);
output(1, 163) <= input(32);
output(1, 164) <= input(0);
output(1, 165) <= input(1);
output(1, 166) <= input(2);
output(1, 167) <= input(3);
output(1, 168) <= input(4);
output(1, 169) <= input(5);
output(1, 170) <= input(6);
output(1, 171) <= input(7);
output(1, 172) <= input(8);
output(1, 173) <= input(9);
output(1, 174) <= input(10);
output(1, 175) <= input(11);
output(1, 176) <= input(38);
output(1, 177) <= input(36);
output(1, 178) <= input(34);
output(1, 179) <= input(32);
output(1, 180) <= input(0);
output(1, 181) <= input(1);
output(1, 182) <= input(2);
output(1, 183) <= input(3);
output(1, 184) <= input(4);
output(1, 185) <= input(5);
output(1, 186) <= input(6);
output(1, 187) <= input(7);
output(1, 188) <= input(8);
output(1, 189) <= input(9);
output(1, 190) <= input(10);
output(1, 191) <= input(11);
output(1, 192) <= input(39);
output(1, 193) <= input(37);
output(1, 194) <= input(35);
output(1, 195) <= input(33);
output(1, 196) <= input(16);
output(1, 197) <= input(17);
output(1, 198) <= input(18);
output(1, 199) <= input(19);
output(1, 200) <= input(20);
output(1, 201) <= input(21);
output(1, 202) <= input(22);
output(1, 203) <= input(23);
output(1, 204) <= input(24);
output(1, 205) <= input(25);
output(1, 206) <= input(26);
output(1, 207) <= input(27);
output(1, 208) <= input(40);
output(1, 209) <= input(38);
output(1, 210) <= input(36);
output(1, 211) <= input(34);
output(1, 212) <= input(32);
output(1, 213) <= input(0);
output(1, 214) <= input(1);
output(1, 215) <= input(2);
output(1, 216) <= input(3);
output(1, 217) <= input(4);
output(1, 218) <= input(5);
output(1, 219) <= input(6);
output(1, 220) <= input(7);
output(1, 221) <= input(8);
output(1, 222) <= input(9);
output(1, 223) <= input(10);
output(1, 224) <= input(41);
output(1, 225) <= input(39);
output(1, 226) <= input(37);
output(1, 227) <= input(35);
output(1, 228) <= input(33);
output(1, 229) <= input(16);
output(1, 230) <= input(17);
output(1, 231) <= input(18);
output(1, 232) <= input(19);
output(1, 233) <= input(20);
output(1, 234) <= input(21);
output(1, 235) <= input(22);
output(1, 236) <= input(23);
output(1, 237) <= input(24);
output(1, 238) <= input(25);
output(1, 239) <= input(26);
output(1, 240) <= input(41);
output(1, 241) <= input(39);
output(1, 242) <= input(37);
output(1, 243) <= input(35);
output(1, 244) <= input(33);
output(1, 245) <= input(16);
output(1, 246) <= input(17);
output(1, 247) <= input(18);
output(1, 248) <= input(19);
output(1, 249) <= input(20);
output(1, 250) <= input(21);
output(1, 251) <= input(22);
output(1, 252) <= input(23);
output(1, 253) <= input(24);
output(1, 254) <= input(25);
output(1, 255) <= input(26);
output(2, 0) <= input(0);
output(2, 1) <= input(1);
output(2, 2) <= input(2);
output(2, 3) <= input(3);
output(2, 4) <= input(4);
output(2, 5) <= input(5);
output(2, 6) <= input(6);
output(2, 7) <= input(7);
output(2, 8) <= input(8);
output(2, 9) <= input(9);
output(2, 10) <= input(10);
output(2, 11) <= input(11);
output(2, 12) <= input(12);
output(2, 13) <= input(13);
output(2, 14) <= input(14);
output(2, 15) <= input(15);
output(2, 16) <= input(16);
output(2, 17) <= input(17);
output(2, 18) <= input(18);
output(2, 19) <= input(19);
output(2, 20) <= input(20);
output(2, 21) <= input(21);
output(2, 22) <= input(22);
output(2, 23) <= input(23);
output(2, 24) <= input(24);
output(2, 25) <= input(25);
output(2, 26) <= input(26);
output(2, 27) <= input(27);
output(2, 28) <= input(28);
output(2, 29) <= input(29);
output(2, 30) <= input(30);
output(2, 31) <= input(31);
output(2, 32) <= input(16);
output(2, 33) <= input(17);
output(2, 34) <= input(18);
output(2, 35) <= input(19);
output(2, 36) <= input(20);
output(2, 37) <= input(21);
output(2, 38) <= input(22);
output(2, 39) <= input(23);
output(2, 40) <= input(24);
output(2, 41) <= input(25);
output(2, 42) <= input(26);
output(2, 43) <= input(27);
output(2, 44) <= input(28);
output(2, 45) <= input(29);
output(2, 46) <= input(30);
output(2, 47) <= input(31);
output(2, 48) <= input(32);
output(2, 49) <= input(0);
output(2, 50) <= input(1);
output(2, 51) <= input(2);
output(2, 52) <= input(3);
output(2, 53) <= input(4);
output(2, 54) <= input(5);
output(2, 55) <= input(6);
output(2, 56) <= input(7);
output(2, 57) <= input(8);
output(2, 58) <= input(9);
output(2, 59) <= input(10);
output(2, 60) <= input(11);
output(2, 61) <= input(12);
output(2, 62) <= input(13);
output(2, 63) <= input(14);
output(2, 64) <= input(33);
output(2, 65) <= input(16);
output(2, 66) <= input(17);
output(2, 67) <= input(18);
output(2, 68) <= input(19);
output(2, 69) <= input(20);
output(2, 70) <= input(21);
output(2, 71) <= input(22);
output(2, 72) <= input(23);
output(2, 73) <= input(24);
output(2, 74) <= input(25);
output(2, 75) <= input(26);
output(2, 76) <= input(27);
output(2, 77) <= input(28);
output(2, 78) <= input(29);
output(2, 79) <= input(30);
output(2, 80) <= input(33);
output(2, 81) <= input(16);
output(2, 82) <= input(17);
output(2, 83) <= input(18);
output(2, 84) <= input(19);
output(2, 85) <= input(20);
output(2, 86) <= input(21);
output(2, 87) <= input(22);
output(2, 88) <= input(23);
output(2, 89) <= input(24);
output(2, 90) <= input(25);
output(2, 91) <= input(26);
output(2, 92) <= input(27);
output(2, 93) <= input(28);
output(2, 94) <= input(29);
output(2, 95) <= input(30);
output(2, 96) <= input(34);
output(2, 97) <= input(32);
output(2, 98) <= input(0);
output(2, 99) <= input(1);
output(2, 100) <= input(2);
output(2, 101) <= input(3);
output(2, 102) <= input(4);
output(2, 103) <= input(5);
output(2, 104) <= input(6);
output(2, 105) <= input(7);
output(2, 106) <= input(8);
output(2, 107) <= input(9);
output(2, 108) <= input(10);
output(2, 109) <= input(11);
output(2, 110) <= input(12);
output(2, 111) <= input(13);
output(2, 112) <= input(34);
output(2, 113) <= input(32);
output(2, 114) <= input(0);
output(2, 115) <= input(1);
output(2, 116) <= input(2);
output(2, 117) <= input(3);
output(2, 118) <= input(4);
output(2, 119) <= input(5);
output(2, 120) <= input(6);
output(2, 121) <= input(7);
output(2, 122) <= input(8);
output(2, 123) <= input(9);
output(2, 124) <= input(10);
output(2, 125) <= input(11);
output(2, 126) <= input(12);
output(2, 127) <= input(13);
output(2, 128) <= input(35);
output(2, 129) <= input(33);
output(2, 130) <= input(16);
output(2, 131) <= input(17);
output(2, 132) <= input(18);
output(2, 133) <= input(19);
output(2, 134) <= input(20);
output(2, 135) <= input(21);
output(2, 136) <= input(22);
output(2, 137) <= input(23);
output(2, 138) <= input(24);
output(2, 139) <= input(25);
output(2, 140) <= input(26);
output(2, 141) <= input(27);
output(2, 142) <= input(28);
output(2, 143) <= input(29);
output(2, 144) <= input(36);
output(2, 145) <= input(34);
output(2, 146) <= input(32);
output(2, 147) <= input(0);
output(2, 148) <= input(1);
output(2, 149) <= input(2);
output(2, 150) <= input(3);
output(2, 151) <= input(4);
output(2, 152) <= input(5);
output(2, 153) <= input(6);
output(2, 154) <= input(7);
output(2, 155) <= input(8);
output(2, 156) <= input(9);
output(2, 157) <= input(10);
output(2, 158) <= input(11);
output(2, 159) <= input(12);
output(2, 160) <= input(36);
output(2, 161) <= input(34);
output(2, 162) <= input(32);
output(2, 163) <= input(0);
output(2, 164) <= input(1);
output(2, 165) <= input(2);
output(2, 166) <= input(3);
output(2, 167) <= input(4);
output(2, 168) <= input(5);
output(2, 169) <= input(6);
output(2, 170) <= input(7);
output(2, 171) <= input(8);
output(2, 172) <= input(9);
output(2, 173) <= input(10);
output(2, 174) <= input(11);
output(2, 175) <= input(12);
output(2, 176) <= input(37);
output(2, 177) <= input(35);
output(2, 178) <= input(33);
output(2, 179) <= input(16);
output(2, 180) <= input(17);
output(2, 181) <= input(18);
output(2, 182) <= input(19);
output(2, 183) <= input(20);
output(2, 184) <= input(21);
output(2, 185) <= input(22);
output(2, 186) <= input(23);
output(2, 187) <= input(24);
output(2, 188) <= input(25);
output(2, 189) <= input(26);
output(2, 190) <= input(27);
output(2, 191) <= input(28);
output(2, 192) <= input(38);
output(2, 193) <= input(36);
output(2, 194) <= input(34);
output(2, 195) <= input(32);
output(2, 196) <= input(0);
output(2, 197) <= input(1);
output(2, 198) <= input(2);
output(2, 199) <= input(3);
output(2, 200) <= input(4);
output(2, 201) <= input(5);
output(2, 202) <= input(6);
output(2, 203) <= input(7);
output(2, 204) <= input(8);
output(2, 205) <= input(9);
output(2, 206) <= input(10);
output(2, 207) <= input(11);
output(2, 208) <= input(38);
output(2, 209) <= input(36);
output(2, 210) <= input(34);
output(2, 211) <= input(32);
output(2, 212) <= input(0);
output(2, 213) <= input(1);
output(2, 214) <= input(2);
output(2, 215) <= input(3);
output(2, 216) <= input(4);
output(2, 217) <= input(5);
output(2, 218) <= input(6);
output(2, 219) <= input(7);
output(2, 220) <= input(8);
output(2, 221) <= input(9);
output(2, 222) <= input(10);
output(2, 223) <= input(11);
output(2, 224) <= input(39);
output(2, 225) <= input(37);
output(2, 226) <= input(35);
output(2, 227) <= input(33);
output(2, 228) <= input(16);
output(2, 229) <= input(17);
output(2, 230) <= input(18);
output(2, 231) <= input(19);
output(2, 232) <= input(20);
output(2, 233) <= input(21);
output(2, 234) <= input(22);
output(2, 235) <= input(23);
output(2, 236) <= input(24);
output(2, 237) <= input(25);
output(2, 238) <= input(26);
output(2, 239) <= input(27);
output(2, 240) <= input(39);
output(2, 241) <= input(37);
output(2, 242) <= input(35);
output(2, 243) <= input(33);
output(2, 244) <= input(16);
output(2, 245) <= input(17);
output(2, 246) <= input(18);
output(2, 247) <= input(19);
output(2, 248) <= input(20);
output(2, 249) <= input(21);
output(2, 250) <= input(22);
output(2, 251) <= input(23);
output(2, 252) <= input(24);
output(2, 253) <= input(25);
output(2, 254) <= input(26);
output(2, 255) <= input(27);
when "1100" =>
output(0, 0) <= input(0);
output(0, 1) <= input(1);
output(0, 2) <= input(2);
output(0, 3) <= input(3);
output(0, 4) <= input(4);
output(0, 5) <= input(5);
output(0, 6) <= input(6);
output(0, 7) <= input(7);
output(0, 8) <= input(8);
output(0, 9) <= input(9);
output(0, 10) <= input(10);
output(0, 11) <= input(11);
output(0, 12) <= input(12);
output(0, 13) <= input(13);
output(0, 14) <= input(14);
output(0, 15) <= input(15);
output(0, 16) <= input(0);
output(0, 17) <= input(1);
output(0, 18) <= input(2);
output(0, 19) <= input(3);
output(0, 20) <= input(4);
output(0, 21) <= input(5);
output(0, 22) <= input(6);
output(0, 23) <= input(7);
output(0, 24) <= input(8);
output(0, 25) <= input(9);
output(0, 26) <= input(10);
output(0, 27) <= input(11);
output(0, 28) <= input(12);
output(0, 29) <= input(13);
output(0, 30) <= input(14);
output(0, 31) <= input(15);
output(0, 32) <= input(16);
output(0, 33) <= input(17);
output(0, 34) <= input(18);
output(0, 35) <= input(19);
output(0, 36) <= input(20);
output(0, 37) <= input(21);
output(0, 38) <= input(22);
output(0, 39) <= input(23);
output(0, 40) <= input(24);
output(0, 41) <= input(25);
output(0, 42) <= input(26);
output(0, 43) <= input(27);
output(0, 44) <= input(28);
output(0, 45) <= input(29);
output(0, 46) <= input(30);
output(0, 47) <= input(31);
output(0, 48) <= input(16);
output(0, 49) <= input(17);
output(0, 50) <= input(18);
output(0, 51) <= input(19);
output(0, 52) <= input(20);
output(0, 53) <= input(21);
output(0, 54) <= input(22);
output(0, 55) <= input(23);
output(0, 56) <= input(24);
output(0, 57) <= input(25);
output(0, 58) <= input(26);
output(0, 59) <= input(27);
output(0, 60) <= input(28);
output(0, 61) <= input(29);
output(0, 62) <= input(30);
output(0, 63) <= input(31);
output(0, 64) <= input(32);
output(0, 65) <= input(0);
output(0, 66) <= input(1);
output(0, 67) <= input(2);
output(0, 68) <= input(3);
output(0, 69) <= input(4);
output(0, 70) <= input(5);
output(0, 71) <= input(6);
output(0, 72) <= input(7);
output(0, 73) <= input(8);
output(0, 74) <= input(9);
output(0, 75) <= input(10);
output(0, 76) <= input(11);
output(0, 77) <= input(12);
output(0, 78) <= input(13);
output(0, 79) <= input(14);
output(0, 80) <= input(32);
output(0, 81) <= input(0);
output(0, 82) <= input(1);
output(0, 83) <= input(2);
output(0, 84) <= input(3);
output(0, 85) <= input(4);
output(0, 86) <= input(5);
output(0, 87) <= input(6);
output(0, 88) <= input(7);
output(0, 89) <= input(8);
output(0, 90) <= input(9);
output(0, 91) <= input(10);
output(0, 92) <= input(11);
output(0, 93) <= input(12);
output(0, 94) <= input(13);
output(0, 95) <= input(14);
output(0, 96) <= input(33);
output(0, 97) <= input(16);
output(0, 98) <= input(17);
output(0, 99) <= input(18);
output(0, 100) <= input(19);
output(0, 101) <= input(20);
output(0, 102) <= input(21);
output(0, 103) <= input(22);
output(0, 104) <= input(23);
output(0, 105) <= input(24);
output(0, 106) <= input(25);
output(0, 107) <= input(26);
output(0, 108) <= input(27);
output(0, 109) <= input(28);
output(0, 110) <= input(29);
output(0, 111) <= input(30);
output(0, 112) <= input(33);
output(0, 113) <= input(16);
output(0, 114) <= input(17);
output(0, 115) <= input(18);
output(0, 116) <= input(19);
output(0, 117) <= input(20);
output(0, 118) <= input(21);
output(0, 119) <= input(22);
output(0, 120) <= input(23);
output(0, 121) <= input(24);
output(0, 122) <= input(25);
output(0, 123) <= input(26);
output(0, 124) <= input(27);
output(0, 125) <= input(28);
output(0, 126) <= input(29);
output(0, 127) <= input(30);
output(0, 128) <= input(34);
output(0, 129) <= input(32);
output(0, 130) <= input(0);
output(0, 131) <= input(1);
output(0, 132) <= input(2);
output(0, 133) <= input(3);
output(0, 134) <= input(4);
output(0, 135) <= input(5);
output(0, 136) <= input(6);
output(0, 137) <= input(7);
output(0, 138) <= input(8);
output(0, 139) <= input(9);
output(0, 140) <= input(10);
output(0, 141) <= input(11);
output(0, 142) <= input(12);
output(0, 143) <= input(13);
output(0, 144) <= input(34);
output(0, 145) <= input(32);
output(0, 146) <= input(0);
output(0, 147) <= input(1);
output(0, 148) <= input(2);
output(0, 149) <= input(3);
output(0, 150) <= input(4);
output(0, 151) <= input(5);
output(0, 152) <= input(6);
output(0, 153) <= input(7);
output(0, 154) <= input(8);
output(0, 155) <= input(9);
output(0, 156) <= input(10);
output(0, 157) <= input(11);
output(0, 158) <= input(12);
output(0, 159) <= input(13);
output(0, 160) <= input(35);
output(0, 161) <= input(33);
output(0, 162) <= input(16);
output(0, 163) <= input(17);
output(0, 164) <= input(18);
output(0, 165) <= input(19);
output(0, 166) <= input(20);
output(0, 167) <= input(21);
output(0, 168) <= input(22);
output(0, 169) <= input(23);
output(0, 170) <= input(24);
output(0, 171) <= input(25);
output(0, 172) <= input(26);
output(0, 173) <= input(27);
output(0, 174) <= input(28);
output(0, 175) <= input(29);
output(0, 176) <= input(35);
output(0, 177) <= input(33);
output(0, 178) <= input(16);
output(0, 179) <= input(17);
output(0, 180) <= input(18);
output(0, 181) <= input(19);
output(0, 182) <= input(20);
output(0, 183) <= input(21);
output(0, 184) <= input(22);
output(0, 185) <= input(23);
output(0, 186) <= input(24);
output(0, 187) <= input(25);
output(0, 188) <= input(26);
output(0, 189) <= input(27);
output(0, 190) <= input(28);
output(0, 191) <= input(29);
output(0, 192) <= input(36);
output(0, 193) <= input(34);
output(0, 194) <= input(32);
output(0, 195) <= input(0);
output(0, 196) <= input(1);
output(0, 197) <= input(2);
output(0, 198) <= input(3);
output(0, 199) <= input(4);
output(0, 200) <= input(5);
output(0, 201) <= input(6);
output(0, 202) <= input(7);
output(0, 203) <= input(8);
output(0, 204) <= input(9);
output(0, 205) <= input(10);
output(0, 206) <= input(11);
output(0, 207) <= input(12);
output(0, 208) <= input(36);
output(0, 209) <= input(34);
output(0, 210) <= input(32);
output(0, 211) <= input(0);
output(0, 212) <= input(1);
output(0, 213) <= input(2);
output(0, 214) <= input(3);
output(0, 215) <= input(4);
output(0, 216) <= input(5);
output(0, 217) <= input(6);
output(0, 218) <= input(7);
output(0, 219) <= input(8);
output(0, 220) <= input(9);
output(0, 221) <= input(10);
output(0, 222) <= input(11);
output(0, 223) <= input(12);
output(0, 224) <= input(37);
output(0, 225) <= input(35);
output(0, 226) <= input(33);
output(0, 227) <= input(16);
output(0, 228) <= input(17);
output(0, 229) <= input(18);
output(0, 230) <= input(19);
output(0, 231) <= input(20);
output(0, 232) <= input(21);
output(0, 233) <= input(22);
output(0, 234) <= input(23);
output(0, 235) <= input(24);
output(0, 236) <= input(25);
output(0, 237) <= input(26);
output(0, 238) <= input(27);
output(0, 239) <= input(28);
output(0, 240) <= input(37);
output(0, 241) <= input(35);
output(0, 242) <= input(33);
output(0, 243) <= input(16);
output(0, 244) <= input(17);
output(0, 245) <= input(18);
output(0, 246) <= input(19);
output(0, 247) <= input(20);
output(0, 248) <= input(21);
output(0, 249) <= input(22);
output(0, 250) <= input(23);
output(0, 251) <= input(24);
output(0, 252) <= input(25);
output(0, 253) <= input(26);
output(0, 254) <= input(27);
output(0, 255) <= input(28);
output(1, 0) <= input(0);
output(1, 1) <= input(1);
output(1, 2) <= input(2);
output(1, 3) <= input(3);
output(1, 4) <= input(4);
output(1, 5) <= input(5);
output(1, 6) <= input(6);
output(1, 7) <= input(7);
output(1, 8) <= input(8);
output(1, 9) <= input(9);
output(1, 10) <= input(10);
output(1, 11) <= input(11);
output(1, 12) <= input(12);
output(1, 13) <= input(13);
output(1, 14) <= input(14);
output(1, 15) <= input(15);
output(1, 16) <= input(0);
output(1, 17) <= input(1);
output(1, 18) <= input(2);
output(1, 19) <= input(3);
output(1, 20) <= input(4);
output(1, 21) <= input(5);
output(1, 22) <= input(6);
output(1, 23) <= input(7);
output(1, 24) <= input(8);
output(1, 25) <= input(9);
output(1, 26) <= input(10);
output(1, 27) <= input(11);
output(1, 28) <= input(12);
output(1, 29) <= input(13);
output(1, 30) <= input(14);
output(1, 31) <= input(15);
output(1, 32) <= input(16);
output(1, 33) <= input(17);
output(1, 34) <= input(18);
output(1, 35) <= input(19);
output(1, 36) <= input(20);
output(1, 37) <= input(21);
output(1, 38) <= input(22);
output(1, 39) <= input(23);
output(1, 40) <= input(24);
output(1, 41) <= input(25);
output(1, 42) <= input(26);
output(1, 43) <= input(27);
output(1, 44) <= input(28);
output(1, 45) <= input(29);
output(1, 46) <= input(30);
output(1, 47) <= input(31);
output(1, 48) <= input(16);
output(1, 49) <= input(17);
output(1, 50) <= input(18);
output(1, 51) <= input(19);
output(1, 52) <= input(20);
output(1, 53) <= input(21);
output(1, 54) <= input(22);
output(1, 55) <= input(23);
output(1, 56) <= input(24);
output(1, 57) <= input(25);
output(1, 58) <= input(26);
output(1, 59) <= input(27);
output(1, 60) <= input(28);
output(1, 61) <= input(29);
output(1, 62) <= input(30);
output(1, 63) <= input(31);
output(1, 64) <= input(16);
output(1, 65) <= input(17);
output(1, 66) <= input(18);
output(1, 67) <= input(19);
output(1, 68) <= input(20);
output(1, 69) <= input(21);
output(1, 70) <= input(22);
output(1, 71) <= input(23);
output(1, 72) <= input(24);
output(1, 73) <= input(25);
output(1, 74) <= input(26);
output(1, 75) <= input(27);
output(1, 76) <= input(28);
output(1, 77) <= input(29);
output(1, 78) <= input(30);
output(1, 79) <= input(31);
output(1, 80) <= input(32);
output(1, 81) <= input(0);
output(1, 82) <= input(1);
output(1, 83) <= input(2);
output(1, 84) <= input(3);
output(1, 85) <= input(4);
output(1, 86) <= input(5);
output(1, 87) <= input(6);
output(1, 88) <= input(7);
output(1, 89) <= input(8);
output(1, 90) <= input(9);
output(1, 91) <= input(10);
output(1, 92) <= input(11);
output(1, 93) <= input(12);
output(1, 94) <= input(13);
output(1, 95) <= input(14);
output(1, 96) <= input(32);
output(1, 97) <= input(0);
output(1, 98) <= input(1);
output(1, 99) <= input(2);
output(1, 100) <= input(3);
output(1, 101) <= input(4);
output(1, 102) <= input(5);
output(1, 103) <= input(6);
output(1, 104) <= input(7);
output(1, 105) <= input(8);
output(1, 106) <= input(9);
output(1, 107) <= input(10);
output(1, 108) <= input(11);
output(1, 109) <= input(12);
output(1, 110) <= input(13);
output(1, 111) <= input(14);
output(1, 112) <= input(32);
output(1, 113) <= input(0);
output(1, 114) <= input(1);
output(1, 115) <= input(2);
output(1, 116) <= input(3);
output(1, 117) <= input(4);
output(1, 118) <= input(5);
output(1, 119) <= input(6);
output(1, 120) <= input(7);
output(1, 121) <= input(8);
output(1, 122) <= input(9);
output(1, 123) <= input(10);
output(1, 124) <= input(11);
output(1, 125) <= input(12);
output(1, 126) <= input(13);
output(1, 127) <= input(14);
output(1, 128) <= input(33);
output(1, 129) <= input(16);
output(1, 130) <= input(17);
output(1, 131) <= input(18);
output(1, 132) <= input(19);
output(1, 133) <= input(20);
output(1, 134) <= input(21);
output(1, 135) <= input(22);
output(1, 136) <= input(23);
output(1, 137) <= input(24);
output(1, 138) <= input(25);
output(1, 139) <= input(26);
output(1, 140) <= input(27);
output(1, 141) <= input(28);
output(1, 142) <= input(29);
output(1, 143) <= input(30);
output(1, 144) <= input(33);
output(1, 145) <= input(16);
output(1, 146) <= input(17);
output(1, 147) <= input(18);
output(1, 148) <= input(19);
output(1, 149) <= input(20);
output(1, 150) <= input(21);
output(1, 151) <= input(22);
output(1, 152) <= input(23);
output(1, 153) <= input(24);
output(1, 154) <= input(25);
output(1, 155) <= input(26);
output(1, 156) <= input(27);
output(1, 157) <= input(28);
output(1, 158) <= input(29);
output(1, 159) <= input(30);
output(1, 160) <= input(34);
output(1, 161) <= input(32);
output(1, 162) <= input(0);
output(1, 163) <= input(1);
output(1, 164) <= input(2);
output(1, 165) <= input(3);
output(1, 166) <= input(4);
output(1, 167) <= input(5);
output(1, 168) <= input(6);
output(1, 169) <= input(7);
output(1, 170) <= input(8);
output(1, 171) <= input(9);
output(1, 172) <= input(10);
output(1, 173) <= input(11);
output(1, 174) <= input(12);
output(1, 175) <= input(13);
output(1, 176) <= input(34);
output(1, 177) <= input(32);
output(1, 178) <= input(0);
output(1, 179) <= input(1);
output(1, 180) <= input(2);
output(1, 181) <= input(3);
output(1, 182) <= input(4);
output(1, 183) <= input(5);
output(1, 184) <= input(6);
output(1, 185) <= input(7);
output(1, 186) <= input(8);
output(1, 187) <= input(9);
output(1, 188) <= input(10);
output(1, 189) <= input(11);
output(1, 190) <= input(12);
output(1, 191) <= input(13);
output(1, 192) <= input(34);
output(1, 193) <= input(32);
output(1, 194) <= input(0);
output(1, 195) <= input(1);
output(1, 196) <= input(2);
output(1, 197) <= input(3);
output(1, 198) <= input(4);
output(1, 199) <= input(5);
output(1, 200) <= input(6);
output(1, 201) <= input(7);
output(1, 202) <= input(8);
output(1, 203) <= input(9);
output(1, 204) <= input(10);
output(1, 205) <= input(11);
output(1, 206) <= input(12);
output(1, 207) <= input(13);
output(1, 208) <= input(35);
output(1, 209) <= input(33);
output(1, 210) <= input(16);
output(1, 211) <= input(17);
output(1, 212) <= input(18);
output(1, 213) <= input(19);
output(1, 214) <= input(20);
output(1, 215) <= input(21);
output(1, 216) <= input(22);
output(1, 217) <= input(23);
output(1, 218) <= input(24);
output(1, 219) <= input(25);
output(1, 220) <= input(26);
output(1, 221) <= input(27);
output(1, 222) <= input(28);
output(1, 223) <= input(29);
output(1, 224) <= input(35);
output(1, 225) <= input(33);
output(1, 226) <= input(16);
output(1, 227) <= input(17);
output(1, 228) <= input(18);
output(1, 229) <= input(19);
output(1, 230) <= input(20);
output(1, 231) <= input(21);
output(1, 232) <= input(22);
output(1, 233) <= input(23);
output(1, 234) <= input(24);
output(1, 235) <= input(25);
output(1, 236) <= input(26);
output(1, 237) <= input(27);
output(1, 238) <= input(28);
output(1, 239) <= input(29);
output(1, 240) <= input(35);
output(1, 241) <= input(33);
output(1, 242) <= input(16);
output(1, 243) <= input(17);
output(1, 244) <= input(18);
output(1, 245) <= input(19);
output(1, 246) <= input(20);
output(1, 247) <= input(21);
output(1, 248) <= input(22);
output(1, 249) <= input(23);
output(1, 250) <= input(24);
output(1, 251) <= input(25);
output(1, 252) <= input(26);
output(1, 253) <= input(27);
output(1, 254) <= input(28);
output(1, 255) <= input(29);
output(2, 0) <= input(0);
output(2, 1) <= input(1);
output(2, 2) <= input(2);
output(2, 3) <= input(3);
output(2, 4) <= input(4);
output(2, 5) <= input(5);
output(2, 6) <= input(6);
output(2, 7) <= input(7);
output(2, 8) <= input(8);
output(2, 9) <= input(9);
output(2, 10) <= input(10);
output(2, 11) <= input(11);
output(2, 12) <= input(12);
output(2, 13) <= input(13);
output(2, 14) <= input(14);
output(2, 15) <= input(15);
output(2, 16) <= input(0);
output(2, 17) <= input(1);
output(2, 18) <= input(2);
output(2, 19) <= input(3);
output(2, 20) <= input(4);
output(2, 21) <= input(5);
output(2, 22) <= input(6);
output(2, 23) <= input(7);
output(2, 24) <= input(8);
output(2, 25) <= input(9);
output(2, 26) <= input(10);
output(2, 27) <= input(11);
output(2, 28) <= input(12);
output(2, 29) <= input(13);
output(2, 30) <= input(14);
output(2, 31) <= input(15);
output(2, 32) <= input(0);
output(2, 33) <= input(1);
output(2, 34) <= input(2);
output(2, 35) <= input(3);
output(2, 36) <= input(4);
output(2, 37) <= input(5);
output(2, 38) <= input(6);
output(2, 39) <= input(7);
output(2, 40) <= input(8);
output(2, 41) <= input(9);
output(2, 42) <= input(10);
output(2, 43) <= input(11);
output(2, 44) <= input(12);
output(2, 45) <= input(13);
output(2, 46) <= input(14);
output(2, 47) <= input(15);
output(2, 48) <= input(0);
output(2, 49) <= input(1);
output(2, 50) <= input(2);
output(2, 51) <= input(3);
output(2, 52) <= input(4);
output(2, 53) <= input(5);
output(2, 54) <= input(6);
output(2, 55) <= input(7);
output(2, 56) <= input(8);
output(2, 57) <= input(9);
output(2, 58) <= input(10);
output(2, 59) <= input(11);
output(2, 60) <= input(12);
output(2, 61) <= input(13);
output(2, 62) <= input(14);
output(2, 63) <= input(15);
output(2, 64) <= input(16);
output(2, 65) <= input(17);
output(2, 66) <= input(18);
output(2, 67) <= input(19);
output(2, 68) <= input(20);
output(2, 69) <= input(21);
output(2, 70) <= input(22);
output(2, 71) <= input(23);
output(2, 72) <= input(24);
output(2, 73) <= input(25);
output(2, 74) <= input(26);
output(2, 75) <= input(27);
output(2, 76) <= input(28);
output(2, 77) <= input(29);
output(2, 78) <= input(30);
output(2, 79) <= input(31);
output(2, 80) <= input(16);
output(2, 81) <= input(17);
output(2, 82) <= input(18);
output(2, 83) <= input(19);
output(2, 84) <= input(20);
output(2, 85) <= input(21);
output(2, 86) <= input(22);
output(2, 87) <= input(23);
output(2, 88) <= input(24);
output(2, 89) <= input(25);
output(2, 90) <= input(26);
output(2, 91) <= input(27);
output(2, 92) <= input(28);
output(2, 93) <= input(29);
output(2, 94) <= input(30);
output(2, 95) <= input(31);
output(2, 96) <= input(16);
output(2, 97) <= input(17);
output(2, 98) <= input(18);
output(2, 99) <= input(19);
output(2, 100) <= input(20);
output(2, 101) <= input(21);
output(2, 102) <= input(22);
output(2, 103) <= input(23);
output(2, 104) <= input(24);
output(2, 105) <= input(25);
output(2, 106) <= input(26);
output(2, 107) <= input(27);
output(2, 108) <= input(28);
output(2, 109) <= input(29);
output(2, 110) <= input(30);
output(2, 111) <= input(31);
output(2, 112) <= input(16);
output(2, 113) <= input(17);
output(2, 114) <= input(18);
output(2, 115) <= input(19);
output(2, 116) <= input(20);
output(2, 117) <= input(21);
output(2, 118) <= input(22);
output(2, 119) <= input(23);
output(2, 120) <= input(24);
output(2, 121) <= input(25);
output(2, 122) <= input(26);
output(2, 123) <= input(27);
output(2, 124) <= input(28);
output(2, 125) <= input(29);
output(2, 126) <= input(30);
output(2, 127) <= input(31);
output(2, 128) <= input(32);
output(2, 129) <= input(0);
output(2, 130) <= input(1);
output(2, 131) <= input(2);
output(2, 132) <= input(3);
output(2, 133) <= input(4);
output(2, 134) <= input(5);
output(2, 135) <= input(6);
output(2, 136) <= input(7);
output(2, 137) <= input(8);
output(2, 138) <= input(9);
output(2, 139) <= input(10);
output(2, 140) <= input(11);
output(2, 141) <= input(12);
output(2, 142) <= input(13);
output(2, 143) <= input(14);
output(2, 144) <= input(32);
output(2, 145) <= input(0);
output(2, 146) <= input(1);
output(2, 147) <= input(2);
output(2, 148) <= input(3);
output(2, 149) <= input(4);
output(2, 150) <= input(5);
output(2, 151) <= input(6);
output(2, 152) <= input(7);
output(2, 153) <= input(8);
output(2, 154) <= input(9);
output(2, 155) <= input(10);
output(2, 156) <= input(11);
output(2, 157) <= input(12);
output(2, 158) <= input(13);
output(2, 159) <= input(14);
output(2, 160) <= input(32);
output(2, 161) <= input(0);
output(2, 162) <= input(1);
output(2, 163) <= input(2);
output(2, 164) <= input(3);
output(2, 165) <= input(4);
output(2, 166) <= input(5);
output(2, 167) <= input(6);
output(2, 168) <= input(7);
output(2, 169) <= input(8);
output(2, 170) <= input(9);
output(2, 171) <= input(10);
output(2, 172) <= input(11);
output(2, 173) <= input(12);
output(2, 174) <= input(13);
output(2, 175) <= input(14);
output(2, 176) <= input(32);
output(2, 177) <= input(0);
output(2, 178) <= input(1);
output(2, 179) <= input(2);
output(2, 180) <= input(3);
output(2, 181) <= input(4);
output(2, 182) <= input(5);
output(2, 183) <= input(6);
output(2, 184) <= input(7);
output(2, 185) <= input(8);
output(2, 186) <= input(9);
output(2, 187) <= input(10);
output(2, 188) <= input(11);
output(2, 189) <= input(12);
output(2, 190) <= input(13);
output(2, 191) <= input(14);
output(2, 192) <= input(33);
output(2, 193) <= input(16);
output(2, 194) <= input(17);
output(2, 195) <= input(18);
output(2, 196) <= input(19);
output(2, 197) <= input(20);
output(2, 198) <= input(21);
output(2, 199) <= input(22);
output(2, 200) <= input(23);
output(2, 201) <= input(24);
output(2, 202) <= input(25);
output(2, 203) <= input(26);
output(2, 204) <= input(27);
output(2, 205) <= input(28);
output(2, 206) <= input(29);
output(2, 207) <= input(30);
output(2, 208) <= input(33);
output(2, 209) <= input(16);
output(2, 210) <= input(17);
output(2, 211) <= input(18);
output(2, 212) <= input(19);
output(2, 213) <= input(20);
output(2, 214) <= input(21);
output(2, 215) <= input(22);
output(2, 216) <= input(23);
output(2, 217) <= input(24);
output(2, 218) <= input(25);
output(2, 219) <= input(26);
output(2, 220) <= input(27);
output(2, 221) <= input(28);
output(2, 222) <= input(29);
output(2, 223) <= input(30);
output(2, 224) <= input(33);
output(2, 225) <= input(16);
output(2, 226) <= input(17);
output(2, 227) <= input(18);
output(2, 228) <= input(19);
output(2, 229) <= input(20);
output(2, 230) <= input(21);
output(2, 231) <= input(22);
output(2, 232) <= input(23);
output(2, 233) <= input(24);
output(2, 234) <= input(25);
output(2, 235) <= input(26);
output(2, 236) <= input(27);
output(2, 237) <= input(28);
output(2, 238) <= input(29);
output(2, 239) <= input(30);
output(2, 240) <= input(33);
output(2, 241) <= input(16);
output(2, 242) <= input(17);
output(2, 243) <= input(18);
output(2, 244) <= input(19);
output(2, 245) <= input(20);
output(2, 246) <= input(21);
output(2, 247) <= input(22);
output(2, 248) <= input(23);
output(2, 249) <= input(24);
output(2, 250) <= input(25);
output(2, 251) <= input(26);
output(2, 252) <= input(27);
output(2, 253) <= input(28);
output(2, 254) <= input(29);
output(2, 255) <= input(30);
when "1101" =>
output(0, 0) <= input(0);
output(0, 1) <= input(1);
output(0, 2) <= input(2);
output(0, 3) <= input(3);
output(0, 4) <= input(4);
output(0, 5) <= input(5);
output(0, 6) <= input(6);
output(0, 7) <= input(7);
output(0, 8) <= input(8);
output(0, 9) <= input(9);
output(0, 10) <= input(10);
output(0, 11) <= input(11);
output(0, 12) <= input(12);
output(0, 13) <= input(13);
output(0, 14) <= input(14);
output(0, 15) <= input(15);
output(0, 16) <= input(0);
output(0, 17) <= input(1);
output(0, 18) <= input(2);
output(0, 19) <= input(3);
output(0, 20) <= input(4);
output(0, 21) <= input(5);
output(0, 22) <= input(6);
output(0, 23) <= input(7);
output(0, 24) <= input(8);
output(0, 25) <= input(9);
output(0, 26) <= input(10);
output(0, 27) <= input(11);
output(0, 28) <= input(12);
output(0, 29) <= input(13);
output(0, 30) <= input(14);
output(0, 31) <= input(15);
output(0, 32) <= input(0);
output(0, 33) <= input(1);
output(0, 34) <= input(2);
output(0, 35) <= input(3);
output(0, 36) <= input(4);
output(0, 37) <= input(5);
output(0, 38) <= input(6);
output(0, 39) <= input(7);
output(0, 40) <= input(8);
output(0, 41) <= input(9);
output(0, 42) <= input(10);
output(0, 43) <= input(11);
output(0, 44) <= input(12);
output(0, 45) <= input(13);
output(0, 46) <= input(14);
output(0, 47) <= input(15);
output(0, 48) <= input(0);
output(0, 49) <= input(1);
output(0, 50) <= input(2);
output(0, 51) <= input(3);
output(0, 52) <= input(4);
output(0, 53) <= input(5);
output(0, 54) <= input(6);
output(0, 55) <= input(7);
output(0, 56) <= input(8);
output(0, 57) <= input(9);
output(0, 58) <= input(10);
output(0, 59) <= input(11);
output(0, 60) <= input(12);
output(0, 61) <= input(13);
output(0, 62) <= input(14);
output(0, 63) <= input(15);
output(0, 64) <= input(0);
output(0, 65) <= input(1);
output(0, 66) <= input(2);
output(0, 67) <= input(3);
output(0, 68) <= input(4);
output(0, 69) <= input(5);
output(0, 70) <= input(6);
output(0, 71) <= input(7);
output(0, 72) <= input(8);
output(0, 73) <= input(9);
output(0, 74) <= input(10);
output(0, 75) <= input(11);
output(0, 76) <= input(12);
output(0, 77) <= input(13);
output(0, 78) <= input(14);
output(0, 79) <= input(15);
output(0, 80) <= input(16);
output(0, 81) <= input(17);
output(0, 82) <= input(18);
output(0, 83) <= input(19);
output(0, 84) <= input(20);
output(0, 85) <= input(21);
output(0, 86) <= input(22);
output(0, 87) <= input(23);
output(0, 88) <= input(24);
output(0, 89) <= input(25);
output(0, 90) <= input(26);
output(0, 91) <= input(27);
output(0, 92) <= input(28);
output(0, 93) <= input(29);
output(0, 94) <= input(30);
output(0, 95) <= input(31);
output(0, 96) <= input(16);
output(0, 97) <= input(17);
output(0, 98) <= input(18);
output(0, 99) <= input(19);
output(0, 100) <= input(20);
output(0, 101) <= input(21);
output(0, 102) <= input(22);
output(0, 103) <= input(23);
output(0, 104) <= input(24);
output(0, 105) <= input(25);
output(0, 106) <= input(26);
output(0, 107) <= input(27);
output(0, 108) <= input(28);
output(0, 109) <= input(29);
output(0, 110) <= input(30);
output(0, 111) <= input(31);
output(0, 112) <= input(16);
output(0, 113) <= input(17);
output(0, 114) <= input(18);
output(0, 115) <= input(19);
output(0, 116) <= input(20);
output(0, 117) <= input(21);
output(0, 118) <= input(22);
output(0, 119) <= input(23);
output(0, 120) <= input(24);
output(0, 121) <= input(25);
output(0, 122) <= input(26);
output(0, 123) <= input(27);
output(0, 124) <= input(28);
output(0, 125) <= input(29);
output(0, 126) <= input(30);
output(0, 127) <= input(31);
output(0, 128) <= input(16);
output(0, 129) <= input(17);
output(0, 130) <= input(18);
output(0, 131) <= input(19);
output(0, 132) <= input(20);
output(0, 133) <= input(21);
output(0, 134) <= input(22);
output(0, 135) <= input(23);
output(0, 136) <= input(24);
output(0, 137) <= input(25);
output(0, 138) <= input(26);
output(0, 139) <= input(27);
output(0, 140) <= input(28);
output(0, 141) <= input(29);
output(0, 142) <= input(30);
output(0, 143) <= input(31);
output(0, 144) <= input(16);
output(0, 145) <= input(17);
output(0, 146) <= input(18);
output(0, 147) <= input(19);
output(0, 148) <= input(20);
output(0, 149) <= input(21);
output(0, 150) <= input(22);
output(0, 151) <= input(23);
output(0, 152) <= input(24);
output(0, 153) <= input(25);
output(0, 154) <= input(26);
output(0, 155) <= input(27);
output(0, 156) <= input(28);
output(0, 157) <= input(29);
output(0, 158) <= input(30);
output(0, 159) <= input(31);
output(0, 160) <= input(32);
output(0, 161) <= input(0);
output(0, 162) <= input(1);
output(0, 163) <= input(2);
output(0, 164) <= input(3);
output(0, 165) <= input(4);
output(0, 166) <= input(5);
output(0, 167) <= input(6);
output(0, 168) <= input(7);
output(0, 169) <= input(8);
output(0, 170) <= input(9);
output(0, 171) <= input(10);
output(0, 172) <= input(11);
output(0, 173) <= input(12);
output(0, 174) <= input(13);
output(0, 175) <= input(14);
output(0, 176) <= input(32);
output(0, 177) <= input(0);
output(0, 178) <= input(1);
output(0, 179) <= input(2);
output(0, 180) <= input(3);
output(0, 181) <= input(4);
output(0, 182) <= input(5);
output(0, 183) <= input(6);
output(0, 184) <= input(7);
output(0, 185) <= input(8);
output(0, 186) <= input(9);
output(0, 187) <= input(10);
output(0, 188) <= input(11);
output(0, 189) <= input(12);
output(0, 190) <= input(13);
output(0, 191) <= input(14);
output(0, 192) <= input(32);
output(0, 193) <= input(0);
output(0, 194) <= input(1);
output(0, 195) <= input(2);
output(0, 196) <= input(3);
output(0, 197) <= input(4);
output(0, 198) <= input(5);
output(0, 199) <= input(6);
output(0, 200) <= input(7);
output(0, 201) <= input(8);
output(0, 202) <= input(9);
output(0, 203) <= input(10);
output(0, 204) <= input(11);
output(0, 205) <= input(12);
output(0, 206) <= input(13);
output(0, 207) <= input(14);
output(0, 208) <= input(32);
output(0, 209) <= input(0);
output(0, 210) <= input(1);
output(0, 211) <= input(2);
output(0, 212) <= input(3);
output(0, 213) <= input(4);
output(0, 214) <= input(5);
output(0, 215) <= input(6);
output(0, 216) <= input(7);
output(0, 217) <= input(8);
output(0, 218) <= input(9);
output(0, 219) <= input(10);
output(0, 220) <= input(11);
output(0, 221) <= input(12);
output(0, 222) <= input(13);
output(0, 223) <= input(14);
output(0, 224) <= input(32);
output(0, 225) <= input(0);
output(0, 226) <= input(1);
output(0, 227) <= input(2);
output(0, 228) <= input(3);
output(0, 229) <= input(4);
output(0, 230) <= input(5);
output(0, 231) <= input(6);
output(0, 232) <= input(7);
output(0, 233) <= input(8);
output(0, 234) <= input(9);
output(0, 235) <= input(10);
output(0, 236) <= input(11);
output(0, 237) <= input(12);
output(0, 238) <= input(13);
output(0, 239) <= input(14);
output(0, 240) <= input(32);
output(0, 241) <= input(0);
output(0, 242) <= input(1);
output(0, 243) <= input(2);
output(0, 244) <= input(3);
output(0, 245) <= input(4);
output(0, 246) <= input(5);
output(0, 247) <= input(6);
output(0, 248) <= input(7);
output(0, 249) <= input(8);
output(0, 250) <= input(9);
output(0, 251) <= input(10);
output(0, 252) <= input(11);
output(0, 253) <= input(12);
output(0, 254) <= input(13);
output(0, 255) <= input(14);
output(1, 0) <= input(0);
output(1, 1) <= input(1);
output(1, 2) <= input(2);
output(1, 3) <= input(3);
output(1, 4) <= input(4);
output(1, 5) <= input(5);
output(1, 6) <= input(6);
output(1, 7) <= input(7);
output(1, 8) <= input(8);
output(1, 9) <= input(9);
output(1, 10) <= input(10);
output(1, 11) <= input(11);
output(1, 12) <= input(12);
output(1, 13) <= input(13);
output(1, 14) <= input(14);
output(1, 15) <= input(15);
output(1, 16) <= input(0);
output(1, 17) <= input(1);
output(1, 18) <= input(2);
output(1, 19) <= input(3);
output(1, 20) <= input(4);
output(1, 21) <= input(5);
output(1, 22) <= input(6);
output(1, 23) <= input(7);
output(1, 24) <= input(8);
output(1, 25) <= input(9);
output(1, 26) <= input(10);
output(1, 27) <= input(11);
output(1, 28) <= input(12);
output(1, 29) <= input(13);
output(1, 30) <= input(14);
output(1, 31) <= input(15);
output(1, 32) <= input(0);
output(1, 33) <= input(1);
output(1, 34) <= input(2);
output(1, 35) <= input(3);
output(1, 36) <= input(4);
output(1, 37) <= input(5);
output(1, 38) <= input(6);
output(1, 39) <= input(7);
output(1, 40) <= input(8);
output(1, 41) <= input(9);
output(1, 42) <= input(10);
output(1, 43) <= input(11);
output(1, 44) <= input(12);
output(1, 45) <= input(13);
output(1, 46) <= input(14);
output(1, 47) <= input(15);
output(1, 48) <= input(0);
output(1, 49) <= input(1);
output(1, 50) <= input(2);
output(1, 51) <= input(3);
output(1, 52) <= input(4);
output(1, 53) <= input(5);
output(1, 54) <= input(6);
output(1, 55) <= input(7);
output(1, 56) <= input(8);
output(1, 57) <= input(9);
output(1, 58) <= input(10);
output(1, 59) <= input(11);
output(1, 60) <= input(12);
output(1, 61) <= input(13);
output(1, 62) <= input(14);
output(1, 63) <= input(15);
output(1, 64) <= input(0);
output(1, 65) <= input(1);
output(1, 66) <= input(2);
output(1, 67) <= input(3);
output(1, 68) <= input(4);
output(1, 69) <= input(5);
output(1, 70) <= input(6);
output(1, 71) <= input(7);
output(1, 72) <= input(8);
output(1, 73) <= input(9);
output(1, 74) <= input(10);
output(1, 75) <= input(11);
output(1, 76) <= input(12);
output(1, 77) <= input(13);
output(1, 78) <= input(14);
output(1, 79) <= input(15);
output(1, 80) <= input(0);
output(1, 81) <= input(1);
output(1, 82) <= input(2);
output(1, 83) <= input(3);
output(1, 84) <= input(4);
output(1, 85) <= input(5);
output(1, 86) <= input(6);
output(1, 87) <= input(7);
output(1, 88) <= input(8);
output(1, 89) <= input(9);
output(1, 90) <= input(10);
output(1, 91) <= input(11);
output(1, 92) <= input(12);
output(1, 93) <= input(13);
output(1, 94) <= input(14);
output(1, 95) <= input(15);
output(1, 96) <= input(0);
output(1, 97) <= input(1);
output(1, 98) <= input(2);
output(1, 99) <= input(3);
output(1, 100) <= input(4);
output(1, 101) <= input(5);
output(1, 102) <= input(6);
output(1, 103) <= input(7);
output(1, 104) <= input(8);
output(1, 105) <= input(9);
output(1, 106) <= input(10);
output(1, 107) <= input(11);
output(1, 108) <= input(12);
output(1, 109) <= input(13);
output(1, 110) <= input(14);
output(1, 111) <= input(15);
output(1, 112) <= input(0);
output(1, 113) <= input(1);
output(1, 114) <= input(2);
output(1, 115) <= input(3);
output(1, 116) <= input(4);
output(1, 117) <= input(5);
output(1, 118) <= input(6);
output(1, 119) <= input(7);
output(1, 120) <= input(8);
output(1, 121) <= input(9);
output(1, 122) <= input(10);
output(1, 123) <= input(11);
output(1, 124) <= input(12);
output(1, 125) <= input(13);
output(1, 126) <= input(14);
output(1, 127) <= input(15);
output(1, 128) <= input(16);
output(1, 129) <= input(17);
output(1, 130) <= input(18);
output(1, 131) <= input(19);
output(1, 132) <= input(20);
output(1, 133) <= input(21);
output(1, 134) <= input(22);
output(1, 135) <= input(23);
output(1, 136) <= input(24);
output(1, 137) <= input(25);
output(1, 138) <= input(26);
output(1, 139) <= input(27);
output(1, 140) <= input(28);
output(1, 141) <= input(29);
output(1, 142) <= input(30);
output(1, 143) <= input(31);
output(1, 144) <= input(16);
output(1, 145) <= input(17);
output(1, 146) <= input(18);
output(1, 147) <= input(19);
output(1, 148) <= input(20);
output(1, 149) <= input(21);
output(1, 150) <= input(22);
output(1, 151) <= input(23);
output(1, 152) <= input(24);
output(1, 153) <= input(25);
output(1, 154) <= input(26);
output(1, 155) <= input(27);
output(1, 156) <= input(28);
output(1, 157) <= input(29);
output(1, 158) <= input(30);
output(1, 159) <= input(31);
output(1, 160) <= input(16);
output(1, 161) <= input(17);
output(1, 162) <= input(18);
output(1, 163) <= input(19);
output(1, 164) <= input(20);
output(1, 165) <= input(21);
output(1, 166) <= input(22);
output(1, 167) <= input(23);
output(1, 168) <= input(24);
output(1, 169) <= input(25);
output(1, 170) <= input(26);
output(1, 171) <= input(27);
output(1, 172) <= input(28);
output(1, 173) <= input(29);
output(1, 174) <= input(30);
output(1, 175) <= input(31);
output(1, 176) <= input(16);
output(1, 177) <= input(17);
output(1, 178) <= input(18);
output(1, 179) <= input(19);
output(1, 180) <= input(20);
output(1, 181) <= input(21);
output(1, 182) <= input(22);
output(1, 183) <= input(23);
output(1, 184) <= input(24);
output(1, 185) <= input(25);
output(1, 186) <= input(26);
output(1, 187) <= input(27);
output(1, 188) <= input(28);
output(1, 189) <= input(29);
output(1, 190) <= input(30);
output(1, 191) <= input(31);
output(1, 192) <= input(16);
output(1, 193) <= input(17);
output(1, 194) <= input(18);
output(1, 195) <= input(19);
output(1, 196) <= input(20);
output(1, 197) <= input(21);
output(1, 198) <= input(22);
output(1, 199) <= input(23);
output(1, 200) <= input(24);
output(1, 201) <= input(25);
output(1, 202) <= input(26);
output(1, 203) <= input(27);
output(1, 204) <= input(28);
output(1, 205) <= input(29);
output(1, 206) <= input(30);
output(1, 207) <= input(31);
output(1, 208) <= input(16);
output(1, 209) <= input(17);
output(1, 210) <= input(18);
output(1, 211) <= input(19);
output(1, 212) <= input(20);
output(1, 213) <= input(21);
output(1, 214) <= input(22);
output(1, 215) <= input(23);
output(1, 216) <= input(24);
output(1, 217) <= input(25);
output(1, 218) <= input(26);
output(1, 219) <= input(27);
output(1, 220) <= input(28);
output(1, 221) <= input(29);
output(1, 222) <= input(30);
output(1, 223) <= input(31);
output(1, 224) <= input(16);
output(1, 225) <= input(17);
output(1, 226) <= input(18);
output(1, 227) <= input(19);
output(1, 228) <= input(20);
output(1, 229) <= input(21);
output(1, 230) <= input(22);
output(1, 231) <= input(23);
output(1, 232) <= input(24);
output(1, 233) <= input(25);
output(1, 234) <= input(26);
output(1, 235) <= input(27);
output(1, 236) <= input(28);
output(1, 237) <= input(29);
output(1, 238) <= input(30);
output(1, 239) <= input(31);
output(1, 240) <= input(16);
output(1, 241) <= input(17);
output(1, 242) <= input(18);
output(1, 243) <= input(19);
output(1, 244) <= input(20);
output(1, 245) <= input(21);
output(1, 246) <= input(22);
output(1, 247) <= input(23);
output(1, 248) <= input(24);
output(1, 249) <= input(25);
output(1, 250) <= input(26);
output(1, 251) <= input(27);
output(1, 252) <= input(28);
output(1, 253) <= input(29);
output(1, 254) <= input(30);
output(1, 255) <= input(31);
output(2, 0) <= input(0);
output(2, 1) <= input(1);
output(2, 2) <= input(2);
output(2, 3) <= input(3);
output(2, 4) <= input(4);
output(2, 5) <= input(5);
output(2, 6) <= input(6);
output(2, 7) <= input(7);
output(2, 8) <= input(8);
output(2, 9) <= input(9);
output(2, 10) <= input(10);
output(2, 11) <= input(11);
output(2, 12) <= input(12);
output(2, 13) <= input(13);
output(2, 14) <= input(14);
output(2, 15) <= input(15);
output(2, 16) <= input(0);
output(2, 17) <= input(1);
output(2, 18) <= input(2);
output(2, 19) <= input(3);
output(2, 20) <= input(4);
output(2, 21) <= input(5);
output(2, 22) <= input(6);
output(2, 23) <= input(7);
output(2, 24) <= input(8);
output(2, 25) <= input(9);
output(2, 26) <= input(10);
output(2, 27) <= input(11);
output(2, 28) <= input(12);
output(2, 29) <= input(13);
output(2, 30) <= input(14);
output(2, 31) <= input(15);
output(2, 32) <= input(0);
output(2, 33) <= input(1);
output(2, 34) <= input(2);
output(2, 35) <= input(3);
output(2, 36) <= input(4);
output(2, 37) <= input(5);
output(2, 38) <= input(6);
output(2, 39) <= input(7);
output(2, 40) <= input(8);
output(2, 41) <= input(9);
output(2, 42) <= input(10);
output(2, 43) <= input(11);
output(2, 44) <= input(12);
output(2, 45) <= input(13);
output(2, 46) <= input(14);
output(2, 47) <= input(15);
output(2, 48) <= input(0);
output(2, 49) <= input(1);
output(2, 50) <= input(2);
output(2, 51) <= input(3);
output(2, 52) <= input(4);
output(2, 53) <= input(5);
output(2, 54) <= input(6);
output(2, 55) <= input(7);
output(2, 56) <= input(8);
output(2, 57) <= input(9);
output(2, 58) <= input(10);
output(2, 59) <= input(11);
output(2, 60) <= input(12);
output(2, 61) <= input(13);
output(2, 62) <= input(14);
output(2, 63) <= input(15);
output(2, 64) <= input(0);
output(2, 65) <= input(1);
output(2, 66) <= input(2);
output(2, 67) <= input(3);
output(2, 68) <= input(4);
output(2, 69) <= input(5);
output(2, 70) <= input(6);
output(2, 71) <= input(7);
output(2, 72) <= input(8);
output(2, 73) <= input(9);
output(2, 74) <= input(10);
output(2, 75) <= input(11);
output(2, 76) <= input(12);
output(2, 77) <= input(13);
output(2, 78) <= input(14);
output(2, 79) <= input(15);
output(2, 80) <= input(0);
output(2, 81) <= input(1);
output(2, 82) <= input(2);
output(2, 83) <= input(3);
output(2, 84) <= input(4);
output(2, 85) <= input(5);
output(2, 86) <= input(6);
output(2, 87) <= input(7);
output(2, 88) <= input(8);
output(2, 89) <= input(9);
output(2, 90) <= input(10);
output(2, 91) <= input(11);
output(2, 92) <= input(12);
output(2, 93) <= input(13);
output(2, 94) <= input(14);
output(2, 95) <= input(15);
output(2, 96) <= input(0);
output(2, 97) <= input(1);
output(2, 98) <= input(2);
output(2, 99) <= input(3);
output(2, 100) <= input(4);
output(2, 101) <= input(5);
output(2, 102) <= input(6);
output(2, 103) <= input(7);
output(2, 104) <= input(8);
output(2, 105) <= input(9);
output(2, 106) <= input(10);
output(2, 107) <= input(11);
output(2, 108) <= input(12);
output(2, 109) <= input(13);
output(2, 110) <= input(14);
output(2, 111) <= input(15);
output(2, 112) <= input(0);
output(2, 113) <= input(1);
output(2, 114) <= input(2);
output(2, 115) <= input(3);
output(2, 116) <= input(4);
output(2, 117) <= input(5);
output(2, 118) <= input(6);
output(2, 119) <= input(7);
output(2, 120) <= input(8);
output(2, 121) <= input(9);
output(2, 122) <= input(10);
output(2, 123) <= input(11);
output(2, 124) <= input(12);
output(2, 125) <= input(13);
output(2, 126) <= input(14);
output(2, 127) <= input(15);
output(2, 128) <= input(0);
output(2, 129) <= input(1);
output(2, 130) <= input(2);
output(2, 131) <= input(3);
output(2, 132) <= input(4);
output(2, 133) <= input(5);
output(2, 134) <= input(6);
output(2, 135) <= input(7);
output(2, 136) <= input(8);
output(2, 137) <= input(9);
output(2, 138) <= input(10);
output(2, 139) <= input(11);
output(2, 140) <= input(12);
output(2, 141) <= input(13);
output(2, 142) <= input(14);
output(2, 143) <= input(15);
output(2, 144) <= input(0);
output(2, 145) <= input(1);
output(2, 146) <= input(2);
output(2, 147) <= input(3);
output(2, 148) <= input(4);
output(2, 149) <= input(5);
output(2, 150) <= input(6);
output(2, 151) <= input(7);
output(2, 152) <= input(8);
output(2, 153) <= input(9);
output(2, 154) <= input(10);
output(2, 155) <= input(11);
output(2, 156) <= input(12);
output(2, 157) <= input(13);
output(2, 158) <= input(14);
output(2, 159) <= input(15);
output(2, 160) <= input(0);
output(2, 161) <= input(1);
output(2, 162) <= input(2);
output(2, 163) <= input(3);
output(2, 164) <= input(4);
output(2, 165) <= input(5);
output(2, 166) <= input(6);
output(2, 167) <= input(7);
output(2, 168) <= input(8);
output(2, 169) <= input(9);
output(2, 170) <= input(10);
output(2, 171) <= input(11);
output(2, 172) <= input(12);
output(2, 173) <= input(13);
output(2, 174) <= input(14);
output(2, 175) <= input(15);
output(2, 176) <= input(0);
output(2, 177) <= input(1);
output(2, 178) <= input(2);
output(2, 179) <= input(3);
output(2, 180) <= input(4);
output(2, 181) <= input(5);
output(2, 182) <= input(6);
output(2, 183) <= input(7);
output(2, 184) <= input(8);
output(2, 185) <= input(9);
output(2, 186) <= input(10);
output(2, 187) <= input(11);
output(2, 188) <= input(12);
output(2, 189) <= input(13);
output(2, 190) <= input(14);
output(2, 191) <= input(15);
output(2, 192) <= input(0);
output(2, 193) <= input(1);
output(2, 194) <= input(2);
output(2, 195) <= input(3);
output(2, 196) <= input(4);
output(2, 197) <= input(5);
output(2, 198) <= input(6);
output(2, 199) <= input(7);
output(2, 200) <= input(8);
output(2, 201) <= input(9);
output(2, 202) <= input(10);
output(2, 203) <= input(11);
output(2, 204) <= input(12);
output(2, 205) <= input(13);
output(2, 206) <= input(14);
output(2, 207) <= input(15);
output(2, 208) <= input(0);
output(2, 209) <= input(1);
output(2, 210) <= input(2);
output(2, 211) <= input(3);
output(2, 212) <= input(4);
output(2, 213) <= input(5);
output(2, 214) <= input(6);
output(2, 215) <= input(7);
output(2, 216) <= input(8);
output(2, 217) <= input(9);
output(2, 218) <= input(10);
output(2, 219) <= input(11);
output(2, 220) <= input(12);
output(2, 221) <= input(13);
output(2, 222) <= input(14);
output(2, 223) <= input(15);
output(2, 224) <= input(0);
output(2, 225) <= input(1);
output(2, 226) <= input(2);
output(2, 227) <= input(3);
output(2, 228) <= input(4);
output(2, 229) <= input(5);
output(2, 230) <= input(6);
output(2, 231) <= input(7);
output(2, 232) <= input(8);
output(2, 233) <= input(9);
output(2, 234) <= input(10);
output(2, 235) <= input(11);
output(2, 236) <= input(12);
output(2, 237) <= input(13);
output(2, 238) <= input(14);
output(2, 239) <= input(15);
output(2, 240) <= input(0);
output(2, 241) <= input(1);
output(2, 242) <= input(2);
output(2, 243) <= input(3);
output(2, 244) <= input(4);
output(2, 245) <= input(5);
output(2, 246) <= input(6);
output(2, 247) <= input(7);
output(2, 248) <= input(8);
output(2, 249) <= input(9);
output(2, 250) <= input(10);
output(2, 251) <= input(11);
output(2, 252) <= input(12);
output(2, 253) <= input(13);
output(2, 254) <= input(14);
output(2, 255) <= input(15);
output(3, 0) <= input(17);
output(3, 1) <= input(18);
output(3, 2) <= input(19);
output(3, 3) <= input(20);
output(3, 4) <= input(21);
output(3, 5) <= input(22);
output(3, 6) <= input(23);
output(3, 7) <= input(24);
output(3, 8) <= input(25);
output(3, 9) <= input(26);
output(3, 10) <= input(27);
output(3, 11) <= input(28);
output(3, 12) <= input(29);
output(3, 13) <= input(30);
output(3, 14) <= input(31);
output(3, 15) <= input(33);
output(3, 16) <= input(17);
output(3, 17) <= input(18);
output(3, 18) <= input(19);
output(3, 19) <= input(20);
output(3, 20) <= input(21);
output(3, 21) <= input(22);
output(3, 22) <= input(23);
output(3, 23) <= input(24);
output(3, 24) <= input(25);
output(3, 25) <= input(26);
output(3, 26) <= input(27);
output(3, 27) <= input(28);
output(3, 28) <= input(29);
output(3, 29) <= input(30);
output(3, 30) <= input(31);
output(3, 31) <= input(33);
output(3, 32) <= input(17);
output(3, 33) <= input(18);
output(3, 34) <= input(19);
output(3, 35) <= input(20);
output(3, 36) <= input(21);
output(3, 37) <= input(22);
output(3, 38) <= input(23);
output(3, 39) <= input(24);
output(3, 40) <= input(25);
output(3, 41) <= input(26);
output(3, 42) <= input(27);
output(3, 43) <= input(28);
output(3, 44) <= input(29);
output(3, 45) <= input(30);
output(3, 46) <= input(31);
output(3, 47) <= input(33);
output(3, 48) <= input(17);
output(3, 49) <= input(18);
output(3, 50) <= input(19);
output(3, 51) <= input(20);
output(3, 52) <= input(21);
output(3, 53) <= input(22);
output(3, 54) <= input(23);
output(3, 55) <= input(24);
output(3, 56) <= input(25);
output(3, 57) <= input(26);
output(3, 58) <= input(27);
output(3, 59) <= input(28);
output(3, 60) <= input(29);
output(3, 61) <= input(30);
output(3, 62) <= input(31);
output(3, 63) <= input(33);
output(3, 64) <= input(17);
output(3, 65) <= input(18);
output(3, 66) <= input(19);
output(3, 67) <= input(20);
output(3, 68) <= input(21);
output(3, 69) <= input(22);
output(3, 70) <= input(23);
output(3, 71) <= input(24);
output(3, 72) <= input(25);
output(3, 73) <= input(26);
output(3, 74) <= input(27);
output(3, 75) <= input(28);
output(3, 76) <= input(29);
output(3, 77) <= input(30);
output(3, 78) <= input(31);
output(3, 79) <= input(33);
output(3, 80) <= input(17);
output(3, 81) <= input(18);
output(3, 82) <= input(19);
output(3, 83) <= input(20);
output(3, 84) <= input(21);
output(3, 85) <= input(22);
output(3, 86) <= input(23);
output(3, 87) <= input(24);
output(3, 88) <= input(25);
output(3, 89) <= input(26);
output(3, 90) <= input(27);
output(3, 91) <= input(28);
output(3, 92) <= input(29);
output(3, 93) <= input(30);
output(3, 94) <= input(31);
output(3, 95) <= input(33);
output(3, 96) <= input(17);
output(3, 97) <= input(18);
output(3, 98) <= input(19);
output(3, 99) <= input(20);
output(3, 100) <= input(21);
output(3, 101) <= input(22);
output(3, 102) <= input(23);
output(3, 103) <= input(24);
output(3, 104) <= input(25);
output(3, 105) <= input(26);
output(3, 106) <= input(27);
output(3, 107) <= input(28);
output(3, 108) <= input(29);
output(3, 109) <= input(30);
output(3, 110) <= input(31);
output(3, 111) <= input(33);
output(3, 112) <= input(17);
output(3, 113) <= input(18);
output(3, 114) <= input(19);
output(3, 115) <= input(20);
output(3, 116) <= input(21);
output(3, 117) <= input(22);
output(3, 118) <= input(23);
output(3, 119) <= input(24);
output(3, 120) <= input(25);
output(3, 121) <= input(26);
output(3, 122) <= input(27);
output(3, 123) <= input(28);
output(3, 124) <= input(29);
output(3, 125) <= input(30);
output(3, 126) <= input(31);
output(3, 127) <= input(33);
output(3, 128) <= input(17);
output(3, 129) <= input(18);
output(3, 130) <= input(19);
output(3, 131) <= input(20);
output(3, 132) <= input(21);
output(3, 133) <= input(22);
output(3, 134) <= input(23);
output(3, 135) <= input(24);
output(3, 136) <= input(25);
output(3, 137) <= input(26);
output(3, 138) <= input(27);
output(3, 139) <= input(28);
output(3, 140) <= input(29);
output(3, 141) <= input(30);
output(3, 142) <= input(31);
output(3, 143) <= input(33);
output(3, 144) <= input(17);
output(3, 145) <= input(18);
output(3, 146) <= input(19);
output(3, 147) <= input(20);
output(3, 148) <= input(21);
output(3, 149) <= input(22);
output(3, 150) <= input(23);
output(3, 151) <= input(24);
output(3, 152) <= input(25);
output(3, 153) <= input(26);
output(3, 154) <= input(27);
output(3, 155) <= input(28);
output(3, 156) <= input(29);
output(3, 157) <= input(30);
output(3, 158) <= input(31);
output(3, 159) <= input(33);
output(3, 160) <= input(17);
output(3, 161) <= input(18);
output(3, 162) <= input(19);
output(3, 163) <= input(20);
output(3, 164) <= input(21);
output(3, 165) <= input(22);
output(3, 166) <= input(23);
output(3, 167) <= input(24);
output(3, 168) <= input(25);
output(3, 169) <= input(26);
output(3, 170) <= input(27);
output(3, 171) <= input(28);
output(3, 172) <= input(29);
output(3, 173) <= input(30);
output(3, 174) <= input(31);
output(3, 175) <= input(33);
output(3, 176) <= input(17);
output(3, 177) <= input(18);
output(3, 178) <= input(19);
output(3, 179) <= input(20);
output(3, 180) <= input(21);
output(3, 181) <= input(22);
output(3, 182) <= input(23);
output(3, 183) <= input(24);
output(3, 184) <= input(25);
output(3, 185) <= input(26);
output(3, 186) <= input(27);
output(3, 187) <= input(28);
output(3, 188) <= input(29);
output(3, 189) <= input(30);
output(3, 190) <= input(31);
output(3, 191) <= input(33);
output(3, 192) <= input(17);
output(3, 193) <= input(18);
output(3, 194) <= input(19);
output(3, 195) <= input(20);
output(3, 196) <= input(21);
output(3, 197) <= input(22);
output(3, 198) <= input(23);
output(3, 199) <= input(24);
output(3, 200) <= input(25);
output(3, 201) <= input(26);
output(3, 202) <= input(27);
output(3, 203) <= input(28);
output(3, 204) <= input(29);
output(3, 205) <= input(30);
output(3, 206) <= input(31);
output(3, 207) <= input(33);
output(3, 208) <= input(17);
output(3, 209) <= input(18);
output(3, 210) <= input(19);
output(3, 211) <= input(20);
output(3, 212) <= input(21);
output(3, 213) <= input(22);
output(3, 214) <= input(23);
output(3, 215) <= input(24);
output(3, 216) <= input(25);
output(3, 217) <= input(26);
output(3, 218) <= input(27);
output(3, 219) <= input(28);
output(3, 220) <= input(29);
output(3, 221) <= input(30);
output(3, 222) <= input(31);
output(3, 223) <= input(33);
output(3, 224) <= input(17);
output(3, 225) <= input(18);
output(3, 226) <= input(19);
output(3, 227) <= input(20);
output(3, 228) <= input(21);
output(3, 229) <= input(22);
output(3, 230) <= input(23);
output(3, 231) <= input(24);
output(3, 232) <= input(25);
output(3, 233) <= input(26);
output(3, 234) <= input(27);
output(3, 235) <= input(28);
output(3, 236) <= input(29);
output(3, 237) <= input(30);
output(3, 238) <= input(31);
output(3, 239) <= input(33);
output(3, 240) <= input(17);
output(3, 241) <= input(18);
output(3, 242) <= input(19);
output(3, 243) <= input(20);
output(3, 244) <= input(21);
output(3, 245) <= input(22);
output(3, 246) <= input(23);
output(3, 247) <= input(24);
output(3, 248) <= input(25);
output(3, 249) <= input(26);
output(3, 250) <= input(27);
output(3, 251) <= input(28);
output(3, 252) <= input(29);
output(3, 253) <= input(30);
output(3, 254) <= input(31);
output(3, 255) <= input(33);
output(4, 0) <= input(17);
output(4, 1) <= input(18);
output(4, 2) <= input(19);
output(4, 3) <= input(20);
output(4, 4) <= input(21);
output(4, 5) <= input(22);
output(4, 6) <= input(23);
output(4, 7) <= input(24);
output(4, 8) <= input(25);
output(4, 9) <= input(26);
output(4, 10) <= input(27);
output(4, 11) <= input(28);
output(4, 12) <= input(29);
output(4, 13) <= input(30);
output(4, 14) <= input(31);
output(4, 15) <= input(33);
output(4, 16) <= input(17);
output(4, 17) <= input(18);
output(4, 18) <= input(19);
output(4, 19) <= input(20);
output(4, 20) <= input(21);
output(4, 21) <= input(22);
output(4, 22) <= input(23);
output(4, 23) <= input(24);
output(4, 24) <= input(25);
output(4, 25) <= input(26);
output(4, 26) <= input(27);
output(4, 27) <= input(28);
output(4, 28) <= input(29);
output(4, 29) <= input(30);
output(4, 30) <= input(31);
output(4, 31) <= input(33);
output(4, 32) <= input(17);
output(4, 33) <= input(18);
output(4, 34) <= input(19);
output(4, 35) <= input(20);
output(4, 36) <= input(21);
output(4, 37) <= input(22);
output(4, 38) <= input(23);
output(4, 39) <= input(24);
output(4, 40) <= input(25);
output(4, 41) <= input(26);
output(4, 42) <= input(27);
output(4, 43) <= input(28);
output(4, 44) <= input(29);
output(4, 45) <= input(30);
output(4, 46) <= input(31);
output(4, 47) <= input(33);
output(4, 48) <= input(17);
output(4, 49) <= input(18);
output(4, 50) <= input(19);
output(4, 51) <= input(20);
output(4, 52) <= input(21);
output(4, 53) <= input(22);
output(4, 54) <= input(23);
output(4, 55) <= input(24);
output(4, 56) <= input(25);
output(4, 57) <= input(26);
output(4, 58) <= input(27);
output(4, 59) <= input(28);
output(4, 60) <= input(29);
output(4, 61) <= input(30);
output(4, 62) <= input(31);
output(4, 63) <= input(33);
output(4, 64) <= input(17);
output(4, 65) <= input(18);
output(4, 66) <= input(19);
output(4, 67) <= input(20);
output(4, 68) <= input(21);
output(4, 69) <= input(22);
output(4, 70) <= input(23);
output(4, 71) <= input(24);
output(4, 72) <= input(25);
output(4, 73) <= input(26);
output(4, 74) <= input(27);
output(4, 75) <= input(28);
output(4, 76) <= input(29);
output(4, 77) <= input(30);
output(4, 78) <= input(31);
output(4, 79) <= input(33);
output(4, 80) <= input(17);
output(4, 81) <= input(18);
output(4, 82) <= input(19);
output(4, 83) <= input(20);
output(4, 84) <= input(21);
output(4, 85) <= input(22);
output(4, 86) <= input(23);
output(4, 87) <= input(24);
output(4, 88) <= input(25);
output(4, 89) <= input(26);
output(4, 90) <= input(27);
output(4, 91) <= input(28);
output(4, 92) <= input(29);
output(4, 93) <= input(30);
output(4, 94) <= input(31);
output(4, 95) <= input(33);
output(4, 96) <= input(17);
output(4, 97) <= input(18);
output(4, 98) <= input(19);
output(4, 99) <= input(20);
output(4, 100) <= input(21);
output(4, 101) <= input(22);
output(4, 102) <= input(23);
output(4, 103) <= input(24);
output(4, 104) <= input(25);
output(4, 105) <= input(26);
output(4, 106) <= input(27);
output(4, 107) <= input(28);
output(4, 108) <= input(29);
output(4, 109) <= input(30);
output(4, 110) <= input(31);
output(4, 111) <= input(33);
output(4, 112) <= input(17);
output(4, 113) <= input(18);
output(4, 114) <= input(19);
output(4, 115) <= input(20);
output(4, 116) <= input(21);
output(4, 117) <= input(22);
output(4, 118) <= input(23);
output(4, 119) <= input(24);
output(4, 120) <= input(25);
output(4, 121) <= input(26);
output(4, 122) <= input(27);
output(4, 123) <= input(28);
output(4, 124) <= input(29);
output(4, 125) <= input(30);
output(4, 126) <= input(31);
output(4, 127) <= input(33);
output(4, 128) <= input(17);
output(4, 129) <= input(18);
output(4, 130) <= input(19);
output(4, 131) <= input(20);
output(4, 132) <= input(21);
output(4, 133) <= input(22);
output(4, 134) <= input(23);
output(4, 135) <= input(24);
output(4, 136) <= input(25);
output(4, 137) <= input(26);
output(4, 138) <= input(27);
output(4, 139) <= input(28);
output(4, 140) <= input(29);
output(4, 141) <= input(30);
output(4, 142) <= input(31);
output(4, 143) <= input(33);
output(4, 144) <= input(17);
output(4, 145) <= input(18);
output(4, 146) <= input(19);
output(4, 147) <= input(20);
output(4, 148) <= input(21);
output(4, 149) <= input(22);
output(4, 150) <= input(23);
output(4, 151) <= input(24);
output(4, 152) <= input(25);
output(4, 153) <= input(26);
output(4, 154) <= input(27);
output(4, 155) <= input(28);
output(4, 156) <= input(29);
output(4, 157) <= input(30);
output(4, 158) <= input(31);
output(4, 159) <= input(33);
output(4, 160) <= input(17);
output(4, 161) <= input(18);
output(4, 162) <= input(19);
output(4, 163) <= input(20);
output(4, 164) <= input(21);
output(4, 165) <= input(22);
output(4, 166) <= input(23);
output(4, 167) <= input(24);
output(4, 168) <= input(25);
output(4, 169) <= input(26);
output(4, 170) <= input(27);
output(4, 171) <= input(28);
output(4, 172) <= input(29);
output(4, 173) <= input(30);
output(4, 174) <= input(31);
output(4, 175) <= input(33);
output(4, 176) <= input(17);
output(4, 177) <= input(18);
output(4, 178) <= input(19);
output(4, 179) <= input(20);
output(4, 180) <= input(21);
output(4, 181) <= input(22);
output(4, 182) <= input(23);
output(4, 183) <= input(24);
output(4, 184) <= input(25);
output(4, 185) <= input(26);
output(4, 186) <= input(27);
output(4, 187) <= input(28);
output(4, 188) <= input(29);
output(4, 189) <= input(30);
output(4, 190) <= input(31);
output(4, 191) <= input(33);
output(4, 192) <= input(17);
output(4, 193) <= input(18);
output(4, 194) <= input(19);
output(4, 195) <= input(20);
output(4, 196) <= input(21);
output(4, 197) <= input(22);
output(4, 198) <= input(23);
output(4, 199) <= input(24);
output(4, 200) <= input(25);
output(4, 201) <= input(26);
output(4, 202) <= input(27);
output(4, 203) <= input(28);
output(4, 204) <= input(29);
output(4, 205) <= input(30);
output(4, 206) <= input(31);
output(4, 207) <= input(33);
output(4, 208) <= input(17);
output(4, 209) <= input(18);
output(4, 210) <= input(19);
output(4, 211) <= input(20);
output(4, 212) <= input(21);
output(4, 213) <= input(22);
output(4, 214) <= input(23);
output(4, 215) <= input(24);
output(4, 216) <= input(25);
output(4, 217) <= input(26);
output(4, 218) <= input(27);
output(4, 219) <= input(28);
output(4, 220) <= input(29);
output(4, 221) <= input(30);
output(4, 222) <= input(31);
output(4, 223) <= input(33);
output(4, 224) <= input(17);
output(4, 225) <= input(18);
output(4, 226) <= input(19);
output(4, 227) <= input(20);
output(4, 228) <= input(21);
output(4, 229) <= input(22);
output(4, 230) <= input(23);
output(4, 231) <= input(24);
output(4, 232) <= input(25);
output(4, 233) <= input(26);
output(4, 234) <= input(27);
output(4, 235) <= input(28);
output(4, 236) <= input(29);
output(4, 237) <= input(30);
output(4, 238) <= input(31);
output(4, 239) <= input(33);
output(4, 240) <= input(1);
output(4, 241) <= input(2);
output(4, 242) <= input(3);
output(4, 243) <= input(4);
output(4, 244) <= input(5);
output(4, 245) <= input(6);
output(4, 246) <= input(7);
output(4, 247) <= input(8);
output(4, 248) <= input(9);
output(4, 249) <= input(10);
output(4, 250) <= input(11);
output(4, 251) <= input(12);
output(4, 252) <= input(13);
output(4, 253) <= input(14);
output(4, 254) <= input(15);
output(4, 255) <= input(34);
output(5, 0) <= input(17);
output(5, 1) <= input(18);
output(5, 2) <= input(19);
output(5, 3) <= input(20);
output(5, 4) <= input(21);
output(5, 5) <= input(22);
output(5, 6) <= input(23);
output(5, 7) <= input(24);
output(5, 8) <= input(25);
output(5, 9) <= input(26);
output(5, 10) <= input(27);
output(5, 11) <= input(28);
output(5, 12) <= input(29);
output(5, 13) <= input(30);
output(5, 14) <= input(31);
output(5, 15) <= input(33);
output(5, 16) <= input(17);
output(5, 17) <= input(18);
output(5, 18) <= input(19);
output(5, 19) <= input(20);
output(5, 20) <= input(21);
output(5, 21) <= input(22);
output(5, 22) <= input(23);
output(5, 23) <= input(24);
output(5, 24) <= input(25);
output(5, 25) <= input(26);
output(5, 26) <= input(27);
output(5, 27) <= input(28);
output(5, 28) <= input(29);
output(5, 29) <= input(30);
output(5, 30) <= input(31);
output(5, 31) <= input(33);
output(5, 32) <= input(17);
output(5, 33) <= input(18);
output(5, 34) <= input(19);
output(5, 35) <= input(20);
output(5, 36) <= input(21);
output(5, 37) <= input(22);
output(5, 38) <= input(23);
output(5, 39) <= input(24);
output(5, 40) <= input(25);
output(5, 41) <= input(26);
output(5, 42) <= input(27);
output(5, 43) <= input(28);
output(5, 44) <= input(29);
output(5, 45) <= input(30);
output(5, 46) <= input(31);
output(5, 47) <= input(33);
output(5, 48) <= input(17);
output(5, 49) <= input(18);
output(5, 50) <= input(19);
output(5, 51) <= input(20);
output(5, 52) <= input(21);
output(5, 53) <= input(22);
output(5, 54) <= input(23);
output(5, 55) <= input(24);
output(5, 56) <= input(25);
output(5, 57) <= input(26);
output(5, 58) <= input(27);
output(5, 59) <= input(28);
output(5, 60) <= input(29);
output(5, 61) <= input(30);
output(5, 62) <= input(31);
output(5, 63) <= input(33);
output(5, 64) <= input(17);
output(5, 65) <= input(18);
output(5, 66) <= input(19);
output(5, 67) <= input(20);
output(5, 68) <= input(21);
output(5, 69) <= input(22);
output(5, 70) <= input(23);
output(5, 71) <= input(24);
output(5, 72) <= input(25);
output(5, 73) <= input(26);
output(5, 74) <= input(27);
output(5, 75) <= input(28);
output(5, 76) <= input(29);
output(5, 77) <= input(30);
output(5, 78) <= input(31);
output(5, 79) <= input(33);
output(5, 80) <= input(17);
output(5, 81) <= input(18);
output(5, 82) <= input(19);
output(5, 83) <= input(20);
output(5, 84) <= input(21);
output(5, 85) <= input(22);
output(5, 86) <= input(23);
output(5, 87) <= input(24);
output(5, 88) <= input(25);
output(5, 89) <= input(26);
output(5, 90) <= input(27);
output(5, 91) <= input(28);
output(5, 92) <= input(29);
output(5, 93) <= input(30);
output(5, 94) <= input(31);
output(5, 95) <= input(33);
output(5, 96) <= input(17);
output(5, 97) <= input(18);
output(5, 98) <= input(19);
output(5, 99) <= input(20);
output(5, 100) <= input(21);
output(5, 101) <= input(22);
output(5, 102) <= input(23);
output(5, 103) <= input(24);
output(5, 104) <= input(25);
output(5, 105) <= input(26);
output(5, 106) <= input(27);
output(5, 107) <= input(28);
output(5, 108) <= input(29);
output(5, 109) <= input(30);
output(5, 110) <= input(31);
output(5, 111) <= input(33);
output(5, 112) <= input(1);
output(5, 113) <= input(2);
output(5, 114) <= input(3);
output(5, 115) <= input(4);
output(5, 116) <= input(5);
output(5, 117) <= input(6);
output(5, 118) <= input(7);
output(5, 119) <= input(8);
output(5, 120) <= input(9);
output(5, 121) <= input(10);
output(5, 122) <= input(11);
output(5, 123) <= input(12);
output(5, 124) <= input(13);
output(5, 125) <= input(14);
output(5, 126) <= input(15);
output(5, 127) <= input(34);
output(5, 128) <= input(1);
output(5, 129) <= input(2);
output(5, 130) <= input(3);
output(5, 131) <= input(4);
output(5, 132) <= input(5);
output(5, 133) <= input(6);
output(5, 134) <= input(7);
output(5, 135) <= input(8);
output(5, 136) <= input(9);
output(5, 137) <= input(10);
output(5, 138) <= input(11);
output(5, 139) <= input(12);
output(5, 140) <= input(13);
output(5, 141) <= input(14);
output(5, 142) <= input(15);
output(5, 143) <= input(34);
output(5, 144) <= input(1);
output(5, 145) <= input(2);
output(5, 146) <= input(3);
output(5, 147) <= input(4);
output(5, 148) <= input(5);
output(5, 149) <= input(6);
output(5, 150) <= input(7);
output(5, 151) <= input(8);
output(5, 152) <= input(9);
output(5, 153) <= input(10);
output(5, 154) <= input(11);
output(5, 155) <= input(12);
output(5, 156) <= input(13);
output(5, 157) <= input(14);
output(5, 158) <= input(15);
output(5, 159) <= input(34);
output(5, 160) <= input(1);
output(5, 161) <= input(2);
output(5, 162) <= input(3);
output(5, 163) <= input(4);
output(5, 164) <= input(5);
output(5, 165) <= input(6);
output(5, 166) <= input(7);
output(5, 167) <= input(8);
output(5, 168) <= input(9);
output(5, 169) <= input(10);
output(5, 170) <= input(11);
output(5, 171) <= input(12);
output(5, 172) <= input(13);
output(5, 173) <= input(14);
output(5, 174) <= input(15);
output(5, 175) <= input(34);
output(5, 176) <= input(1);
output(5, 177) <= input(2);
output(5, 178) <= input(3);
output(5, 179) <= input(4);
output(5, 180) <= input(5);
output(5, 181) <= input(6);
output(5, 182) <= input(7);
output(5, 183) <= input(8);
output(5, 184) <= input(9);
output(5, 185) <= input(10);
output(5, 186) <= input(11);
output(5, 187) <= input(12);
output(5, 188) <= input(13);
output(5, 189) <= input(14);
output(5, 190) <= input(15);
output(5, 191) <= input(34);
output(5, 192) <= input(1);
output(5, 193) <= input(2);
output(5, 194) <= input(3);
output(5, 195) <= input(4);
output(5, 196) <= input(5);
output(5, 197) <= input(6);
output(5, 198) <= input(7);
output(5, 199) <= input(8);
output(5, 200) <= input(9);
output(5, 201) <= input(10);
output(5, 202) <= input(11);
output(5, 203) <= input(12);
output(5, 204) <= input(13);
output(5, 205) <= input(14);
output(5, 206) <= input(15);
output(5, 207) <= input(34);
output(5, 208) <= input(1);
output(5, 209) <= input(2);
output(5, 210) <= input(3);
output(5, 211) <= input(4);
output(5, 212) <= input(5);
output(5, 213) <= input(6);
output(5, 214) <= input(7);
output(5, 215) <= input(8);
output(5, 216) <= input(9);
output(5, 217) <= input(10);
output(5, 218) <= input(11);
output(5, 219) <= input(12);
output(5, 220) <= input(13);
output(5, 221) <= input(14);
output(5, 222) <= input(15);
output(5, 223) <= input(34);
output(5, 224) <= input(1);
output(5, 225) <= input(2);
output(5, 226) <= input(3);
output(5, 227) <= input(4);
output(5, 228) <= input(5);
output(5, 229) <= input(6);
output(5, 230) <= input(7);
output(5, 231) <= input(8);
output(5, 232) <= input(9);
output(5, 233) <= input(10);
output(5, 234) <= input(11);
output(5, 235) <= input(12);
output(5, 236) <= input(13);
output(5, 237) <= input(14);
output(5, 238) <= input(15);
output(5, 239) <= input(34);
output(5, 240) <= input(18);
output(5, 241) <= input(19);
output(5, 242) <= input(20);
output(5, 243) <= input(21);
output(5, 244) <= input(22);
output(5, 245) <= input(23);
output(5, 246) <= input(24);
output(5, 247) <= input(25);
output(5, 248) <= input(26);
output(5, 249) <= input(27);
output(5, 250) <= input(28);
output(5, 251) <= input(29);
output(5, 252) <= input(30);
output(5, 253) <= input(31);
output(5, 254) <= input(33);
output(5, 255) <= input(35);
output(6, 0) <= input(17);
output(6, 1) <= input(18);
output(6, 2) <= input(19);
output(6, 3) <= input(20);
output(6, 4) <= input(21);
output(6, 5) <= input(22);
output(6, 6) <= input(23);
output(6, 7) <= input(24);
output(6, 8) <= input(25);
output(6, 9) <= input(26);
output(6, 10) <= input(27);
output(6, 11) <= input(28);
output(6, 12) <= input(29);
output(6, 13) <= input(30);
output(6, 14) <= input(31);
output(6, 15) <= input(33);
output(6, 16) <= input(17);
output(6, 17) <= input(18);
output(6, 18) <= input(19);
output(6, 19) <= input(20);
output(6, 20) <= input(21);
output(6, 21) <= input(22);
output(6, 22) <= input(23);
output(6, 23) <= input(24);
output(6, 24) <= input(25);
output(6, 25) <= input(26);
output(6, 26) <= input(27);
output(6, 27) <= input(28);
output(6, 28) <= input(29);
output(6, 29) <= input(30);
output(6, 30) <= input(31);
output(6, 31) <= input(33);
output(6, 32) <= input(17);
output(6, 33) <= input(18);
output(6, 34) <= input(19);
output(6, 35) <= input(20);
output(6, 36) <= input(21);
output(6, 37) <= input(22);
output(6, 38) <= input(23);
output(6, 39) <= input(24);
output(6, 40) <= input(25);
output(6, 41) <= input(26);
output(6, 42) <= input(27);
output(6, 43) <= input(28);
output(6, 44) <= input(29);
output(6, 45) <= input(30);
output(6, 46) <= input(31);
output(6, 47) <= input(33);
output(6, 48) <= input(17);
output(6, 49) <= input(18);
output(6, 50) <= input(19);
output(6, 51) <= input(20);
output(6, 52) <= input(21);
output(6, 53) <= input(22);
output(6, 54) <= input(23);
output(6, 55) <= input(24);
output(6, 56) <= input(25);
output(6, 57) <= input(26);
output(6, 58) <= input(27);
output(6, 59) <= input(28);
output(6, 60) <= input(29);
output(6, 61) <= input(30);
output(6, 62) <= input(31);
output(6, 63) <= input(33);
output(6, 64) <= input(17);
output(6, 65) <= input(18);
output(6, 66) <= input(19);
output(6, 67) <= input(20);
output(6, 68) <= input(21);
output(6, 69) <= input(22);
output(6, 70) <= input(23);
output(6, 71) <= input(24);
output(6, 72) <= input(25);
output(6, 73) <= input(26);
output(6, 74) <= input(27);
output(6, 75) <= input(28);
output(6, 76) <= input(29);
output(6, 77) <= input(30);
output(6, 78) <= input(31);
output(6, 79) <= input(33);
output(6, 80) <= input(1);
output(6, 81) <= input(2);
output(6, 82) <= input(3);
output(6, 83) <= input(4);
output(6, 84) <= input(5);
output(6, 85) <= input(6);
output(6, 86) <= input(7);
output(6, 87) <= input(8);
output(6, 88) <= input(9);
output(6, 89) <= input(10);
output(6, 90) <= input(11);
output(6, 91) <= input(12);
output(6, 92) <= input(13);
output(6, 93) <= input(14);
output(6, 94) <= input(15);
output(6, 95) <= input(34);
output(6, 96) <= input(1);
output(6, 97) <= input(2);
output(6, 98) <= input(3);
output(6, 99) <= input(4);
output(6, 100) <= input(5);
output(6, 101) <= input(6);
output(6, 102) <= input(7);
output(6, 103) <= input(8);
output(6, 104) <= input(9);
output(6, 105) <= input(10);
output(6, 106) <= input(11);
output(6, 107) <= input(12);
output(6, 108) <= input(13);
output(6, 109) <= input(14);
output(6, 110) <= input(15);
output(6, 111) <= input(34);
output(6, 112) <= input(1);
output(6, 113) <= input(2);
output(6, 114) <= input(3);
output(6, 115) <= input(4);
output(6, 116) <= input(5);
output(6, 117) <= input(6);
output(6, 118) <= input(7);
output(6, 119) <= input(8);
output(6, 120) <= input(9);
output(6, 121) <= input(10);
output(6, 122) <= input(11);
output(6, 123) <= input(12);
output(6, 124) <= input(13);
output(6, 125) <= input(14);
output(6, 126) <= input(15);
output(6, 127) <= input(34);
output(6, 128) <= input(1);
output(6, 129) <= input(2);
output(6, 130) <= input(3);
output(6, 131) <= input(4);
output(6, 132) <= input(5);
output(6, 133) <= input(6);
output(6, 134) <= input(7);
output(6, 135) <= input(8);
output(6, 136) <= input(9);
output(6, 137) <= input(10);
output(6, 138) <= input(11);
output(6, 139) <= input(12);
output(6, 140) <= input(13);
output(6, 141) <= input(14);
output(6, 142) <= input(15);
output(6, 143) <= input(34);
output(6, 144) <= input(1);
output(6, 145) <= input(2);
output(6, 146) <= input(3);
output(6, 147) <= input(4);
output(6, 148) <= input(5);
output(6, 149) <= input(6);
output(6, 150) <= input(7);
output(6, 151) <= input(8);
output(6, 152) <= input(9);
output(6, 153) <= input(10);
output(6, 154) <= input(11);
output(6, 155) <= input(12);
output(6, 156) <= input(13);
output(6, 157) <= input(14);
output(6, 158) <= input(15);
output(6, 159) <= input(34);
output(6, 160) <= input(18);
output(6, 161) <= input(19);
output(6, 162) <= input(20);
output(6, 163) <= input(21);
output(6, 164) <= input(22);
output(6, 165) <= input(23);
output(6, 166) <= input(24);
output(6, 167) <= input(25);
output(6, 168) <= input(26);
output(6, 169) <= input(27);
output(6, 170) <= input(28);
output(6, 171) <= input(29);
output(6, 172) <= input(30);
output(6, 173) <= input(31);
output(6, 174) <= input(33);
output(6, 175) <= input(35);
output(6, 176) <= input(18);
output(6, 177) <= input(19);
output(6, 178) <= input(20);
output(6, 179) <= input(21);
output(6, 180) <= input(22);
output(6, 181) <= input(23);
output(6, 182) <= input(24);
output(6, 183) <= input(25);
output(6, 184) <= input(26);
output(6, 185) <= input(27);
output(6, 186) <= input(28);
output(6, 187) <= input(29);
output(6, 188) <= input(30);
output(6, 189) <= input(31);
output(6, 190) <= input(33);
output(6, 191) <= input(35);
output(6, 192) <= input(18);
output(6, 193) <= input(19);
output(6, 194) <= input(20);
output(6, 195) <= input(21);
output(6, 196) <= input(22);
output(6, 197) <= input(23);
output(6, 198) <= input(24);
output(6, 199) <= input(25);
output(6, 200) <= input(26);
output(6, 201) <= input(27);
output(6, 202) <= input(28);
output(6, 203) <= input(29);
output(6, 204) <= input(30);
output(6, 205) <= input(31);
output(6, 206) <= input(33);
output(6, 207) <= input(35);
output(6, 208) <= input(18);
output(6, 209) <= input(19);
output(6, 210) <= input(20);
output(6, 211) <= input(21);
output(6, 212) <= input(22);
output(6, 213) <= input(23);
output(6, 214) <= input(24);
output(6, 215) <= input(25);
output(6, 216) <= input(26);
output(6, 217) <= input(27);
output(6, 218) <= input(28);
output(6, 219) <= input(29);
output(6, 220) <= input(30);
output(6, 221) <= input(31);
output(6, 222) <= input(33);
output(6, 223) <= input(35);
output(6, 224) <= input(18);
output(6, 225) <= input(19);
output(6, 226) <= input(20);
output(6, 227) <= input(21);
output(6, 228) <= input(22);
output(6, 229) <= input(23);
output(6, 230) <= input(24);
output(6, 231) <= input(25);
output(6, 232) <= input(26);
output(6, 233) <= input(27);
output(6, 234) <= input(28);
output(6, 235) <= input(29);
output(6, 236) <= input(30);
output(6, 237) <= input(31);
output(6, 238) <= input(33);
output(6, 239) <= input(35);
output(6, 240) <= input(2);
output(6, 241) <= input(3);
output(6, 242) <= input(4);
output(6, 243) <= input(5);
output(6, 244) <= input(6);
output(6, 245) <= input(7);
output(6, 246) <= input(8);
output(6, 247) <= input(9);
output(6, 248) <= input(10);
output(6, 249) <= input(11);
output(6, 250) <= input(12);
output(6, 251) <= input(13);
output(6, 252) <= input(14);
output(6, 253) <= input(15);
output(6, 254) <= input(34);
output(6, 255) <= input(36);
output(7, 0) <= input(17);
output(7, 1) <= input(18);
output(7, 2) <= input(19);
output(7, 3) <= input(20);
output(7, 4) <= input(21);
output(7, 5) <= input(22);
output(7, 6) <= input(23);
output(7, 7) <= input(24);
output(7, 8) <= input(25);
output(7, 9) <= input(26);
output(7, 10) <= input(27);
output(7, 11) <= input(28);
output(7, 12) <= input(29);
output(7, 13) <= input(30);
output(7, 14) <= input(31);
output(7, 15) <= input(33);
output(7, 16) <= input(17);
output(7, 17) <= input(18);
output(7, 18) <= input(19);
output(7, 19) <= input(20);
output(7, 20) <= input(21);
output(7, 21) <= input(22);
output(7, 22) <= input(23);
output(7, 23) <= input(24);
output(7, 24) <= input(25);
output(7, 25) <= input(26);
output(7, 26) <= input(27);
output(7, 27) <= input(28);
output(7, 28) <= input(29);
output(7, 29) <= input(30);
output(7, 30) <= input(31);
output(7, 31) <= input(33);
output(7, 32) <= input(17);
output(7, 33) <= input(18);
output(7, 34) <= input(19);
output(7, 35) <= input(20);
output(7, 36) <= input(21);
output(7, 37) <= input(22);
output(7, 38) <= input(23);
output(7, 39) <= input(24);
output(7, 40) <= input(25);
output(7, 41) <= input(26);
output(7, 42) <= input(27);
output(7, 43) <= input(28);
output(7, 44) <= input(29);
output(7, 45) <= input(30);
output(7, 46) <= input(31);
output(7, 47) <= input(33);
output(7, 48) <= input(1);
output(7, 49) <= input(2);
output(7, 50) <= input(3);
output(7, 51) <= input(4);
output(7, 52) <= input(5);
output(7, 53) <= input(6);
output(7, 54) <= input(7);
output(7, 55) <= input(8);
output(7, 56) <= input(9);
output(7, 57) <= input(10);
output(7, 58) <= input(11);
output(7, 59) <= input(12);
output(7, 60) <= input(13);
output(7, 61) <= input(14);
output(7, 62) <= input(15);
output(7, 63) <= input(34);
output(7, 64) <= input(1);
output(7, 65) <= input(2);
output(7, 66) <= input(3);
output(7, 67) <= input(4);
output(7, 68) <= input(5);
output(7, 69) <= input(6);
output(7, 70) <= input(7);
output(7, 71) <= input(8);
output(7, 72) <= input(9);
output(7, 73) <= input(10);
output(7, 74) <= input(11);
output(7, 75) <= input(12);
output(7, 76) <= input(13);
output(7, 77) <= input(14);
output(7, 78) <= input(15);
output(7, 79) <= input(34);
output(7, 80) <= input(1);
output(7, 81) <= input(2);
output(7, 82) <= input(3);
output(7, 83) <= input(4);
output(7, 84) <= input(5);
output(7, 85) <= input(6);
output(7, 86) <= input(7);
output(7, 87) <= input(8);
output(7, 88) <= input(9);
output(7, 89) <= input(10);
output(7, 90) <= input(11);
output(7, 91) <= input(12);
output(7, 92) <= input(13);
output(7, 93) <= input(14);
output(7, 94) <= input(15);
output(7, 95) <= input(34);
output(7, 96) <= input(1);
output(7, 97) <= input(2);
output(7, 98) <= input(3);
output(7, 99) <= input(4);
output(7, 100) <= input(5);
output(7, 101) <= input(6);
output(7, 102) <= input(7);
output(7, 103) <= input(8);
output(7, 104) <= input(9);
output(7, 105) <= input(10);
output(7, 106) <= input(11);
output(7, 107) <= input(12);
output(7, 108) <= input(13);
output(7, 109) <= input(14);
output(7, 110) <= input(15);
output(7, 111) <= input(34);
output(7, 112) <= input(18);
output(7, 113) <= input(19);
output(7, 114) <= input(20);
output(7, 115) <= input(21);
output(7, 116) <= input(22);
output(7, 117) <= input(23);
output(7, 118) <= input(24);
output(7, 119) <= input(25);
output(7, 120) <= input(26);
output(7, 121) <= input(27);
output(7, 122) <= input(28);
output(7, 123) <= input(29);
output(7, 124) <= input(30);
output(7, 125) <= input(31);
output(7, 126) <= input(33);
output(7, 127) <= input(35);
output(7, 128) <= input(18);
output(7, 129) <= input(19);
output(7, 130) <= input(20);
output(7, 131) <= input(21);
output(7, 132) <= input(22);
output(7, 133) <= input(23);
output(7, 134) <= input(24);
output(7, 135) <= input(25);
output(7, 136) <= input(26);
output(7, 137) <= input(27);
output(7, 138) <= input(28);
output(7, 139) <= input(29);
output(7, 140) <= input(30);
output(7, 141) <= input(31);
output(7, 142) <= input(33);
output(7, 143) <= input(35);
output(7, 144) <= input(18);
output(7, 145) <= input(19);
output(7, 146) <= input(20);
output(7, 147) <= input(21);
output(7, 148) <= input(22);
output(7, 149) <= input(23);
output(7, 150) <= input(24);
output(7, 151) <= input(25);
output(7, 152) <= input(26);
output(7, 153) <= input(27);
output(7, 154) <= input(28);
output(7, 155) <= input(29);
output(7, 156) <= input(30);
output(7, 157) <= input(31);
output(7, 158) <= input(33);
output(7, 159) <= input(35);
output(7, 160) <= input(18);
output(7, 161) <= input(19);
output(7, 162) <= input(20);
output(7, 163) <= input(21);
output(7, 164) <= input(22);
output(7, 165) <= input(23);
output(7, 166) <= input(24);
output(7, 167) <= input(25);
output(7, 168) <= input(26);
output(7, 169) <= input(27);
output(7, 170) <= input(28);
output(7, 171) <= input(29);
output(7, 172) <= input(30);
output(7, 173) <= input(31);
output(7, 174) <= input(33);
output(7, 175) <= input(35);
output(7, 176) <= input(2);
output(7, 177) <= input(3);
output(7, 178) <= input(4);
output(7, 179) <= input(5);
output(7, 180) <= input(6);
output(7, 181) <= input(7);
output(7, 182) <= input(8);
output(7, 183) <= input(9);
output(7, 184) <= input(10);
output(7, 185) <= input(11);
output(7, 186) <= input(12);
output(7, 187) <= input(13);
output(7, 188) <= input(14);
output(7, 189) <= input(15);
output(7, 190) <= input(34);
output(7, 191) <= input(36);
output(7, 192) <= input(2);
output(7, 193) <= input(3);
output(7, 194) <= input(4);
output(7, 195) <= input(5);
output(7, 196) <= input(6);
output(7, 197) <= input(7);
output(7, 198) <= input(8);
output(7, 199) <= input(9);
output(7, 200) <= input(10);
output(7, 201) <= input(11);
output(7, 202) <= input(12);
output(7, 203) <= input(13);
output(7, 204) <= input(14);
output(7, 205) <= input(15);
output(7, 206) <= input(34);
output(7, 207) <= input(36);
output(7, 208) <= input(2);
output(7, 209) <= input(3);
output(7, 210) <= input(4);
output(7, 211) <= input(5);
output(7, 212) <= input(6);
output(7, 213) <= input(7);
output(7, 214) <= input(8);
output(7, 215) <= input(9);
output(7, 216) <= input(10);
output(7, 217) <= input(11);
output(7, 218) <= input(12);
output(7, 219) <= input(13);
output(7, 220) <= input(14);
output(7, 221) <= input(15);
output(7, 222) <= input(34);
output(7, 223) <= input(36);
output(7, 224) <= input(2);
output(7, 225) <= input(3);
output(7, 226) <= input(4);
output(7, 227) <= input(5);
output(7, 228) <= input(6);
output(7, 229) <= input(7);
output(7, 230) <= input(8);
output(7, 231) <= input(9);
output(7, 232) <= input(10);
output(7, 233) <= input(11);
output(7, 234) <= input(12);
output(7, 235) <= input(13);
output(7, 236) <= input(14);
output(7, 237) <= input(15);
output(7, 238) <= input(34);
output(7, 239) <= input(36);
output(7, 240) <= input(19);
output(7, 241) <= input(20);
output(7, 242) <= input(21);
output(7, 243) <= input(22);
output(7, 244) <= input(23);
output(7, 245) <= input(24);
output(7, 246) <= input(25);
output(7, 247) <= input(26);
output(7, 248) <= input(27);
output(7, 249) <= input(28);
output(7, 250) <= input(29);
output(7, 251) <= input(30);
output(7, 252) <= input(31);
output(7, 253) <= input(33);
output(7, 254) <= input(35);
output(7, 255) <= input(37);
when "1110" =>
output(0, 0) <= input(0);
output(0, 1) <= input(1);
output(0, 2) <= input(2);
output(0, 3) <= input(3);
output(0, 4) <= input(4);
output(0, 5) <= input(5);
output(0, 6) <= input(6);
output(0, 7) <= input(7);
output(0, 8) <= input(8);
output(0, 9) <= input(9);
output(0, 10) <= input(10);
output(0, 11) <= input(11);
output(0, 12) <= input(12);
output(0, 13) <= input(13);
output(0, 14) <= input(14);
output(0, 15) <= input(15);
output(0, 16) <= input(0);
output(0, 17) <= input(1);
output(0, 18) <= input(2);
output(0, 19) <= input(3);
output(0, 20) <= input(4);
output(0, 21) <= input(5);
output(0, 22) <= input(6);
output(0, 23) <= input(7);
output(0, 24) <= input(8);
output(0, 25) <= input(9);
output(0, 26) <= input(10);
output(0, 27) <= input(11);
output(0, 28) <= input(12);
output(0, 29) <= input(13);
output(0, 30) <= input(14);
output(0, 31) <= input(15);
output(0, 32) <= input(16);
output(0, 33) <= input(17);
output(0, 34) <= input(18);
output(0, 35) <= input(19);
output(0, 36) <= input(20);
output(0, 37) <= input(21);
output(0, 38) <= input(22);
output(0, 39) <= input(23);
output(0, 40) <= input(24);
output(0, 41) <= input(25);
output(0, 42) <= input(26);
output(0, 43) <= input(27);
output(0, 44) <= input(28);
output(0, 45) <= input(29);
output(0, 46) <= input(30);
output(0, 47) <= input(31);
output(0, 48) <= input(16);
output(0, 49) <= input(17);
output(0, 50) <= input(18);
output(0, 51) <= input(19);
output(0, 52) <= input(20);
output(0, 53) <= input(21);
output(0, 54) <= input(22);
output(0, 55) <= input(23);
output(0, 56) <= input(24);
output(0, 57) <= input(25);
output(0, 58) <= input(26);
output(0, 59) <= input(27);
output(0, 60) <= input(28);
output(0, 61) <= input(29);
output(0, 62) <= input(30);
output(0, 63) <= input(31);
output(0, 64) <= input(16);
output(0, 65) <= input(17);
output(0, 66) <= input(18);
output(0, 67) <= input(19);
output(0, 68) <= input(20);
output(0, 69) <= input(21);
output(0, 70) <= input(22);
output(0, 71) <= input(23);
output(0, 72) <= input(24);
output(0, 73) <= input(25);
output(0, 74) <= input(26);
output(0, 75) <= input(27);
output(0, 76) <= input(28);
output(0, 77) <= input(29);
output(0, 78) <= input(30);
output(0, 79) <= input(31);
output(0, 80) <= input(1);
output(0, 81) <= input(2);
output(0, 82) <= input(3);
output(0, 83) <= input(4);
output(0, 84) <= input(5);
output(0, 85) <= input(6);
output(0, 86) <= input(7);
output(0, 87) <= input(8);
output(0, 88) <= input(9);
output(0, 89) <= input(10);
output(0, 90) <= input(11);
output(0, 91) <= input(12);
output(0, 92) <= input(13);
output(0, 93) <= input(14);
output(0, 94) <= input(15);
output(0, 95) <= input(32);
output(0, 96) <= input(1);
output(0, 97) <= input(2);
output(0, 98) <= input(3);
output(0, 99) <= input(4);
output(0, 100) <= input(5);
output(0, 101) <= input(6);
output(0, 102) <= input(7);
output(0, 103) <= input(8);
output(0, 104) <= input(9);
output(0, 105) <= input(10);
output(0, 106) <= input(11);
output(0, 107) <= input(12);
output(0, 108) <= input(13);
output(0, 109) <= input(14);
output(0, 110) <= input(15);
output(0, 111) <= input(32);
output(0, 112) <= input(17);
output(0, 113) <= input(18);
output(0, 114) <= input(19);
output(0, 115) <= input(20);
output(0, 116) <= input(21);
output(0, 117) <= input(22);
output(0, 118) <= input(23);
output(0, 119) <= input(24);
output(0, 120) <= input(25);
output(0, 121) <= input(26);
output(0, 122) <= input(27);
output(0, 123) <= input(28);
output(0, 124) <= input(29);
output(0, 125) <= input(30);
output(0, 126) <= input(31);
output(0, 127) <= input(33);
output(0, 128) <= input(17);
output(0, 129) <= input(18);
output(0, 130) <= input(19);
output(0, 131) <= input(20);
output(0, 132) <= input(21);
output(0, 133) <= input(22);
output(0, 134) <= input(23);
output(0, 135) <= input(24);
output(0, 136) <= input(25);
output(0, 137) <= input(26);
output(0, 138) <= input(27);
output(0, 139) <= input(28);
output(0, 140) <= input(29);
output(0, 141) <= input(30);
output(0, 142) <= input(31);
output(0, 143) <= input(33);
output(0, 144) <= input(17);
output(0, 145) <= input(18);
output(0, 146) <= input(19);
output(0, 147) <= input(20);
output(0, 148) <= input(21);
output(0, 149) <= input(22);
output(0, 150) <= input(23);
output(0, 151) <= input(24);
output(0, 152) <= input(25);
output(0, 153) <= input(26);
output(0, 154) <= input(27);
output(0, 155) <= input(28);
output(0, 156) <= input(29);
output(0, 157) <= input(30);
output(0, 158) <= input(31);
output(0, 159) <= input(33);
output(0, 160) <= input(2);
output(0, 161) <= input(3);
output(0, 162) <= input(4);
output(0, 163) <= input(5);
output(0, 164) <= input(6);
output(0, 165) <= input(7);
output(0, 166) <= input(8);
output(0, 167) <= input(9);
output(0, 168) <= input(10);
output(0, 169) <= input(11);
output(0, 170) <= input(12);
output(0, 171) <= input(13);
output(0, 172) <= input(14);
output(0, 173) <= input(15);
output(0, 174) <= input(32);
output(0, 175) <= input(34);
output(0, 176) <= input(2);
output(0, 177) <= input(3);
output(0, 178) <= input(4);
output(0, 179) <= input(5);
output(0, 180) <= input(6);
output(0, 181) <= input(7);
output(0, 182) <= input(8);
output(0, 183) <= input(9);
output(0, 184) <= input(10);
output(0, 185) <= input(11);
output(0, 186) <= input(12);
output(0, 187) <= input(13);
output(0, 188) <= input(14);
output(0, 189) <= input(15);
output(0, 190) <= input(32);
output(0, 191) <= input(34);
output(0, 192) <= input(2);
output(0, 193) <= input(3);
output(0, 194) <= input(4);
output(0, 195) <= input(5);
output(0, 196) <= input(6);
output(0, 197) <= input(7);
output(0, 198) <= input(8);
output(0, 199) <= input(9);
output(0, 200) <= input(10);
output(0, 201) <= input(11);
output(0, 202) <= input(12);
output(0, 203) <= input(13);
output(0, 204) <= input(14);
output(0, 205) <= input(15);
output(0, 206) <= input(32);
output(0, 207) <= input(34);
output(0, 208) <= input(18);
output(0, 209) <= input(19);
output(0, 210) <= input(20);
output(0, 211) <= input(21);
output(0, 212) <= input(22);
output(0, 213) <= input(23);
output(0, 214) <= input(24);
output(0, 215) <= input(25);
output(0, 216) <= input(26);
output(0, 217) <= input(27);
output(0, 218) <= input(28);
output(0, 219) <= input(29);
output(0, 220) <= input(30);
output(0, 221) <= input(31);
output(0, 222) <= input(33);
output(0, 223) <= input(35);
output(0, 224) <= input(18);
output(0, 225) <= input(19);
output(0, 226) <= input(20);
output(0, 227) <= input(21);
output(0, 228) <= input(22);
output(0, 229) <= input(23);
output(0, 230) <= input(24);
output(0, 231) <= input(25);
output(0, 232) <= input(26);
output(0, 233) <= input(27);
output(0, 234) <= input(28);
output(0, 235) <= input(29);
output(0, 236) <= input(30);
output(0, 237) <= input(31);
output(0, 238) <= input(33);
output(0, 239) <= input(35);
output(0, 240) <= input(3);
output(0, 241) <= input(4);
output(0, 242) <= input(5);
output(0, 243) <= input(6);
output(0, 244) <= input(7);
output(0, 245) <= input(8);
output(0, 246) <= input(9);
output(0, 247) <= input(10);
output(0, 248) <= input(11);
output(0, 249) <= input(12);
output(0, 250) <= input(13);
output(0, 251) <= input(14);
output(0, 252) <= input(15);
output(0, 253) <= input(32);
output(0, 254) <= input(34);
output(0, 255) <= input(36);
output(1, 0) <= input(0);
output(1, 1) <= input(1);
output(1, 2) <= input(2);
output(1, 3) <= input(3);
output(1, 4) <= input(4);
output(1, 5) <= input(5);
output(1, 6) <= input(6);
output(1, 7) <= input(7);
output(1, 8) <= input(8);
output(1, 9) <= input(9);
output(1, 10) <= input(10);
output(1, 11) <= input(11);
output(1, 12) <= input(12);
output(1, 13) <= input(13);
output(1, 14) <= input(14);
output(1, 15) <= input(15);
output(1, 16) <= input(16);
output(1, 17) <= input(17);
output(1, 18) <= input(18);
output(1, 19) <= input(19);
output(1, 20) <= input(20);
output(1, 21) <= input(21);
output(1, 22) <= input(22);
output(1, 23) <= input(23);
output(1, 24) <= input(24);
output(1, 25) <= input(25);
output(1, 26) <= input(26);
output(1, 27) <= input(27);
output(1, 28) <= input(28);
output(1, 29) <= input(29);
output(1, 30) <= input(30);
output(1, 31) <= input(31);
output(1, 32) <= input(16);
output(1, 33) <= input(17);
output(1, 34) <= input(18);
output(1, 35) <= input(19);
output(1, 36) <= input(20);
output(1, 37) <= input(21);
output(1, 38) <= input(22);
output(1, 39) <= input(23);
output(1, 40) <= input(24);
output(1, 41) <= input(25);
output(1, 42) <= input(26);
output(1, 43) <= input(27);
output(1, 44) <= input(28);
output(1, 45) <= input(29);
output(1, 46) <= input(30);
output(1, 47) <= input(31);
output(1, 48) <= input(1);
output(1, 49) <= input(2);
output(1, 50) <= input(3);
output(1, 51) <= input(4);
output(1, 52) <= input(5);
output(1, 53) <= input(6);
output(1, 54) <= input(7);
output(1, 55) <= input(8);
output(1, 56) <= input(9);
output(1, 57) <= input(10);
output(1, 58) <= input(11);
output(1, 59) <= input(12);
output(1, 60) <= input(13);
output(1, 61) <= input(14);
output(1, 62) <= input(15);
output(1, 63) <= input(32);
output(1, 64) <= input(1);
output(1, 65) <= input(2);
output(1, 66) <= input(3);
output(1, 67) <= input(4);
output(1, 68) <= input(5);
output(1, 69) <= input(6);
output(1, 70) <= input(7);
output(1, 71) <= input(8);
output(1, 72) <= input(9);
output(1, 73) <= input(10);
output(1, 74) <= input(11);
output(1, 75) <= input(12);
output(1, 76) <= input(13);
output(1, 77) <= input(14);
output(1, 78) <= input(15);
output(1, 79) <= input(32);
output(1, 80) <= input(17);
output(1, 81) <= input(18);
output(1, 82) <= input(19);
output(1, 83) <= input(20);
output(1, 84) <= input(21);
output(1, 85) <= input(22);
output(1, 86) <= input(23);
output(1, 87) <= input(24);
output(1, 88) <= input(25);
output(1, 89) <= input(26);
output(1, 90) <= input(27);
output(1, 91) <= input(28);
output(1, 92) <= input(29);
output(1, 93) <= input(30);
output(1, 94) <= input(31);
output(1, 95) <= input(33);
output(1, 96) <= input(17);
output(1, 97) <= input(18);
output(1, 98) <= input(19);
output(1, 99) <= input(20);
output(1, 100) <= input(21);
output(1, 101) <= input(22);
output(1, 102) <= input(23);
output(1, 103) <= input(24);
output(1, 104) <= input(25);
output(1, 105) <= input(26);
output(1, 106) <= input(27);
output(1, 107) <= input(28);
output(1, 108) <= input(29);
output(1, 109) <= input(30);
output(1, 110) <= input(31);
output(1, 111) <= input(33);
output(1, 112) <= input(2);
output(1, 113) <= input(3);
output(1, 114) <= input(4);
output(1, 115) <= input(5);
output(1, 116) <= input(6);
output(1, 117) <= input(7);
output(1, 118) <= input(8);
output(1, 119) <= input(9);
output(1, 120) <= input(10);
output(1, 121) <= input(11);
output(1, 122) <= input(12);
output(1, 123) <= input(13);
output(1, 124) <= input(14);
output(1, 125) <= input(15);
output(1, 126) <= input(32);
output(1, 127) <= input(34);
output(1, 128) <= input(2);
output(1, 129) <= input(3);
output(1, 130) <= input(4);
output(1, 131) <= input(5);
output(1, 132) <= input(6);
output(1, 133) <= input(7);
output(1, 134) <= input(8);
output(1, 135) <= input(9);
output(1, 136) <= input(10);
output(1, 137) <= input(11);
output(1, 138) <= input(12);
output(1, 139) <= input(13);
output(1, 140) <= input(14);
output(1, 141) <= input(15);
output(1, 142) <= input(32);
output(1, 143) <= input(34);
output(1, 144) <= input(18);
output(1, 145) <= input(19);
output(1, 146) <= input(20);
output(1, 147) <= input(21);
output(1, 148) <= input(22);
output(1, 149) <= input(23);
output(1, 150) <= input(24);
output(1, 151) <= input(25);
output(1, 152) <= input(26);
output(1, 153) <= input(27);
output(1, 154) <= input(28);
output(1, 155) <= input(29);
output(1, 156) <= input(30);
output(1, 157) <= input(31);
output(1, 158) <= input(33);
output(1, 159) <= input(35);
output(1, 160) <= input(18);
output(1, 161) <= input(19);
output(1, 162) <= input(20);
output(1, 163) <= input(21);
output(1, 164) <= input(22);
output(1, 165) <= input(23);
output(1, 166) <= input(24);
output(1, 167) <= input(25);
output(1, 168) <= input(26);
output(1, 169) <= input(27);
output(1, 170) <= input(28);
output(1, 171) <= input(29);
output(1, 172) <= input(30);
output(1, 173) <= input(31);
output(1, 174) <= input(33);
output(1, 175) <= input(35);
output(1, 176) <= input(3);
output(1, 177) <= input(4);
output(1, 178) <= input(5);
output(1, 179) <= input(6);
output(1, 180) <= input(7);
output(1, 181) <= input(8);
output(1, 182) <= input(9);
output(1, 183) <= input(10);
output(1, 184) <= input(11);
output(1, 185) <= input(12);
output(1, 186) <= input(13);
output(1, 187) <= input(14);
output(1, 188) <= input(15);
output(1, 189) <= input(32);
output(1, 190) <= input(34);
output(1, 191) <= input(36);
output(1, 192) <= input(3);
output(1, 193) <= input(4);
output(1, 194) <= input(5);
output(1, 195) <= input(6);
output(1, 196) <= input(7);
output(1, 197) <= input(8);
output(1, 198) <= input(9);
output(1, 199) <= input(10);
output(1, 200) <= input(11);
output(1, 201) <= input(12);
output(1, 202) <= input(13);
output(1, 203) <= input(14);
output(1, 204) <= input(15);
output(1, 205) <= input(32);
output(1, 206) <= input(34);
output(1, 207) <= input(36);
output(1, 208) <= input(19);
output(1, 209) <= input(20);
output(1, 210) <= input(21);
output(1, 211) <= input(22);
output(1, 212) <= input(23);
output(1, 213) <= input(24);
output(1, 214) <= input(25);
output(1, 215) <= input(26);
output(1, 216) <= input(27);
output(1, 217) <= input(28);
output(1, 218) <= input(29);
output(1, 219) <= input(30);
output(1, 220) <= input(31);
output(1, 221) <= input(33);
output(1, 222) <= input(35);
output(1, 223) <= input(37);
output(1, 224) <= input(19);
output(1, 225) <= input(20);
output(1, 226) <= input(21);
output(1, 227) <= input(22);
output(1, 228) <= input(23);
output(1, 229) <= input(24);
output(1, 230) <= input(25);
output(1, 231) <= input(26);
output(1, 232) <= input(27);
output(1, 233) <= input(28);
output(1, 234) <= input(29);
output(1, 235) <= input(30);
output(1, 236) <= input(31);
output(1, 237) <= input(33);
output(1, 238) <= input(35);
output(1, 239) <= input(37);
output(1, 240) <= input(4);
output(1, 241) <= input(5);
output(1, 242) <= input(6);
output(1, 243) <= input(7);
output(1, 244) <= input(8);
output(1, 245) <= input(9);
output(1, 246) <= input(10);
output(1, 247) <= input(11);
output(1, 248) <= input(12);
output(1, 249) <= input(13);
output(1, 250) <= input(14);
output(1, 251) <= input(15);
output(1, 252) <= input(32);
output(1, 253) <= input(34);
output(1, 254) <= input(36);
output(1, 255) <= input(38);
output(2, 0) <= input(0);
output(2, 1) <= input(1);
output(2, 2) <= input(2);
output(2, 3) <= input(3);
output(2, 4) <= input(4);
output(2, 5) <= input(5);
output(2, 6) <= input(6);
output(2, 7) <= input(7);
output(2, 8) <= input(8);
output(2, 9) <= input(9);
output(2, 10) <= input(10);
output(2, 11) <= input(11);
output(2, 12) <= input(12);
output(2, 13) <= input(13);
output(2, 14) <= input(14);
output(2, 15) <= input(15);
output(2, 16) <= input(16);
output(2, 17) <= input(17);
output(2, 18) <= input(18);
output(2, 19) <= input(19);
output(2, 20) <= input(20);
output(2, 21) <= input(21);
output(2, 22) <= input(22);
output(2, 23) <= input(23);
output(2, 24) <= input(24);
output(2, 25) <= input(25);
output(2, 26) <= input(26);
output(2, 27) <= input(27);
output(2, 28) <= input(28);
output(2, 29) <= input(29);
output(2, 30) <= input(30);
output(2, 31) <= input(31);
output(2, 32) <= input(16);
output(2, 33) <= input(17);
output(2, 34) <= input(18);
output(2, 35) <= input(19);
output(2, 36) <= input(20);
output(2, 37) <= input(21);
output(2, 38) <= input(22);
output(2, 39) <= input(23);
output(2, 40) <= input(24);
output(2, 41) <= input(25);
output(2, 42) <= input(26);
output(2, 43) <= input(27);
output(2, 44) <= input(28);
output(2, 45) <= input(29);
output(2, 46) <= input(30);
output(2, 47) <= input(31);
output(2, 48) <= input(1);
output(2, 49) <= input(2);
output(2, 50) <= input(3);
output(2, 51) <= input(4);
output(2, 52) <= input(5);
output(2, 53) <= input(6);
output(2, 54) <= input(7);
output(2, 55) <= input(8);
output(2, 56) <= input(9);
output(2, 57) <= input(10);
output(2, 58) <= input(11);
output(2, 59) <= input(12);
output(2, 60) <= input(13);
output(2, 61) <= input(14);
output(2, 62) <= input(15);
output(2, 63) <= input(32);
output(2, 64) <= input(17);
output(2, 65) <= input(18);
output(2, 66) <= input(19);
output(2, 67) <= input(20);
output(2, 68) <= input(21);
output(2, 69) <= input(22);
output(2, 70) <= input(23);
output(2, 71) <= input(24);
output(2, 72) <= input(25);
output(2, 73) <= input(26);
output(2, 74) <= input(27);
output(2, 75) <= input(28);
output(2, 76) <= input(29);
output(2, 77) <= input(30);
output(2, 78) <= input(31);
output(2, 79) <= input(33);
output(2, 80) <= input(17);
output(2, 81) <= input(18);
output(2, 82) <= input(19);
output(2, 83) <= input(20);
output(2, 84) <= input(21);
output(2, 85) <= input(22);
output(2, 86) <= input(23);
output(2, 87) <= input(24);
output(2, 88) <= input(25);
output(2, 89) <= input(26);
output(2, 90) <= input(27);
output(2, 91) <= input(28);
output(2, 92) <= input(29);
output(2, 93) <= input(30);
output(2, 94) <= input(31);
output(2, 95) <= input(33);
output(2, 96) <= input(2);
output(2, 97) <= input(3);
output(2, 98) <= input(4);
output(2, 99) <= input(5);
output(2, 100) <= input(6);
output(2, 101) <= input(7);
output(2, 102) <= input(8);
output(2, 103) <= input(9);
output(2, 104) <= input(10);
output(2, 105) <= input(11);
output(2, 106) <= input(12);
output(2, 107) <= input(13);
output(2, 108) <= input(14);
output(2, 109) <= input(15);
output(2, 110) <= input(32);
output(2, 111) <= input(34);
output(2, 112) <= input(18);
output(2, 113) <= input(19);
output(2, 114) <= input(20);
output(2, 115) <= input(21);
output(2, 116) <= input(22);
output(2, 117) <= input(23);
output(2, 118) <= input(24);
output(2, 119) <= input(25);
output(2, 120) <= input(26);
output(2, 121) <= input(27);
output(2, 122) <= input(28);
output(2, 123) <= input(29);
output(2, 124) <= input(30);
output(2, 125) <= input(31);
output(2, 126) <= input(33);
output(2, 127) <= input(35);
output(2, 128) <= input(18);
output(2, 129) <= input(19);
output(2, 130) <= input(20);
output(2, 131) <= input(21);
output(2, 132) <= input(22);
output(2, 133) <= input(23);
output(2, 134) <= input(24);
output(2, 135) <= input(25);
output(2, 136) <= input(26);
output(2, 137) <= input(27);
output(2, 138) <= input(28);
output(2, 139) <= input(29);
output(2, 140) <= input(30);
output(2, 141) <= input(31);
output(2, 142) <= input(33);
output(2, 143) <= input(35);
output(2, 144) <= input(3);
output(2, 145) <= input(4);
output(2, 146) <= input(5);
output(2, 147) <= input(6);
output(2, 148) <= input(7);
output(2, 149) <= input(8);
output(2, 150) <= input(9);
output(2, 151) <= input(10);
output(2, 152) <= input(11);
output(2, 153) <= input(12);
output(2, 154) <= input(13);
output(2, 155) <= input(14);
output(2, 156) <= input(15);
output(2, 157) <= input(32);
output(2, 158) <= input(34);
output(2, 159) <= input(36);
output(2, 160) <= input(3);
output(2, 161) <= input(4);
output(2, 162) <= input(5);
output(2, 163) <= input(6);
output(2, 164) <= input(7);
output(2, 165) <= input(8);
output(2, 166) <= input(9);
output(2, 167) <= input(10);
output(2, 168) <= input(11);
output(2, 169) <= input(12);
output(2, 170) <= input(13);
output(2, 171) <= input(14);
output(2, 172) <= input(15);
output(2, 173) <= input(32);
output(2, 174) <= input(34);
output(2, 175) <= input(36);
output(2, 176) <= input(19);
output(2, 177) <= input(20);
output(2, 178) <= input(21);
output(2, 179) <= input(22);
output(2, 180) <= input(23);
output(2, 181) <= input(24);
output(2, 182) <= input(25);
output(2, 183) <= input(26);
output(2, 184) <= input(27);
output(2, 185) <= input(28);
output(2, 186) <= input(29);
output(2, 187) <= input(30);
output(2, 188) <= input(31);
output(2, 189) <= input(33);
output(2, 190) <= input(35);
output(2, 191) <= input(37);
output(2, 192) <= input(4);
output(2, 193) <= input(5);
output(2, 194) <= input(6);
output(2, 195) <= input(7);
output(2, 196) <= input(8);
output(2, 197) <= input(9);
output(2, 198) <= input(10);
output(2, 199) <= input(11);
output(2, 200) <= input(12);
output(2, 201) <= input(13);
output(2, 202) <= input(14);
output(2, 203) <= input(15);
output(2, 204) <= input(32);
output(2, 205) <= input(34);
output(2, 206) <= input(36);
output(2, 207) <= input(38);
output(2, 208) <= input(4);
output(2, 209) <= input(5);
output(2, 210) <= input(6);
output(2, 211) <= input(7);
output(2, 212) <= input(8);
output(2, 213) <= input(9);
output(2, 214) <= input(10);
output(2, 215) <= input(11);
output(2, 216) <= input(12);
output(2, 217) <= input(13);
output(2, 218) <= input(14);
output(2, 219) <= input(15);
output(2, 220) <= input(32);
output(2, 221) <= input(34);
output(2, 222) <= input(36);
output(2, 223) <= input(38);
output(2, 224) <= input(20);
output(2, 225) <= input(21);
output(2, 226) <= input(22);
output(2, 227) <= input(23);
output(2, 228) <= input(24);
output(2, 229) <= input(25);
output(2, 230) <= input(26);
output(2, 231) <= input(27);
output(2, 232) <= input(28);
output(2, 233) <= input(29);
output(2, 234) <= input(30);
output(2, 235) <= input(31);
output(2, 236) <= input(33);
output(2, 237) <= input(35);
output(2, 238) <= input(37);
output(2, 239) <= input(39);
output(2, 240) <= input(5);
output(2, 241) <= input(6);
output(2, 242) <= input(7);
output(2, 243) <= input(8);
output(2, 244) <= input(9);
output(2, 245) <= input(10);
output(2, 246) <= input(11);
output(2, 247) <= input(12);
output(2, 248) <= input(13);
output(2, 249) <= input(14);
output(2, 250) <= input(15);
output(2, 251) <= input(32);
output(2, 252) <= input(34);
output(2, 253) <= input(36);
output(2, 254) <= input(38);
output(2, 255) <= input(40);
output(3, 0) <= input(0);
output(3, 1) <= input(1);
output(3, 2) <= input(2);
output(3, 3) <= input(3);
output(3, 4) <= input(4);
output(3, 5) <= input(5);
output(3, 6) <= input(6);
output(3, 7) <= input(7);
output(3, 8) <= input(8);
output(3, 9) <= input(9);
output(3, 10) <= input(10);
output(3, 11) <= input(11);
output(3, 12) <= input(12);
output(3, 13) <= input(13);
output(3, 14) <= input(14);
output(3, 15) <= input(15);
output(3, 16) <= input(16);
output(3, 17) <= input(17);
output(3, 18) <= input(18);
output(3, 19) <= input(19);
output(3, 20) <= input(20);
output(3, 21) <= input(21);
output(3, 22) <= input(22);
output(3, 23) <= input(23);
output(3, 24) <= input(24);
output(3, 25) <= input(25);
output(3, 26) <= input(26);
output(3, 27) <= input(27);
output(3, 28) <= input(28);
output(3, 29) <= input(29);
output(3, 30) <= input(30);
output(3, 31) <= input(31);
output(3, 32) <= input(1);
output(3, 33) <= input(2);
output(3, 34) <= input(3);
output(3, 35) <= input(4);
output(3, 36) <= input(5);
output(3, 37) <= input(6);
output(3, 38) <= input(7);
output(3, 39) <= input(8);
output(3, 40) <= input(9);
output(3, 41) <= input(10);
output(3, 42) <= input(11);
output(3, 43) <= input(12);
output(3, 44) <= input(13);
output(3, 45) <= input(14);
output(3, 46) <= input(15);
output(3, 47) <= input(32);
output(3, 48) <= input(17);
output(3, 49) <= input(18);
output(3, 50) <= input(19);
output(3, 51) <= input(20);
output(3, 52) <= input(21);
output(3, 53) <= input(22);
output(3, 54) <= input(23);
output(3, 55) <= input(24);
output(3, 56) <= input(25);
output(3, 57) <= input(26);
output(3, 58) <= input(27);
output(3, 59) <= input(28);
output(3, 60) <= input(29);
output(3, 61) <= input(30);
output(3, 62) <= input(31);
output(3, 63) <= input(33);
output(3, 64) <= input(17);
output(3, 65) <= input(18);
output(3, 66) <= input(19);
output(3, 67) <= input(20);
output(3, 68) <= input(21);
output(3, 69) <= input(22);
output(3, 70) <= input(23);
output(3, 71) <= input(24);
output(3, 72) <= input(25);
output(3, 73) <= input(26);
output(3, 74) <= input(27);
output(3, 75) <= input(28);
output(3, 76) <= input(29);
output(3, 77) <= input(30);
output(3, 78) <= input(31);
output(3, 79) <= input(33);
output(3, 80) <= input(2);
output(3, 81) <= input(3);
output(3, 82) <= input(4);
output(3, 83) <= input(5);
output(3, 84) <= input(6);
output(3, 85) <= input(7);
output(3, 86) <= input(8);
output(3, 87) <= input(9);
output(3, 88) <= input(10);
output(3, 89) <= input(11);
output(3, 90) <= input(12);
output(3, 91) <= input(13);
output(3, 92) <= input(14);
output(3, 93) <= input(15);
output(3, 94) <= input(32);
output(3, 95) <= input(34);
output(3, 96) <= input(18);
output(3, 97) <= input(19);
output(3, 98) <= input(20);
output(3, 99) <= input(21);
output(3, 100) <= input(22);
output(3, 101) <= input(23);
output(3, 102) <= input(24);
output(3, 103) <= input(25);
output(3, 104) <= input(26);
output(3, 105) <= input(27);
output(3, 106) <= input(28);
output(3, 107) <= input(29);
output(3, 108) <= input(30);
output(3, 109) <= input(31);
output(3, 110) <= input(33);
output(3, 111) <= input(35);
output(3, 112) <= input(3);
output(3, 113) <= input(4);
output(3, 114) <= input(5);
output(3, 115) <= input(6);
output(3, 116) <= input(7);
output(3, 117) <= input(8);
output(3, 118) <= input(9);
output(3, 119) <= input(10);
output(3, 120) <= input(11);
output(3, 121) <= input(12);
output(3, 122) <= input(13);
output(3, 123) <= input(14);
output(3, 124) <= input(15);
output(3, 125) <= input(32);
output(3, 126) <= input(34);
output(3, 127) <= input(36);
output(3, 128) <= input(3);
output(3, 129) <= input(4);
output(3, 130) <= input(5);
output(3, 131) <= input(6);
output(3, 132) <= input(7);
output(3, 133) <= input(8);
output(3, 134) <= input(9);
output(3, 135) <= input(10);
output(3, 136) <= input(11);
output(3, 137) <= input(12);
output(3, 138) <= input(13);
output(3, 139) <= input(14);
output(3, 140) <= input(15);
output(3, 141) <= input(32);
output(3, 142) <= input(34);
output(3, 143) <= input(36);
output(3, 144) <= input(19);
output(3, 145) <= input(20);
output(3, 146) <= input(21);
output(3, 147) <= input(22);
output(3, 148) <= input(23);
output(3, 149) <= input(24);
output(3, 150) <= input(25);
output(3, 151) <= input(26);
output(3, 152) <= input(27);
output(3, 153) <= input(28);
output(3, 154) <= input(29);
output(3, 155) <= input(30);
output(3, 156) <= input(31);
output(3, 157) <= input(33);
output(3, 158) <= input(35);
output(3, 159) <= input(37);
output(3, 160) <= input(4);
output(3, 161) <= input(5);
output(3, 162) <= input(6);
output(3, 163) <= input(7);
output(3, 164) <= input(8);
output(3, 165) <= input(9);
output(3, 166) <= input(10);
output(3, 167) <= input(11);
output(3, 168) <= input(12);
output(3, 169) <= input(13);
output(3, 170) <= input(14);
output(3, 171) <= input(15);
output(3, 172) <= input(32);
output(3, 173) <= input(34);
output(3, 174) <= input(36);
output(3, 175) <= input(38);
output(3, 176) <= input(20);
output(3, 177) <= input(21);
output(3, 178) <= input(22);
output(3, 179) <= input(23);
output(3, 180) <= input(24);
output(3, 181) <= input(25);
output(3, 182) <= input(26);
output(3, 183) <= input(27);
output(3, 184) <= input(28);
output(3, 185) <= input(29);
output(3, 186) <= input(30);
output(3, 187) <= input(31);
output(3, 188) <= input(33);
output(3, 189) <= input(35);
output(3, 190) <= input(37);
output(3, 191) <= input(39);
output(3, 192) <= input(20);
output(3, 193) <= input(21);
output(3, 194) <= input(22);
output(3, 195) <= input(23);
output(3, 196) <= input(24);
output(3, 197) <= input(25);
output(3, 198) <= input(26);
output(3, 199) <= input(27);
output(3, 200) <= input(28);
output(3, 201) <= input(29);
output(3, 202) <= input(30);
output(3, 203) <= input(31);
output(3, 204) <= input(33);
output(3, 205) <= input(35);
output(3, 206) <= input(37);
output(3, 207) <= input(39);
output(3, 208) <= input(5);
output(3, 209) <= input(6);
output(3, 210) <= input(7);
output(3, 211) <= input(8);
output(3, 212) <= input(9);
output(3, 213) <= input(10);
output(3, 214) <= input(11);
output(3, 215) <= input(12);
output(3, 216) <= input(13);
output(3, 217) <= input(14);
output(3, 218) <= input(15);
output(3, 219) <= input(32);
output(3, 220) <= input(34);
output(3, 221) <= input(36);
output(3, 222) <= input(38);
output(3, 223) <= input(40);
output(3, 224) <= input(21);
output(3, 225) <= input(22);
output(3, 226) <= input(23);
output(3, 227) <= input(24);
output(3, 228) <= input(25);
output(3, 229) <= input(26);
output(3, 230) <= input(27);
output(3, 231) <= input(28);
output(3, 232) <= input(29);
output(3, 233) <= input(30);
output(3, 234) <= input(31);
output(3, 235) <= input(33);
output(3, 236) <= input(35);
output(3, 237) <= input(37);
output(3, 238) <= input(39);
output(3, 239) <= input(41);
output(3, 240) <= input(6);
output(3, 241) <= input(7);
output(3, 242) <= input(8);
output(3, 243) <= input(9);
output(3, 244) <= input(10);
output(3, 245) <= input(11);
output(3, 246) <= input(12);
output(3, 247) <= input(13);
output(3, 248) <= input(14);
output(3, 249) <= input(15);
output(3, 250) <= input(32);
output(3, 251) <= input(34);
output(3, 252) <= input(36);
output(3, 253) <= input(38);
output(3, 254) <= input(40);
output(3, 255) <= input(42);
output(4, 0) <= input(0);
output(4, 1) <= input(1);
output(4, 2) <= input(2);
output(4, 3) <= input(3);
output(4, 4) <= input(4);
output(4, 5) <= input(5);
output(4, 6) <= input(6);
output(4, 7) <= input(7);
output(4, 8) <= input(8);
output(4, 9) <= input(9);
output(4, 10) <= input(10);
output(4, 11) <= input(11);
output(4, 12) <= input(12);
output(4, 13) <= input(13);
output(4, 14) <= input(14);
output(4, 15) <= input(15);
output(4, 16) <= input(16);
output(4, 17) <= input(17);
output(4, 18) <= input(18);
output(4, 19) <= input(19);
output(4, 20) <= input(20);
output(4, 21) <= input(21);
output(4, 22) <= input(22);
output(4, 23) <= input(23);
output(4, 24) <= input(24);
output(4, 25) <= input(25);
output(4, 26) <= input(26);
output(4, 27) <= input(27);
output(4, 28) <= input(28);
output(4, 29) <= input(29);
output(4, 30) <= input(30);
output(4, 31) <= input(31);
output(4, 32) <= input(1);
output(4, 33) <= input(2);
output(4, 34) <= input(3);
output(4, 35) <= input(4);
output(4, 36) <= input(5);
output(4, 37) <= input(6);
output(4, 38) <= input(7);
output(4, 39) <= input(8);
output(4, 40) <= input(9);
output(4, 41) <= input(10);
output(4, 42) <= input(11);
output(4, 43) <= input(12);
output(4, 44) <= input(13);
output(4, 45) <= input(14);
output(4, 46) <= input(15);
output(4, 47) <= input(32);
output(4, 48) <= input(17);
output(4, 49) <= input(18);
output(4, 50) <= input(19);
output(4, 51) <= input(20);
output(4, 52) <= input(21);
output(4, 53) <= input(22);
output(4, 54) <= input(23);
output(4, 55) <= input(24);
output(4, 56) <= input(25);
output(4, 57) <= input(26);
output(4, 58) <= input(27);
output(4, 59) <= input(28);
output(4, 60) <= input(29);
output(4, 61) <= input(30);
output(4, 62) <= input(31);
output(4, 63) <= input(33);
output(4, 64) <= input(2);
output(4, 65) <= input(3);
output(4, 66) <= input(4);
output(4, 67) <= input(5);
output(4, 68) <= input(6);
output(4, 69) <= input(7);
output(4, 70) <= input(8);
output(4, 71) <= input(9);
output(4, 72) <= input(10);
output(4, 73) <= input(11);
output(4, 74) <= input(12);
output(4, 75) <= input(13);
output(4, 76) <= input(14);
output(4, 77) <= input(15);
output(4, 78) <= input(32);
output(4, 79) <= input(34);
output(4, 80) <= input(18);
output(4, 81) <= input(19);
output(4, 82) <= input(20);
output(4, 83) <= input(21);
output(4, 84) <= input(22);
output(4, 85) <= input(23);
output(4, 86) <= input(24);
output(4, 87) <= input(25);
output(4, 88) <= input(26);
output(4, 89) <= input(27);
output(4, 90) <= input(28);
output(4, 91) <= input(29);
output(4, 92) <= input(30);
output(4, 93) <= input(31);
output(4, 94) <= input(33);
output(4, 95) <= input(35);
output(4, 96) <= input(3);
output(4, 97) <= input(4);
output(4, 98) <= input(5);
output(4, 99) <= input(6);
output(4, 100) <= input(7);
output(4, 101) <= input(8);
output(4, 102) <= input(9);
output(4, 103) <= input(10);
output(4, 104) <= input(11);
output(4, 105) <= input(12);
output(4, 106) <= input(13);
output(4, 107) <= input(14);
output(4, 108) <= input(15);
output(4, 109) <= input(32);
output(4, 110) <= input(34);
output(4, 111) <= input(36);
output(4, 112) <= input(19);
output(4, 113) <= input(20);
output(4, 114) <= input(21);
output(4, 115) <= input(22);
output(4, 116) <= input(23);
output(4, 117) <= input(24);
output(4, 118) <= input(25);
output(4, 119) <= input(26);
output(4, 120) <= input(27);
output(4, 121) <= input(28);
output(4, 122) <= input(29);
output(4, 123) <= input(30);
output(4, 124) <= input(31);
output(4, 125) <= input(33);
output(4, 126) <= input(35);
output(4, 127) <= input(37);
output(4, 128) <= input(19);
output(4, 129) <= input(20);
output(4, 130) <= input(21);
output(4, 131) <= input(22);
output(4, 132) <= input(23);
output(4, 133) <= input(24);
output(4, 134) <= input(25);
output(4, 135) <= input(26);
output(4, 136) <= input(27);
output(4, 137) <= input(28);
output(4, 138) <= input(29);
output(4, 139) <= input(30);
output(4, 140) <= input(31);
output(4, 141) <= input(33);
output(4, 142) <= input(35);
output(4, 143) <= input(37);
output(4, 144) <= input(4);
output(4, 145) <= input(5);
output(4, 146) <= input(6);
output(4, 147) <= input(7);
output(4, 148) <= input(8);
output(4, 149) <= input(9);
output(4, 150) <= input(10);
output(4, 151) <= input(11);
output(4, 152) <= input(12);
output(4, 153) <= input(13);
output(4, 154) <= input(14);
output(4, 155) <= input(15);
output(4, 156) <= input(32);
output(4, 157) <= input(34);
output(4, 158) <= input(36);
output(4, 159) <= input(38);
output(4, 160) <= input(20);
output(4, 161) <= input(21);
output(4, 162) <= input(22);
output(4, 163) <= input(23);
output(4, 164) <= input(24);
output(4, 165) <= input(25);
output(4, 166) <= input(26);
output(4, 167) <= input(27);
output(4, 168) <= input(28);
output(4, 169) <= input(29);
output(4, 170) <= input(30);
output(4, 171) <= input(31);
output(4, 172) <= input(33);
output(4, 173) <= input(35);
output(4, 174) <= input(37);
output(4, 175) <= input(39);
output(4, 176) <= input(5);
output(4, 177) <= input(6);
output(4, 178) <= input(7);
output(4, 179) <= input(8);
output(4, 180) <= input(9);
output(4, 181) <= input(10);
output(4, 182) <= input(11);
output(4, 183) <= input(12);
output(4, 184) <= input(13);
output(4, 185) <= input(14);
output(4, 186) <= input(15);
output(4, 187) <= input(32);
output(4, 188) <= input(34);
output(4, 189) <= input(36);
output(4, 190) <= input(38);
output(4, 191) <= input(40);
output(4, 192) <= input(21);
output(4, 193) <= input(22);
output(4, 194) <= input(23);
output(4, 195) <= input(24);
output(4, 196) <= input(25);
output(4, 197) <= input(26);
output(4, 198) <= input(27);
output(4, 199) <= input(28);
output(4, 200) <= input(29);
output(4, 201) <= input(30);
output(4, 202) <= input(31);
output(4, 203) <= input(33);
output(4, 204) <= input(35);
output(4, 205) <= input(37);
output(4, 206) <= input(39);
output(4, 207) <= input(41);
output(4, 208) <= input(6);
output(4, 209) <= input(7);
output(4, 210) <= input(8);
output(4, 211) <= input(9);
output(4, 212) <= input(10);
output(4, 213) <= input(11);
output(4, 214) <= input(12);
output(4, 215) <= input(13);
output(4, 216) <= input(14);
output(4, 217) <= input(15);
output(4, 218) <= input(32);
output(4, 219) <= input(34);
output(4, 220) <= input(36);
output(4, 221) <= input(38);
output(4, 222) <= input(40);
output(4, 223) <= input(42);
output(4, 224) <= input(22);
output(4, 225) <= input(23);
output(4, 226) <= input(24);
output(4, 227) <= input(25);
output(4, 228) <= input(26);
output(4, 229) <= input(27);
output(4, 230) <= input(28);
output(4, 231) <= input(29);
output(4, 232) <= input(30);
output(4, 233) <= input(31);
output(4, 234) <= input(33);
output(4, 235) <= input(35);
output(4, 236) <= input(37);
output(4, 237) <= input(39);
output(4, 238) <= input(41);
output(4, 239) <= input(43);
output(4, 240) <= input(7);
output(4, 241) <= input(8);
output(4, 242) <= input(9);
output(4, 243) <= input(10);
output(4, 244) <= input(11);
output(4, 245) <= input(12);
output(4, 246) <= input(13);
output(4, 247) <= input(14);
output(4, 248) <= input(15);
output(4, 249) <= input(32);
output(4, 250) <= input(34);
output(4, 251) <= input(36);
output(4, 252) <= input(38);
output(4, 253) <= input(40);
output(4, 254) <= input(42);
output(4, 255) <= input(44);
output(5, 0) <= input(16);
output(5, 1) <= input(17);
output(5, 2) <= input(18);
output(5, 3) <= input(19);
output(5, 4) <= input(20);
output(5, 5) <= input(21);
output(5, 6) <= input(22);
output(5, 7) <= input(23);
output(5, 8) <= input(24);
output(5, 9) <= input(25);
output(5, 10) <= input(26);
output(5, 11) <= input(27);
output(5, 12) <= input(28);
output(5, 13) <= input(29);
output(5, 14) <= input(30);
output(5, 15) <= input(31);
output(5, 16) <= input(1);
output(5, 17) <= input(2);
output(5, 18) <= input(3);
output(5, 19) <= input(4);
output(5, 20) <= input(5);
output(5, 21) <= input(6);
output(5, 22) <= input(7);
output(5, 23) <= input(8);
output(5, 24) <= input(9);
output(5, 25) <= input(10);
output(5, 26) <= input(11);
output(5, 27) <= input(12);
output(5, 28) <= input(13);
output(5, 29) <= input(14);
output(5, 30) <= input(15);
output(5, 31) <= input(32);
output(5, 32) <= input(17);
output(5, 33) <= input(18);
output(5, 34) <= input(19);
output(5, 35) <= input(20);
output(5, 36) <= input(21);
output(5, 37) <= input(22);
output(5, 38) <= input(23);
output(5, 39) <= input(24);
output(5, 40) <= input(25);
output(5, 41) <= input(26);
output(5, 42) <= input(27);
output(5, 43) <= input(28);
output(5, 44) <= input(29);
output(5, 45) <= input(30);
output(5, 46) <= input(31);
output(5, 47) <= input(33);
output(5, 48) <= input(2);
output(5, 49) <= input(3);
output(5, 50) <= input(4);
output(5, 51) <= input(5);
output(5, 52) <= input(6);
output(5, 53) <= input(7);
output(5, 54) <= input(8);
output(5, 55) <= input(9);
output(5, 56) <= input(10);
output(5, 57) <= input(11);
output(5, 58) <= input(12);
output(5, 59) <= input(13);
output(5, 60) <= input(14);
output(5, 61) <= input(15);
output(5, 62) <= input(32);
output(5, 63) <= input(34);
output(5, 64) <= input(18);
output(5, 65) <= input(19);
output(5, 66) <= input(20);
output(5, 67) <= input(21);
output(5, 68) <= input(22);
output(5, 69) <= input(23);
output(5, 70) <= input(24);
output(5, 71) <= input(25);
output(5, 72) <= input(26);
output(5, 73) <= input(27);
output(5, 74) <= input(28);
output(5, 75) <= input(29);
output(5, 76) <= input(30);
output(5, 77) <= input(31);
output(5, 78) <= input(33);
output(5, 79) <= input(35);
output(5, 80) <= input(3);
output(5, 81) <= input(4);
output(5, 82) <= input(5);
output(5, 83) <= input(6);
output(5, 84) <= input(7);
output(5, 85) <= input(8);
output(5, 86) <= input(9);
output(5, 87) <= input(10);
output(5, 88) <= input(11);
output(5, 89) <= input(12);
output(5, 90) <= input(13);
output(5, 91) <= input(14);
output(5, 92) <= input(15);
output(5, 93) <= input(32);
output(5, 94) <= input(34);
output(5, 95) <= input(36);
output(5, 96) <= input(19);
output(5, 97) <= input(20);
output(5, 98) <= input(21);
output(5, 99) <= input(22);
output(5, 100) <= input(23);
output(5, 101) <= input(24);
output(5, 102) <= input(25);
output(5, 103) <= input(26);
output(5, 104) <= input(27);
output(5, 105) <= input(28);
output(5, 106) <= input(29);
output(5, 107) <= input(30);
output(5, 108) <= input(31);
output(5, 109) <= input(33);
output(5, 110) <= input(35);
output(5, 111) <= input(37);
output(5, 112) <= input(4);
output(5, 113) <= input(5);
output(5, 114) <= input(6);
output(5, 115) <= input(7);
output(5, 116) <= input(8);
output(5, 117) <= input(9);
output(5, 118) <= input(10);
output(5, 119) <= input(11);
output(5, 120) <= input(12);
output(5, 121) <= input(13);
output(5, 122) <= input(14);
output(5, 123) <= input(15);
output(5, 124) <= input(32);
output(5, 125) <= input(34);
output(5, 126) <= input(36);
output(5, 127) <= input(38);
output(5, 128) <= input(20);
output(5, 129) <= input(21);
output(5, 130) <= input(22);
output(5, 131) <= input(23);
output(5, 132) <= input(24);
output(5, 133) <= input(25);
output(5, 134) <= input(26);
output(5, 135) <= input(27);
output(5, 136) <= input(28);
output(5, 137) <= input(29);
output(5, 138) <= input(30);
output(5, 139) <= input(31);
output(5, 140) <= input(33);
output(5, 141) <= input(35);
output(5, 142) <= input(37);
output(5, 143) <= input(39);
output(5, 144) <= input(5);
output(5, 145) <= input(6);
output(5, 146) <= input(7);
output(5, 147) <= input(8);
output(5, 148) <= input(9);
output(5, 149) <= input(10);
output(5, 150) <= input(11);
output(5, 151) <= input(12);
output(5, 152) <= input(13);
output(5, 153) <= input(14);
output(5, 154) <= input(15);
output(5, 155) <= input(32);
output(5, 156) <= input(34);
output(5, 157) <= input(36);
output(5, 158) <= input(38);
output(5, 159) <= input(40);
output(5, 160) <= input(21);
output(5, 161) <= input(22);
output(5, 162) <= input(23);
output(5, 163) <= input(24);
output(5, 164) <= input(25);
output(5, 165) <= input(26);
output(5, 166) <= input(27);
output(5, 167) <= input(28);
output(5, 168) <= input(29);
output(5, 169) <= input(30);
output(5, 170) <= input(31);
output(5, 171) <= input(33);
output(5, 172) <= input(35);
output(5, 173) <= input(37);
output(5, 174) <= input(39);
output(5, 175) <= input(41);
output(5, 176) <= input(6);
output(5, 177) <= input(7);
output(5, 178) <= input(8);
output(5, 179) <= input(9);
output(5, 180) <= input(10);
output(5, 181) <= input(11);
output(5, 182) <= input(12);
output(5, 183) <= input(13);
output(5, 184) <= input(14);
output(5, 185) <= input(15);
output(5, 186) <= input(32);
output(5, 187) <= input(34);
output(5, 188) <= input(36);
output(5, 189) <= input(38);
output(5, 190) <= input(40);
output(5, 191) <= input(42);
output(5, 192) <= input(22);
output(5, 193) <= input(23);
output(5, 194) <= input(24);
output(5, 195) <= input(25);
output(5, 196) <= input(26);
output(5, 197) <= input(27);
output(5, 198) <= input(28);
output(5, 199) <= input(29);
output(5, 200) <= input(30);
output(5, 201) <= input(31);
output(5, 202) <= input(33);
output(5, 203) <= input(35);
output(5, 204) <= input(37);
output(5, 205) <= input(39);
output(5, 206) <= input(41);
output(5, 207) <= input(43);
output(5, 208) <= input(7);
output(5, 209) <= input(8);
output(5, 210) <= input(9);
output(5, 211) <= input(10);
output(5, 212) <= input(11);
output(5, 213) <= input(12);
output(5, 214) <= input(13);
output(5, 215) <= input(14);
output(5, 216) <= input(15);
output(5, 217) <= input(32);
output(5, 218) <= input(34);
output(5, 219) <= input(36);
output(5, 220) <= input(38);
output(5, 221) <= input(40);
output(5, 222) <= input(42);
output(5, 223) <= input(44);
output(5, 224) <= input(23);
output(5, 225) <= input(24);
output(5, 226) <= input(25);
output(5, 227) <= input(26);
output(5, 228) <= input(27);
output(5, 229) <= input(28);
output(5, 230) <= input(29);
output(5, 231) <= input(30);
output(5, 232) <= input(31);
output(5, 233) <= input(33);
output(5, 234) <= input(35);
output(5, 235) <= input(37);
output(5, 236) <= input(39);
output(5, 237) <= input(41);
output(5, 238) <= input(43);
output(5, 239) <= input(45);
output(5, 240) <= input(8);
output(5, 241) <= input(9);
output(5, 242) <= input(10);
output(5, 243) <= input(11);
output(5, 244) <= input(12);
output(5, 245) <= input(13);
output(5, 246) <= input(14);
output(5, 247) <= input(15);
output(5, 248) <= input(32);
output(5, 249) <= input(34);
output(5, 250) <= input(36);
output(5, 251) <= input(38);
output(5, 252) <= input(40);
output(5, 253) <= input(42);
output(5, 254) <= input(44);
output(5, 255) <= input(46);
when "1111" =>
output(0, 0) <= input(0);
output(0, 1) <= input(1);
output(0, 2) <= input(2);
output(0, 3) <= input(3);
output(0, 4) <= input(4);
output(0, 5) <= input(5);
output(0, 6) <= input(6);
output(0, 7) <= input(7);
output(0, 8) <= input(8);
output(0, 9) <= input(9);
output(0, 10) <= input(10);
output(0, 11) <= input(11);
output(0, 12) <= input(12);
output(0, 13) <= input(13);
output(0, 14) <= input(14);
output(0, 15) <= input(15);
output(0, 16) <= input(16);
output(0, 17) <= input(17);
output(0, 18) <= input(18);
output(0, 19) <= input(19);
output(0, 20) <= input(20);
output(0, 21) <= input(21);
output(0, 22) <= input(22);
output(0, 23) <= input(23);
output(0, 24) <= input(24);
output(0, 25) <= input(25);
output(0, 26) <= input(26);
output(0, 27) <= input(27);
output(0, 28) <= input(28);
output(0, 29) <= input(29);
output(0, 30) <= input(30);
output(0, 31) <= input(31);
output(0, 32) <= input(1);
output(0, 33) <= input(2);
output(0, 34) <= input(3);
output(0, 35) <= input(4);
output(0, 36) <= input(5);
output(0, 37) <= input(6);
output(0, 38) <= input(7);
output(0, 39) <= input(8);
output(0, 40) <= input(9);
output(0, 41) <= input(10);
output(0, 42) <= input(11);
output(0, 43) <= input(12);
output(0, 44) <= input(13);
output(0, 45) <= input(14);
output(0, 46) <= input(15);
output(0, 47) <= input(32);
output(0, 48) <= input(17);
output(0, 49) <= input(18);
output(0, 50) <= input(19);
output(0, 51) <= input(20);
output(0, 52) <= input(21);
output(0, 53) <= input(22);
output(0, 54) <= input(23);
output(0, 55) <= input(24);
output(0, 56) <= input(25);
output(0, 57) <= input(26);
output(0, 58) <= input(27);
output(0, 59) <= input(28);
output(0, 60) <= input(29);
output(0, 61) <= input(30);
output(0, 62) <= input(31);
output(0, 63) <= input(33);
output(0, 64) <= input(2);
output(0, 65) <= input(3);
output(0, 66) <= input(4);
output(0, 67) <= input(5);
output(0, 68) <= input(6);
output(0, 69) <= input(7);
output(0, 70) <= input(8);
output(0, 71) <= input(9);
output(0, 72) <= input(10);
output(0, 73) <= input(11);
output(0, 74) <= input(12);
output(0, 75) <= input(13);
output(0, 76) <= input(14);
output(0, 77) <= input(15);
output(0, 78) <= input(32);
output(0, 79) <= input(34);
output(0, 80) <= input(18);
output(0, 81) <= input(19);
output(0, 82) <= input(20);
output(0, 83) <= input(21);
output(0, 84) <= input(22);
output(0, 85) <= input(23);
output(0, 86) <= input(24);
output(0, 87) <= input(25);
output(0, 88) <= input(26);
output(0, 89) <= input(27);
output(0, 90) <= input(28);
output(0, 91) <= input(29);
output(0, 92) <= input(30);
output(0, 93) <= input(31);
output(0, 94) <= input(33);
output(0, 95) <= input(35);
output(0, 96) <= input(3);
output(0, 97) <= input(4);
output(0, 98) <= input(5);
output(0, 99) <= input(6);
output(0, 100) <= input(7);
output(0, 101) <= input(8);
output(0, 102) <= input(9);
output(0, 103) <= input(10);
output(0, 104) <= input(11);
output(0, 105) <= input(12);
output(0, 106) <= input(13);
output(0, 107) <= input(14);
output(0, 108) <= input(15);
output(0, 109) <= input(32);
output(0, 110) <= input(34);
output(0, 111) <= input(36);
output(0, 112) <= input(4);
output(0, 113) <= input(5);
output(0, 114) <= input(6);
output(0, 115) <= input(7);
output(0, 116) <= input(8);
output(0, 117) <= input(9);
output(0, 118) <= input(10);
output(0, 119) <= input(11);
output(0, 120) <= input(12);
output(0, 121) <= input(13);
output(0, 122) <= input(14);
output(0, 123) <= input(15);
output(0, 124) <= input(32);
output(0, 125) <= input(34);
output(0, 126) <= input(36);
output(0, 127) <= input(37);
output(0, 128) <= input(20);
output(0, 129) <= input(21);
output(0, 130) <= input(22);
output(0, 131) <= input(23);
output(0, 132) <= input(24);
output(0, 133) <= input(25);
output(0, 134) <= input(26);
output(0, 135) <= input(27);
output(0, 136) <= input(28);
output(0, 137) <= input(29);
output(0, 138) <= input(30);
output(0, 139) <= input(31);
output(0, 140) <= input(33);
output(0, 141) <= input(35);
output(0, 142) <= input(38);
output(0, 143) <= input(39);
output(0, 144) <= input(5);
output(0, 145) <= input(6);
output(0, 146) <= input(7);
output(0, 147) <= input(8);
output(0, 148) <= input(9);
output(0, 149) <= input(10);
output(0, 150) <= input(11);
output(0, 151) <= input(12);
output(0, 152) <= input(13);
output(0, 153) <= input(14);
output(0, 154) <= input(15);
output(0, 155) <= input(32);
output(0, 156) <= input(34);
output(0, 157) <= input(36);
output(0, 158) <= input(37);
output(0, 159) <= input(40);
output(0, 160) <= input(21);
output(0, 161) <= input(22);
output(0, 162) <= input(23);
output(0, 163) <= input(24);
output(0, 164) <= input(25);
output(0, 165) <= input(26);
output(0, 166) <= input(27);
output(0, 167) <= input(28);
output(0, 168) <= input(29);
output(0, 169) <= input(30);
output(0, 170) <= input(31);
output(0, 171) <= input(33);
output(0, 172) <= input(35);
output(0, 173) <= input(38);
output(0, 174) <= input(39);
output(0, 175) <= input(41);
output(0, 176) <= input(6);
output(0, 177) <= input(7);
output(0, 178) <= input(8);
output(0, 179) <= input(9);
output(0, 180) <= input(10);
output(0, 181) <= input(11);
output(0, 182) <= input(12);
output(0, 183) <= input(13);
output(0, 184) <= input(14);
output(0, 185) <= input(15);
output(0, 186) <= input(32);
output(0, 187) <= input(34);
output(0, 188) <= input(36);
output(0, 189) <= input(37);
output(0, 190) <= input(40);
output(0, 191) <= input(42);
output(0, 192) <= input(22);
output(0, 193) <= input(23);
output(0, 194) <= input(24);
output(0, 195) <= input(25);
output(0, 196) <= input(26);
output(0, 197) <= input(27);
output(0, 198) <= input(28);
output(0, 199) <= input(29);
output(0, 200) <= input(30);
output(0, 201) <= input(31);
output(0, 202) <= input(33);
output(0, 203) <= input(35);
output(0, 204) <= input(38);
output(0, 205) <= input(39);
output(0, 206) <= input(41);
output(0, 207) <= input(43);
output(0, 208) <= input(7);
output(0, 209) <= input(8);
output(0, 210) <= input(9);
output(0, 211) <= input(10);
output(0, 212) <= input(11);
output(0, 213) <= input(12);
output(0, 214) <= input(13);
output(0, 215) <= input(14);
output(0, 216) <= input(15);
output(0, 217) <= input(32);
output(0, 218) <= input(34);
output(0, 219) <= input(36);
output(0, 220) <= input(37);
output(0, 221) <= input(40);
output(0, 222) <= input(42);
output(0, 223) <= input(44);
output(0, 224) <= input(23);
output(0, 225) <= input(24);
output(0, 226) <= input(25);
output(0, 227) <= input(26);
output(0, 228) <= input(27);
output(0, 229) <= input(28);
output(0, 230) <= input(29);
output(0, 231) <= input(30);
output(0, 232) <= input(31);
output(0, 233) <= input(33);
output(0, 234) <= input(35);
output(0, 235) <= input(38);
output(0, 236) <= input(39);
output(0, 237) <= input(41);
output(0, 238) <= input(43);
output(0, 239) <= input(45);
output(0, 240) <= input(24);
output(0, 241) <= input(25);
output(0, 242) <= input(26);
output(0, 243) <= input(27);
output(0, 244) <= input(28);
output(0, 245) <= input(29);
output(0, 246) <= input(30);
output(0, 247) <= input(31);
output(0, 248) <= input(33);
output(0, 249) <= input(35);
output(0, 250) <= input(38);
output(0, 251) <= input(39);
output(0, 252) <= input(41);
output(0, 253) <= input(43);
output(0, 254) <= input(45);
output(0, 255) <= input(46);
output(1, 0) <= input(0);
output(1, 1) <= input(1);
output(1, 2) <= input(2);
output(1, 3) <= input(3);
output(1, 4) <= input(4);
output(1, 5) <= input(5);
output(1, 6) <= input(6);
output(1, 7) <= input(7);
output(1, 8) <= input(8);
output(1, 9) <= input(9);
output(1, 10) <= input(10);
output(1, 11) <= input(11);
output(1, 12) <= input(12);
output(1, 13) <= input(13);
output(1, 14) <= input(14);
output(1, 15) <= input(15);
output(1, 16) <= input(16);
output(1, 17) <= input(17);
output(1, 18) <= input(18);
output(1, 19) <= input(19);
output(1, 20) <= input(20);
output(1, 21) <= input(21);
output(1, 22) <= input(22);
output(1, 23) <= input(23);
output(1, 24) <= input(24);
output(1, 25) <= input(25);
output(1, 26) <= input(26);
output(1, 27) <= input(27);
output(1, 28) <= input(28);
output(1, 29) <= input(29);
output(1, 30) <= input(30);
output(1, 31) <= input(31);
output(1, 32) <= input(1);
output(1, 33) <= input(2);
output(1, 34) <= input(3);
output(1, 35) <= input(4);
output(1, 36) <= input(5);
output(1, 37) <= input(6);
output(1, 38) <= input(7);
output(1, 39) <= input(8);
output(1, 40) <= input(9);
output(1, 41) <= input(10);
output(1, 42) <= input(11);
output(1, 43) <= input(12);
output(1, 44) <= input(13);
output(1, 45) <= input(14);
output(1, 46) <= input(15);
output(1, 47) <= input(32);
output(1, 48) <= input(2);
output(1, 49) <= input(3);
output(1, 50) <= input(4);
output(1, 51) <= input(5);
output(1, 52) <= input(6);
output(1, 53) <= input(7);
output(1, 54) <= input(8);
output(1, 55) <= input(9);
output(1, 56) <= input(10);
output(1, 57) <= input(11);
output(1, 58) <= input(12);
output(1, 59) <= input(13);
output(1, 60) <= input(14);
output(1, 61) <= input(15);
output(1, 62) <= input(32);
output(1, 63) <= input(34);
output(1, 64) <= input(18);
output(1, 65) <= input(19);
output(1, 66) <= input(20);
output(1, 67) <= input(21);
output(1, 68) <= input(22);
output(1, 69) <= input(23);
output(1, 70) <= input(24);
output(1, 71) <= input(25);
output(1, 72) <= input(26);
output(1, 73) <= input(27);
output(1, 74) <= input(28);
output(1, 75) <= input(29);
output(1, 76) <= input(30);
output(1, 77) <= input(31);
output(1, 78) <= input(33);
output(1, 79) <= input(35);
output(1, 80) <= input(3);
output(1, 81) <= input(4);
output(1, 82) <= input(5);
output(1, 83) <= input(6);
output(1, 84) <= input(7);
output(1, 85) <= input(8);
output(1, 86) <= input(9);
output(1, 87) <= input(10);
output(1, 88) <= input(11);
output(1, 89) <= input(12);
output(1, 90) <= input(13);
output(1, 91) <= input(14);
output(1, 92) <= input(15);
output(1, 93) <= input(32);
output(1, 94) <= input(34);
output(1, 95) <= input(36);
output(1, 96) <= input(19);
output(1, 97) <= input(20);
output(1, 98) <= input(21);
output(1, 99) <= input(22);
output(1, 100) <= input(23);
output(1, 101) <= input(24);
output(1, 102) <= input(25);
output(1, 103) <= input(26);
output(1, 104) <= input(27);
output(1, 105) <= input(28);
output(1, 106) <= input(29);
output(1, 107) <= input(30);
output(1, 108) <= input(31);
output(1, 109) <= input(33);
output(1, 110) <= input(35);
output(1, 111) <= input(38);
output(1, 112) <= input(20);
output(1, 113) <= input(21);
output(1, 114) <= input(22);
output(1, 115) <= input(23);
output(1, 116) <= input(24);
output(1, 117) <= input(25);
output(1, 118) <= input(26);
output(1, 119) <= input(27);
output(1, 120) <= input(28);
output(1, 121) <= input(29);
output(1, 122) <= input(30);
output(1, 123) <= input(31);
output(1, 124) <= input(33);
output(1, 125) <= input(35);
output(1, 126) <= input(38);
output(1, 127) <= input(39);
output(1, 128) <= input(5);
output(1, 129) <= input(6);
output(1, 130) <= input(7);
output(1, 131) <= input(8);
output(1, 132) <= input(9);
output(1, 133) <= input(10);
output(1, 134) <= input(11);
output(1, 135) <= input(12);
output(1, 136) <= input(13);
output(1, 137) <= input(14);
output(1, 138) <= input(15);
output(1, 139) <= input(32);
output(1, 140) <= input(34);
output(1, 141) <= input(36);
output(1, 142) <= input(37);
output(1, 143) <= input(40);
output(1, 144) <= input(21);
output(1, 145) <= input(22);
output(1, 146) <= input(23);
output(1, 147) <= input(24);
output(1, 148) <= input(25);
output(1, 149) <= input(26);
output(1, 150) <= input(27);
output(1, 151) <= input(28);
output(1, 152) <= input(29);
output(1, 153) <= input(30);
output(1, 154) <= input(31);
output(1, 155) <= input(33);
output(1, 156) <= input(35);
output(1, 157) <= input(38);
output(1, 158) <= input(39);
output(1, 159) <= input(41);
output(1, 160) <= input(6);
output(1, 161) <= input(7);
output(1, 162) <= input(8);
output(1, 163) <= input(9);
output(1, 164) <= input(10);
output(1, 165) <= input(11);
output(1, 166) <= input(12);
output(1, 167) <= input(13);
output(1, 168) <= input(14);
output(1, 169) <= input(15);
output(1, 170) <= input(32);
output(1, 171) <= input(34);
output(1, 172) <= input(36);
output(1, 173) <= input(37);
output(1, 174) <= input(40);
output(1, 175) <= input(42);
output(1, 176) <= input(7);
output(1, 177) <= input(8);
output(1, 178) <= input(9);
output(1, 179) <= input(10);
output(1, 180) <= input(11);
output(1, 181) <= input(12);
output(1, 182) <= input(13);
output(1, 183) <= input(14);
output(1, 184) <= input(15);
output(1, 185) <= input(32);
output(1, 186) <= input(34);
output(1, 187) <= input(36);
output(1, 188) <= input(37);
output(1, 189) <= input(40);
output(1, 190) <= input(42);
output(1, 191) <= input(44);
output(1, 192) <= input(23);
output(1, 193) <= input(24);
output(1, 194) <= input(25);
output(1, 195) <= input(26);
output(1, 196) <= input(27);
output(1, 197) <= input(28);
output(1, 198) <= input(29);
output(1, 199) <= input(30);
output(1, 200) <= input(31);
output(1, 201) <= input(33);
output(1, 202) <= input(35);
output(1, 203) <= input(38);
output(1, 204) <= input(39);
output(1, 205) <= input(41);
output(1, 206) <= input(43);
output(1, 207) <= input(45);
output(1, 208) <= input(8);
output(1, 209) <= input(9);
output(1, 210) <= input(10);
output(1, 211) <= input(11);
output(1, 212) <= input(12);
output(1, 213) <= input(13);
output(1, 214) <= input(14);
output(1, 215) <= input(15);
output(1, 216) <= input(32);
output(1, 217) <= input(34);
output(1, 218) <= input(36);
output(1, 219) <= input(37);
output(1, 220) <= input(40);
output(1, 221) <= input(42);
output(1, 222) <= input(44);
output(1, 223) <= input(47);
output(1, 224) <= input(24);
output(1, 225) <= input(25);
output(1, 226) <= input(26);
output(1, 227) <= input(27);
output(1, 228) <= input(28);
output(1, 229) <= input(29);
output(1, 230) <= input(30);
output(1, 231) <= input(31);
output(1, 232) <= input(33);
output(1, 233) <= input(35);
output(1, 234) <= input(38);
output(1, 235) <= input(39);
output(1, 236) <= input(41);
output(1, 237) <= input(43);
output(1, 238) <= input(45);
output(1, 239) <= input(46);
output(1, 240) <= input(25);
output(1, 241) <= input(26);
output(1, 242) <= input(27);
output(1, 243) <= input(28);
output(1, 244) <= input(29);
output(1, 245) <= input(30);
output(1, 246) <= input(31);
output(1, 247) <= input(33);
output(1, 248) <= input(35);
output(1, 249) <= input(38);
output(1, 250) <= input(39);
output(1, 251) <= input(41);
output(1, 252) <= input(43);
output(1, 253) <= input(45);
output(1, 254) <= input(46);
output(1, 255) <= input(48);
output(2, 0) <= input(0);
output(2, 1) <= input(1);
output(2, 2) <= input(2);
output(2, 3) <= input(3);
output(2, 4) <= input(4);
output(2, 5) <= input(5);
output(2, 6) <= input(6);
output(2, 7) <= input(7);
output(2, 8) <= input(8);
output(2, 9) <= input(9);
output(2, 10) <= input(10);
output(2, 11) <= input(11);
output(2, 12) <= input(12);
output(2, 13) <= input(13);
output(2, 14) <= input(14);
output(2, 15) <= input(15);
output(2, 16) <= input(16);
output(2, 17) <= input(17);
output(2, 18) <= input(18);
output(2, 19) <= input(19);
output(2, 20) <= input(20);
output(2, 21) <= input(21);
output(2, 22) <= input(22);
output(2, 23) <= input(23);
output(2, 24) <= input(24);
output(2, 25) <= input(25);
output(2, 26) <= input(26);
output(2, 27) <= input(27);
output(2, 28) <= input(28);
output(2, 29) <= input(29);
output(2, 30) <= input(30);
output(2, 31) <= input(31);
output(2, 32) <= input(17);
output(2, 33) <= input(18);
output(2, 34) <= input(19);
output(2, 35) <= input(20);
output(2, 36) <= input(21);
output(2, 37) <= input(22);
output(2, 38) <= input(23);
output(2, 39) <= input(24);
output(2, 40) <= input(25);
output(2, 41) <= input(26);
output(2, 42) <= input(27);
output(2, 43) <= input(28);
output(2, 44) <= input(29);
output(2, 45) <= input(30);
output(2, 46) <= input(31);
output(2, 47) <= input(33);
output(2, 48) <= input(2);
output(2, 49) <= input(3);
output(2, 50) <= input(4);
output(2, 51) <= input(5);
output(2, 52) <= input(6);
output(2, 53) <= input(7);
output(2, 54) <= input(8);
output(2, 55) <= input(9);
output(2, 56) <= input(10);
output(2, 57) <= input(11);
output(2, 58) <= input(12);
output(2, 59) <= input(13);
output(2, 60) <= input(14);
output(2, 61) <= input(15);
output(2, 62) <= input(32);
output(2, 63) <= input(34);
output(2, 64) <= input(3);
output(2, 65) <= input(4);
output(2, 66) <= input(5);
output(2, 67) <= input(6);
output(2, 68) <= input(7);
output(2, 69) <= input(8);
output(2, 70) <= input(9);
output(2, 71) <= input(10);
output(2, 72) <= input(11);
output(2, 73) <= input(12);
output(2, 74) <= input(13);
output(2, 75) <= input(14);
output(2, 76) <= input(15);
output(2, 77) <= input(32);
output(2, 78) <= input(34);
output(2, 79) <= input(36);
output(2, 80) <= input(19);
output(2, 81) <= input(20);
output(2, 82) <= input(21);
output(2, 83) <= input(22);
output(2, 84) <= input(23);
output(2, 85) <= input(24);
output(2, 86) <= input(25);
output(2, 87) <= input(26);
output(2, 88) <= input(27);
output(2, 89) <= input(28);
output(2, 90) <= input(29);
output(2, 91) <= input(30);
output(2, 92) <= input(31);
output(2, 93) <= input(33);
output(2, 94) <= input(35);
output(2, 95) <= input(38);
output(2, 96) <= input(20);
output(2, 97) <= input(21);
output(2, 98) <= input(22);
output(2, 99) <= input(23);
output(2, 100) <= input(24);
output(2, 101) <= input(25);
output(2, 102) <= input(26);
output(2, 103) <= input(27);
output(2, 104) <= input(28);
output(2, 105) <= input(29);
output(2, 106) <= input(30);
output(2, 107) <= input(31);
output(2, 108) <= input(33);
output(2, 109) <= input(35);
output(2, 110) <= input(38);
output(2, 111) <= input(39);
output(2, 112) <= input(5);
output(2, 113) <= input(6);
output(2, 114) <= input(7);
output(2, 115) <= input(8);
output(2, 116) <= input(9);
output(2, 117) <= input(10);
output(2, 118) <= input(11);
output(2, 119) <= input(12);
output(2, 120) <= input(13);
output(2, 121) <= input(14);
output(2, 122) <= input(15);
output(2, 123) <= input(32);
output(2, 124) <= input(34);
output(2, 125) <= input(36);
output(2, 126) <= input(37);
output(2, 127) <= input(40);
output(2, 128) <= input(21);
output(2, 129) <= input(22);
output(2, 130) <= input(23);
output(2, 131) <= input(24);
output(2, 132) <= input(25);
output(2, 133) <= input(26);
output(2, 134) <= input(27);
output(2, 135) <= input(28);
output(2, 136) <= input(29);
output(2, 137) <= input(30);
output(2, 138) <= input(31);
output(2, 139) <= input(33);
output(2, 140) <= input(35);
output(2, 141) <= input(38);
output(2, 142) <= input(39);
output(2, 143) <= input(41);
output(2, 144) <= input(22);
output(2, 145) <= input(23);
output(2, 146) <= input(24);
output(2, 147) <= input(25);
output(2, 148) <= input(26);
output(2, 149) <= input(27);
output(2, 150) <= input(28);
output(2, 151) <= input(29);
output(2, 152) <= input(30);
output(2, 153) <= input(31);
output(2, 154) <= input(33);
output(2, 155) <= input(35);
output(2, 156) <= input(38);
output(2, 157) <= input(39);
output(2, 158) <= input(41);
output(2, 159) <= input(43);
output(2, 160) <= input(7);
output(2, 161) <= input(8);
output(2, 162) <= input(9);
output(2, 163) <= input(10);
output(2, 164) <= input(11);
output(2, 165) <= input(12);
output(2, 166) <= input(13);
output(2, 167) <= input(14);
output(2, 168) <= input(15);
output(2, 169) <= input(32);
output(2, 170) <= input(34);
output(2, 171) <= input(36);
output(2, 172) <= input(37);
output(2, 173) <= input(40);
output(2, 174) <= input(42);
output(2, 175) <= input(44);
output(2, 176) <= input(8);
output(2, 177) <= input(9);
output(2, 178) <= input(10);
output(2, 179) <= input(11);
output(2, 180) <= input(12);
output(2, 181) <= input(13);
output(2, 182) <= input(14);
output(2, 183) <= input(15);
output(2, 184) <= input(32);
output(2, 185) <= input(34);
output(2, 186) <= input(36);
output(2, 187) <= input(37);
output(2, 188) <= input(40);
output(2, 189) <= input(42);
output(2, 190) <= input(44);
output(2, 191) <= input(47);
output(2, 192) <= input(24);
output(2, 193) <= input(25);
output(2, 194) <= input(26);
output(2, 195) <= input(27);
output(2, 196) <= input(28);
output(2, 197) <= input(29);
output(2, 198) <= input(30);
output(2, 199) <= input(31);
output(2, 200) <= input(33);
output(2, 201) <= input(35);
output(2, 202) <= input(38);
output(2, 203) <= input(39);
output(2, 204) <= input(41);
output(2, 205) <= input(43);
output(2, 206) <= input(45);
output(2, 207) <= input(46);
output(2, 208) <= input(25);
output(2, 209) <= input(26);
output(2, 210) <= input(27);
output(2, 211) <= input(28);
output(2, 212) <= input(29);
output(2, 213) <= input(30);
output(2, 214) <= input(31);
output(2, 215) <= input(33);
output(2, 216) <= input(35);
output(2, 217) <= input(38);
output(2, 218) <= input(39);
output(2, 219) <= input(41);
output(2, 220) <= input(43);
output(2, 221) <= input(45);
output(2, 222) <= input(46);
output(2, 223) <= input(48);
output(2, 224) <= input(10);
output(2, 225) <= input(11);
output(2, 226) <= input(12);
output(2, 227) <= input(13);
output(2, 228) <= input(14);
output(2, 229) <= input(15);
output(2, 230) <= input(32);
output(2, 231) <= input(34);
output(2, 232) <= input(36);
output(2, 233) <= input(37);
output(2, 234) <= input(40);
output(2, 235) <= input(42);
output(2, 236) <= input(44);
output(2, 237) <= input(47);
output(2, 238) <= input(49);
output(2, 239) <= input(50);
output(2, 240) <= input(11);
output(2, 241) <= input(12);
output(2, 242) <= input(13);
output(2, 243) <= input(14);
output(2, 244) <= input(15);
output(2, 245) <= input(32);
output(2, 246) <= input(34);
output(2, 247) <= input(36);
output(2, 248) <= input(37);
output(2, 249) <= input(40);
output(2, 250) <= input(42);
output(2, 251) <= input(44);
output(2, 252) <= input(47);
output(2, 253) <= input(49);
output(2, 254) <= input(50);
output(2, 255) <= input(51);
output(3, 0) <= input(0);
output(3, 1) <= input(1);
output(3, 2) <= input(2);
output(3, 3) <= input(3);
output(3, 4) <= input(4);
output(3, 5) <= input(5);
output(3, 6) <= input(6);
output(3, 7) <= input(7);
output(3, 8) <= input(8);
output(3, 9) <= input(9);
output(3, 10) <= input(10);
output(3, 11) <= input(11);
output(3, 12) <= input(12);
output(3, 13) <= input(13);
output(3, 14) <= input(14);
output(3, 15) <= input(15);
output(3, 16) <= input(1);
output(3, 17) <= input(2);
output(3, 18) <= input(3);
output(3, 19) <= input(4);
output(3, 20) <= input(5);
output(3, 21) <= input(6);
output(3, 22) <= input(7);
output(3, 23) <= input(8);
output(3, 24) <= input(9);
output(3, 25) <= input(10);
output(3, 26) <= input(11);
output(3, 27) <= input(12);
output(3, 28) <= input(13);
output(3, 29) <= input(14);
output(3, 30) <= input(15);
output(3, 31) <= input(32);
output(3, 32) <= input(17);
output(3, 33) <= input(18);
output(3, 34) <= input(19);
output(3, 35) <= input(20);
output(3, 36) <= input(21);
output(3, 37) <= input(22);
output(3, 38) <= input(23);
output(3, 39) <= input(24);
output(3, 40) <= input(25);
output(3, 41) <= input(26);
output(3, 42) <= input(27);
output(3, 43) <= input(28);
output(3, 44) <= input(29);
output(3, 45) <= input(30);
output(3, 46) <= input(31);
output(3, 47) <= input(33);
output(3, 48) <= input(18);
output(3, 49) <= input(19);
output(3, 50) <= input(20);
output(3, 51) <= input(21);
output(3, 52) <= input(22);
output(3, 53) <= input(23);
output(3, 54) <= input(24);
output(3, 55) <= input(25);
output(3, 56) <= input(26);
output(3, 57) <= input(27);
output(3, 58) <= input(28);
output(3, 59) <= input(29);
output(3, 60) <= input(30);
output(3, 61) <= input(31);
output(3, 62) <= input(33);
output(3, 63) <= input(35);
output(3, 64) <= input(19);
output(3, 65) <= input(20);
output(3, 66) <= input(21);
output(3, 67) <= input(22);
output(3, 68) <= input(23);
output(3, 69) <= input(24);
output(3, 70) <= input(25);
output(3, 71) <= input(26);
output(3, 72) <= input(27);
output(3, 73) <= input(28);
output(3, 74) <= input(29);
output(3, 75) <= input(30);
output(3, 76) <= input(31);
output(3, 77) <= input(33);
output(3, 78) <= input(35);
output(3, 79) <= input(38);
output(3, 80) <= input(4);
output(3, 81) <= input(5);
output(3, 82) <= input(6);
output(3, 83) <= input(7);
output(3, 84) <= input(8);
output(3, 85) <= input(9);
output(3, 86) <= input(10);
output(3, 87) <= input(11);
output(3, 88) <= input(12);
output(3, 89) <= input(13);
output(3, 90) <= input(14);
output(3, 91) <= input(15);
output(3, 92) <= input(32);
output(3, 93) <= input(34);
output(3, 94) <= input(36);
output(3, 95) <= input(37);
output(3, 96) <= input(5);
output(3, 97) <= input(6);
output(3, 98) <= input(7);
output(3, 99) <= input(8);
output(3, 100) <= input(9);
output(3, 101) <= input(10);
output(3, 102) <= input(11);
output(3, 103) <= input(12);
output(3, 104) <= input(13);
output(3, 105) <= input(14);
output(3, 106) <= input(15);
output(3, 107) <= input(32);
output(3, 108) <= input(34);
output(3, 109) <= input(36);
output(3, 110) <= input(37);
output(3, 111) <= input(40);
output(3, 112) <= input(6);
output(3, 113) <= input(7);
output(3, 114) <= input(8);
output(3, 115) <= input(9);
output(3, 116) <= input(10);
output(3, 117) <= input(11);
output(3, 118) <= input(12);
output(3, 119) <= input(13);
output(3, 120) <= input(14);
output(3, 121) <= input(15);
output(3, 122) <= input(32);
output(3, 123) <= input(34);
output(3, 124) <= input(36);
output(3, 125) <= input(37);
output(3, 126) <= input(40);
output(3, 127) <= input(42);
output(3, 128) <= input(22);
output(3, 129) <= input(23);
output(3, 130) <= input(24);
output(3, 131) <= input(25);
output(3, 132) <= input(26);
output(3, 133) <= input(27);
output(3, 134) <= input(28);
output(3, 135) <= input(29);
output(3, 136) <= input(30);
output(3, 137) <= input(31);
output(3, 138) <= input(33);
output(3, 139) <= input(35);
output(3, 140) <= input(38);
output(3, 141) <= input(39);
output(3, 142) <= input(41);
output(3, 143) <= input(43);
output(3, 144) <= input(23);
output(3, 145) <= input(24);
output(3, 146) <= input(25);
output(3, 147) <= input(26);
output(3, 148) <= input(27);
output(3, 149) <= input(28);
output(3, 150) <= input(29);
output(3, 151) <= input(30);
output(3, 152) <= input(31);
output(3, 153) <= input(33);
output(3, 154) <= input(35);
output(3, 155) <= input(38);
output(3, 156) <= input(39);
output(3, 157) <= input(41);
output(3, 158) <= input(43);
output(3, 159) <= input(45);
output(3, 160) <= input(8);
output(3, 161) <= input(9);
output(3, 162) <= input(10);
output(3, 163) <= input(11);
output(3, 164) <= input(12);
output(3, 165) <= input(13);
output(3, 166) <= input(14);
output(3, 167) <= input(15);
output(3, 168) <= input(32);
output(3, 169) <= input(34);
output(3, 170) <= input(36);
output(3, 171) <= input(37);
output(3, 172) <= input(40);
output(3, 173) <= input(42);
output(3, 174) <= input(44);
output(3, 175) <= input(47);
output(3, 176) <= input(9);
output(3, 177) <= input(10);
output(3, 178) <= input(11);
output(3, 179) <= input(12);
output(3, 180) <= input(13);
output(3, 181) <= input(14);
output(3, 182) <= input(15);
output(3, 183) <= input(32);
output(3, 184) <= input(34);
output(3, 185) <= input(36);
output(3, 186) <= input(37);
output(3, 187) <= input(40);
output(3, 188) <= input(42);
output(3, 189) <= input(44);
output(3, 190) <= input(47);
output(3, 191) <= input(49);
output(3, 192) <= input(10);
output(3, 193) <= input(11);
output(3, 194) <= input(12);
output(3, 195) <= input(13);
output(3, 196) <= input(14);
output(3, 197) <= input(15);
output(3, 198) <= input(32);
output(3, 199) <= input(34);
output(3, 200) <= input(36);
output(3, 201) <= input(37);
output(3, 202) <= input(40);
output(3, 203) <= input(42);
output(3, 204) <= input(44);
output(3, 205) <= input(47);
output(3, 206) <= input(49);
output(3, 207) <= input(50);
output(3, 208) <= input(26);
output(3, 209) <= input(27);
output(3, 210) <= input(28);
output(3, 211) <= input(29);
output(3, 212) <= input(30);
output(3, 213) <= input(31);
output(3, 214) <= input(33);
output(3, 215) <= input(35);
output(3, 216) <= input(38);
output(3, 217) <= input(39);
output(3, 218) <= input(41);
output(3, 219) <= input(43);
output(3, 220) <= input(45);
output(3, 221) <= input(46);
output(3, 222) <= input(48);
output(3, 223) <= input(52);
output(3, 224) <= input(27);
output(3, 225) <= input(28);
output(3, 226) <= input(29);
output(3, 227) <= input(30);
output(3, 228) <= input(31);
output(3, 229) <= input(33);
output(3, 230) <= input(35);
output(3, 231) <= input(38);
output(3, 232) <= input(39);
output(3, 233) <= input(41);
output(3, 234) <= input(43);
output(3, 235) <= input(45);
output(3, 236) <= input(46);
output(3, 237) <= input(48);
output(3, 238) <= input(52);
output(3, 239) <= input(53);
output(3, 240) <= input(28);
output(3, 241) <= input(29);
output(3, 242) <= input(30);
output(3, 243) <= input(31);
output(3, 244) <= input(33);
output(3, 245) <= input(35);
output(3, 246) <= input(38);
output(3, 247) <= input(39);
output(3, 248) <= input(41);
output(3, 249) <= input(43);
output(3, 250) <= input(45);
output(3, 251) <= input(46);
output(3, 252) <= input(48);
output(3, 253) <= input(52);
output(3, 254) <= input(53);
output(3, 255) <= input(54);
output(4, 0) <= input(0);
output(4, 1) <= input(1);
output(4, 2) <= input(2);
output(4, 3) <= input(3);
output(4, 4) <= input(4);
output(4, 5) <= input(5);
output(4, 6) <= input(6);
output(4, 7) <= input(7);
output(4, 8) <= input(8);
output(4, 9) <= input(9);
output(4, 10) <= input(10);
output(4, 11) <= input(11);
output(4, 12) <= input(12);
output(4, 13) <= input(13);
output(4, 14) <= input(14);
output(4, 15) <= input(15);
output(4, 16) <= input(1);
output(4, 17) <= input(2);
output(4, 18) <= input(3);
output(4, 19) <= input(4);
output(4, 20) <= input(5);
output(4, 21) <= input(6);
output(4, 22) <= input(7);
output(4, 23) <= input(8);
output(4, 24) <= input(9);
output(4, 25) <= input(10);
output(4, 26) <= input(11);
output(4, 27) <= input(12);
output(4, 28) <= input(13);
output(4, 29) <= input(14);
output(4, 30) <= input(15);
output(4, 31) <= input(32);
output(4, 32) <= input(2);
output(4, 33) <= input(3);
output(4, 34) <= input(4);
output(4, 35) <= input(5);
output(4, 36) <= input(6);
output(4, 37) <= input(7);
output(4, 38) <= input(8);
output(4, 39) <= input(9);
output(4, 40) <= input(10);
output(4, 41) <= input(11);
output(4, 42) <= input(12);
output(4, 43) <= input(13);
output(4, 44) <= input(14);
output(4, 45) <= input(15);
output(4, 46) <= input(32);
output(4, 47) <= input(34);
output(4, 48) <= input(3);
output(4, 49) <= input(4);
output(4, 50) <= input(5);
output(4, 51) <= input(6);
output(4, 52) <= input(7);
output(4, 53) <= input(8);
output(4, 54) <= input(9);
output(4, 55) <= input(10);
output(4, 56) <= input(11);
output(4, 57) <= input(12);
output(4, 58) <= input(13);
output(4, 59) <= input(14);
output(4, 60) <= input(15);
output(4, 61) <= input(32);
output(4, 62) <= input(34);
output(4, 63) <= input(36);
output(4, 64) <= input(4);
output(4, 65) <= input(5);
output(4, 66) <= input(6);
output(4, 67) <= input(7);
output(4, 68) <= input(8);
output(4, 69) <= input(9);
output(4, 70) <= input(10);
output(4, 71) <= input(11);
output(4, 72) <= input(12);
output(4, 73) <= input(13);
output(4, 74) <= input(14);
output(4, 75) <= input(15);
output(4, 76) <= input(32);
output(4, 77) <= input(34);
output(4, 78) <= input(36);
output(4, 79) <= input(37);
output(4, 80) <= input(20);
output(4, 81) <= input(21);
output(4, 82) <= input(22);
output(4, 83) <= input(23);
output(4, 84) <= input(24);
output(4, 85) <= input(25);
output(4, 86) <= input(26);
output(4, 87) <= input(27);
output(4, 88) <= input(28);
output(4, 89) <= input(29);
output(4, 90) <= input(30);
output(4, 91) <= input(31);
output(4, 92) <= input(33);
output(4, 93) <= input(35);
output(4, 94) <= input(38);
output(4, 95) <= input(39);
output(4, 96) <= input(21);
output(4, 97) <= input(22);
output(4, 98) <= input(23);
output(4, 99) <= input(24);
output(4, 100) <= input(25);
output(4, 101) <= input(26);
output(4, 102) <= input(27);
output(4, 103) <= input(28);
output(4, 104) <= input(29);
output(4, 105) <= input(30);
output(4, 106) <= input(31);
output(4, 107) <= input(33);
output(4, 108) <= input(35);
output(4, 109) <= input(38);
output(4, 110) <= input(39);
output(4, 111) <= input(41);
output(4, 112) <= input(22);
output(4, 113) <= input(23);
output(4, 114) <= input(24);
output(4, 115) <= input(25);
output(4, 116) <= input(26);
output(4, 117) <= input(27);
output(4, 118) <= input(28);
output(4, 119) <= input(29);
output(4, 120) <= input(30);
output(4, 121) <= input(31);
output(4, 122) <= input(33);
output(4, 123) <= input(35);
output(4, 124) <= input(38);
output(4, 125) <= input(39);
output(4, 126) <= input(41);
output(4, 127) <= input(43);
output(4, 128) <= input(23);
output(4, 129) <= input(24);
output(4, 130) <= input(25);
output(4, 131) <= input(26);
output(4, 132) <= input(27);
output(4, 133) <= input(28);
output(4, 134) <= input(29);
output(4, 135) <= input(30);
output(4, 136) <= input(31);
output(4, 137) <= input(33);
output(4, 138) <= input(35);
output(4, 139) <= input(38);
output(4, 140) <= input(39);
output(4, 141) <= input(41);
output(4, 142) <= input(43);
output(4, 143) <= input(45);
output(4, 144) <= input(24);
output(4, 145) <= input(25);
output(4, 146) <= input(26);
output(4, 147) <= input(27);
output(4, 148) <= input(28);
output(4, 149) <= input(29);
output(4, 150) <= input(30);
output(4, 151) <= input(31);
output(4, 152) <= input(33);
output(4, 153) <= input(35);
output(4, 154) <= input(38);
output(4, 155) <= input(39);
output(4, 156) <= input(41);
output(4, 157) <= input(43);
output(4, 158) <= input(45);
output(4, 159) <= input(46);
output(4, 160) <= input(9);
output(4, 161) <= input(10);
output(4, 162) <= input(11);
output(4, 163) <= input(12);
output(4, 164) <= input(13);
output(4, 165) <= input(14);
output(4, 166) <= input(15);
output(4, 167) <= input(32);
output(4, 168) <= input(34);
output(4, 169) <= input(36);
output(4, 170) <= input(37);
output(4, 171) <= input(40);
output(4, 172) <= input(42);
output(4, 173) <= input(44);
output(4, 174) <= input(47);
output(4, 175) <= input(49);
output(4, 176) <= input(10);
output(4, 177) <= input(11);
output(4, 178) <= input(12);
output(4, 179) <= input(13);
output(4, 180) <= input(14);
output(4, 181) <= input(15);
output(4, 182) <= input(32);
output(4, 183) <= input(34);
output(4, 184) <= input(36);
output(4, 185) <= input(37);
output(4, 186) <= input(40);
output(4, 187) <= input(42);
output(4, 188) <= input(44);
output(4, 189) <= input(47);
output(4, 190) <= input(49);
output(4, 191) <= input(50);
output(4, 192) <= input(11);
output(4, 193) <= input(12);
output(4, 194) <= input(13);
output(4, 195) <= input(14);
output(4, 196) <= input(15);
output(4, 197) <= input(32);
output(4, 198) <= input(34);
output(4, 199) <= input(36);
output(4, 200) <= input(37);
output(4, 201) <= input(40);
output(4, 202) <= input(42);
output(4, 203) <= input(44);
output(4, 204) <= input(47);
output(4, 205) <= input(49);
output(4, 206) <= input(50);
output(4, 207) <= input(51);
output(4, 208) <= input(12);
output(4, 209) <= input(13);
output(4, 210) <= input(14);
output(4, 211) <= input(15);
output(4, 212) <= input(32);
output(4, 213) <= input(34);
output(4, 214) <= input(36);
output(4, 215) <= input(37);
output(4, 216) <= input(40);
output(4, 217) <= input(42);
output(4, 218) <= input(44);
output(4, 219) <= input(47);
output(4, 220) <= input(49);
output(4, 221) <= input(50);
output(4, 222) <= input(51);
output(4, 223) <= input(55);
output(4, 224) <= input(13);
output(4, 225) <= input(14);
output(4, 226) <= input(15);
output(4, 227) <= input(32);
output(4, 228) <= input(34);
output(4, 229) <= input(36);
output(4, 230) <= input(37);
output(4, 231) <= input(40);
output(4, 232) <= input(42);
output(4, 233) <= input(44);
output(4, 234) <= input(47);
output(4, 235) <= input(49);
output(4, 236) <= input(50);
output(4, 237) <= input(51);
output(4, 238) <= input(55);
output(4, 239) <= input(56);
output(4, 240) <= input(14);
output(4, 241) <= input(15);
output(4, 242) <= input(32);
output(4, 243) <= input(34);
output(4, 244) <= input(36);
output(4, 245) <= input(37);
output(4, 246) <= input(40);
output(4, 247) <= input(42);
output(4, 248) <= input(44);
output(4, 249) <= input(47);
output(4, 250) <= input(49);
output(4, 251) <= input(50);
output(4, 252) <= input(51);
output(4, 253) <= input(55);
output(4, 254) <= input(56);
output(4, 255) <= input(57);
output(5, 0) <= input(16);
output(5, 1) <= input(17);
output(5, 2) <= input(18);
output(5, 3) <= input(19);
output(5, 4) <= input(20);
output(5, 5) <= input(21);
output(5, 6) <= input(22);
output(5, 7) <= input(23);
output(5, 8) <= input(24);
output(5, 9) <= input(25);
output(5, 10) <= input(26);
output(5, 11) <= input(27);
output(5, 12) <= input(28);
output(5, 13) <= input(29);
output(5, 14) <= input(30);
output(5, 15) <= input(31);
output(5, 16) <= input(17);
output(5, 17) <= input(18);
output(5, 18) <= input(19);
output(5, 19) <= input(20);
output(5, 20) <= input(21);
output(5, 21) <= input(22);
output(5, 22) <= input(23);
output(5, 23) <= input(24);
output(5, 24) <= input(25);
output(5, 25) <= input(26);
output(5, 26) <= input(27);
output(5, 27) <= input(28);
output(5, 28) <= input(29);
output(5, 29) <= input(30);
output(5, 30) <= input(31);
output(5, 31) <= input(33);
output(5, 32) <= input(18);
output(5, 33) <= input(19);
output(5, 34) <= input(20);
output(5, 35) <= input(21);
output(5, 36) <= input(22);
output(5, 37) <= input(23);
output(5, 38) <= input(24);
output(5, 39) <= input(25);
output(5, 40) <= input(26);
output(5, 41) <= input(27);
output(5, 42) <= input(28);
output(5, 43) <= input(29);
output(5, 44) <= input(30);
output(5, 45) <= input(31);
output(5, 46) <= input(33);
output(5, 47) <= input(35);
output(5, 48) <= input(19);
output(5, 49) <= input(20);
output(5, 50) <= input(21);
output(5, 51) <= input(22);
output(5, 52) <= input(23);
output(5, 53) <= input(24);
output(5, 54) <= input(25);
output(5, 55) <= input(26);
output(5, 56) <= input(27);
output(5, 57) <= input(28);
output(5, 58) <= input(29);
output(5, 59) <= input(30);
output(5, 60) <= input(31);
output(5, 61) <= input(33);
output(5, 62) <= input(35);
output(5, 63) <= input(38);
output(5, 64) <= input(20);
output(5, 65) <= input(21);
output(5, 66) <= input(22);
output(5, 67) <= input(23);
output(5, 68) <= input(24);
output(5, 69) <= input(25);
output(5, 70) <= input(26);
output(5, 71) <= input(27);
output(5, 72) <= input(28);
output(5, 73) <= input(29);
output(5, 74) <= input(30);
output(5, 75) <= input(31);
output(5, 76) <= input(33);
output(5, 77) <= input(35);
output(5, 78) <= input(38);
output(5, 79) <= input(39);
output(5, 80) <= input(21);
output(5, 81) <= input(22);
output(5, 82) <= input(23);
output(5, 83) <= input(24);
output(5, 84) <= input(25);
output(5, 85) <= input(26);
output(5, 86) <= input(27);
output(5, 87) <= input(28);
output(5, 88) <= input(29);
output(5, 89) <= input(30);
output(5, 90) <= input(31);
output(5, 91) <= input(33);
output(5, 92) <= input(35);
output(5, 93) <= input(38);
output(5, 94) <= input(39);
output(5, 95) <= input(41);
output(5, 96) <= input(22);
output(5, 97) <= input(23);
output(5, 98) <= input(24);
output(5, 99) <= input(25);
output(5, 100) <= input(26);
output(5, 101) <= input(27);
output(5, 102) <= input(28);
output(5, 103) <= input(29);
output(5, 104) <= input(30);
output(5, 105) <= input(31);
output(5, 106) <= input(33);
output(5, 107) <= input(35);
output(5, 108) <= input(38);
output(5, 109) <= input(39);
output(5, 110) <= input(41);
output(5, 111) <= input(43);
output(5, 112) <= input(23);
output(5, 113) <= input(24);
output(5, 114) <= input(25);
output(5, 115) <= input(26);
output(5, 116) <= input(27);
output(5, 117) <= input(28);
output(5, 118) <= input(29);
output(5, 119) <= input(30);
output(5, 120) <= input(31);
output(5, 121) <= input(33);
output(5, 122) <= input(35);
output(5, 123) <= input(38);
output(5, 124) <= input(39);
output(5, 125) <= input(41);
output(5, 126) <= input(43);
output(5, 127) <= input(45);
output(5, 128) <= input(24);
output(5, 129) <= input(25);
output(5, 130) <= input(26);
output(5, 131) <= input(27);
output(5, 132) <= input(28);
output(5, 133) <= input(29);
output(5, 134) <= input(30);
output(5, 135) <= input(31);
output(5, 136) <= input(33);
output(5, 137) <= input(35);
output(5, 138) <= input(38);
output(5, 139) <= input(39);
output(5, 140) <= input(41);
output(5, 141) <= input(43);
output(5, 142) <= input(45);
output(5, 143) <= input(46);
output(5, 144) <= input(25);
output(5, 145) <= input(26);
output(5, 146) <= input(27);
output(5, 147) <= input(28);
output(5, 148) <= input(29);
output(5, 149) <= input(30);
output(5, 150) <= input(31);
output(5, 151) <= input(33);
output(5, 152) <= input(35);
output(5, 153) <= input(38);
output(5, 154) <= input(39);
output(5, 155) <= input(41);
output(5, 156) <= input(43);
output(5, 157) <= input(45);
output(5, 158) <= input(46);
output(5, 159) <= input(48);
output(5, 160) <= input(26);
output(5, 161) <= input(27);
output(5, 162) <= input(28);
output(5, 163) <= input(29);
output(5, 164) <= input(30);
output(5, 165) <= input(31);
output(5, 166) <= input(33);
output(5, 167) <= input(35);
output(5, 168) <= input(38);
output(5, 169) <= input(39);
output(5, 170) <= input(41);
output(5, 171) <= input(43);
output(5, 172) <= input(45);
output(5, 173) <= input(46);
output(5, 174) <= input(48);
output(5, 175) <= input(52);
output(5, 176) <= input(27);
output(5, 177) <= input(28);
output(5, 178) <= input(29);
output(5, 179) <= input(30);
output(5, 180) <= input(31);
output(5, 181) <= input(33);
output(5, 182) <= input(35);
output(5, 183) <= input(38);
output(5, 184) <= input(39);
output(5, 185) <= input(41);
output(5, 186) <= input(43);
output(5, 187) <= input(45);
output(5, 188) <= input(46);
output(5, 189) <= input(48);
output(5, 190) <= input(52);
output(5, 191) <= input(53);
output(5, 192) <= input(28);
output(5, 193) <= input(29);
output(5, 194) <= input(30);
output(5, 195) <= input(31);
output(5, 196) <= input(33);
output(5, 197) <= input(35);
output(5, 198) <= input(38);
output(5, 199) <= input(39);
output(5, 200) <= input(41);
output(5, 201) <= input(43);
output(5, 202) <= input(45);
output(5, 203) <= input(46);
output(5, 204) <= input(48);
output(5, 205) <= input(52);
output(5, 206) <= input(53);
output(5, 207) <= input(54);
output(5, 208) <= input(29);
output(5, 209) <= input(30);
output(5, 210) <= input(31);
output(5, 211) <= input(33);
output(5, 212) <= input(35);
output(5, 213) <= input(38);
output(5, 214) <= input(39);
output(5, 215) <= input(41);
output(5, 216) <= input(43);
output(5, 217) <= input(45);
output(5, 218) <= input(46);
output(5, 219) <= input(48);
output(5, 220) <= input(52);
output(5, 221) <= input(53);
output(5, 222) <= input(54);
output(5, 223) <= input(58);
output(5, 224) <= input(30);
output(5, 225) <= input(31);
output(5, 226) <= input(33);
output(5, 227) <= input(35);
output(5, 228) <= input(38);
output(5, 229) <= input(39);
output(5, 230) <= input(41);
output(5, 231) <= input(43);
output(5, 232) <= input(45);
output(5, 233) <= input(46);
output(5, 234) <= input(48);
output(5, 235) <= input(52);
output(5, 236) <= input(53);
output(5, 237) <= input(54);
output(5, 238) <= input(58);
output(5, 239) <= input(59);
output(5, 240) <= input(31);
output(5, 241) <= input(33);
output(5, 242) <= input(35);
output(5, 243) <= input(38);
output(5, 244) <= input(39);
output(5, 245) <= input(41);
output(5, 246) <= input(43);
output(5, 247) <= input(45);
output(5, 248) <= input(46);
output(5, 249) <= input(48);
output(5, 250) <= input(52);
output(5, 251) <= input(53);
output(5, 252) <= input(54);
output(5, 253) <= input(58);
output(5, 254) <= input(59);
output(5, 255) <= input(60);
when others => for i in 0 to 7 loop for j in 0 to 255 loop output(i,j) <= "00000000"; end loop; end loop;
end case;
elsif control = "100" then 
case iteration_control is
when "0000" =>
output(0, 0) <= input(0);
output(0, 1) <= input(1);
output(0, 2) <= input(2);
output(0, 3) <= input(3);
output(0, 4) <= input(4);
output(0, 5) <= input(5);
output(0, 6) <= input(6);
output(0, 7) <= input(7);
output(0, 8) <= input(8);
output(0, 9) <= input(9);
output(0, 10) <= input(10);
output(0, 11) <= input(11);
output(0, 12) <= input(12);
output(0, 13) <= input(13);
output(0, 14) <= input(14);
output(0, 15) <= input(15);
output(0, 16) <= input(1);
output(0, 17) <= input(2);
output(0, 18) <= input(3);
output(0, 19) <= input(4);
output(0, 20) <= input(5);
output(0, 21) <= input(6);
output(0, 22) <= input(7);
output(0, 23) <= input(8);
output(0, 24) <= input(9);
output(0, 25) <= input(10);
output(0, 26) <= input(11);
output(0, 27) <= input(12);
output(0, 28) <= input(13);
output(0, 29) <= input(14);
output(0, 30) <= input(15);
output(0, 31) <= input(16);
output(0, 32) <= input(2);
output(0, 33) <= input(3);
output(0, 34) <= input(4);
output(0, 35) <= input(5);
output(0, 36) <= input(6);
output(0, 37) <= input(7);
output(0, 38) <= input(8);
output(0, 39) <= input(9);
output(0, 40) <= input(10);
output(0, 41) <= input(11);
output(0, 42) <= input(12);
output(0, 43) <= input(13);
output(0, 44) <= input(14);
output(0, 45) <= input(15);
output(0, 46) <= input(16);
output(0, 47) <= input(17);
output(0, 48) <= input(3);
output(0, 49) <= input(4);
output(0, 50) <= input(5);
output(0, 51) <= input(6);
output(0, 52) <= input(7);
output(0, 53) <= input(8);
output(0, 54) <= input(9);
output(0, 55) <= input(10);
output(0, 56) <= input(11);
output(0, 57) <= input(12);
output(0, 58) <= input(13);
output(0, 59) <= input(14);
output(0, 60) <= input(15);
output(0, 61) <= input(16);
output(0, 62) <= input(17);
output(0, 63) <= input(18);
output(0, 64) <= input(4);
output(0, 65) <= input(5);
output(0, 66) <= input(6);
output(0, 67) <= input(7);
output(0, 68) <= input(8);
output(0, 69) <= input(9);
output(0, 70) <= input(10);
output(0, 71) <= input(11);
output(0, 72) <= input(12);
output(0, 73) <= input(13);
output(0, 74) <= input(14);
output(0, 75) <= input(15);
output(0, 76) <= input(16);
output(0, 77) <= input(17);
output(0, 78) <= input(18);
output(0, 79) <= input(19);
output(0, 80) <= input(5);
output(0, 81) <= input(6);
output(0, 82) <= input(7);
output(0, 83) <= input(8);
output(0, 84) <= input(9);
output(0, 85) <= input(10);
output(0, 86) <= input(11);
output(0, 87) <= input(12);
output(0, 88) <= input(13);
output(0, 89) <= input(14);
output(0, 90) <= input(15);
output(0, 91) <= input(16);
output(0, 92) <= input(17);
output(0, 93) <= input(18);
output(0, 94) <= input(19);
output(0, 95) <= input(20);
output(0, 96) <= input(6);
output(0, 97) <= input(7);
output(0, 98) <= input(8);
output(0, 99) <= input(9);
output(0, 100) <= input(10);
output(0, 101) <= input(11);
output(0, 102) <= input(12);
output(0, 103) <= input(13);
output(0, 104) <= input(14);
output(0, 105) <= input(15);
output(0, 106) <= input(16);
output(0, 107) <= input(17);
output(0, 108) <= input(18);
output(0, 109) <= input(19);
output(0, 110) <= input(20);
output(0, 111) <= input(21);
output(0, 112) <= input(7);
output(0, 113) <= input(8);
output(0, 114) <= input(9);
output(0, 115) <= input(10);
output(0, 116) <= input(11);
output(0, 117) <= input(12);
output(0, 118) <= input(13);
output(0, 119) <= input(14);
output(0, 120) <= input(15);
output(0, 121) <= input(16);
output(0, 122) <= input(17);
output(0, 123) <= input(18);
output(0, 124) <= input(19);
output(0, 125) <= input(20);
output(0, 126) <= input(21);
output(0, 127) <= input(22);
output(0, 128) <= input(8);
output(0, 129) <= input(9);
output(0, 130) <= input(10);
output(0, 131) <= input(11);
output(0, 132) <= input(12);
output(0, 133) <= input(13);
output(0, 134) <= input(14);
output(0, 135) <= input(15);
output(0, 136) <= input(16);
output(0, 137) <= input(17);
output(0, 138) <= input(18);
output(0, 139) <= input(19);
output(0, 140) <= input(20);
output(0, 141) <= input(21);
output(0, 142) <= input(22);
output(0, 143) <= input(23);
output(0, 144) <= input(9);
output(0, 145) <= input(10);
output(0, 146) <= input(11);
output(0, 147) <= input(12);
output(0, 148) <= input(13);
output(0, 149) <= input(14);
output(0, 150) <= input(15);
output(0, 151) <= input(16);
output(0, 152) <= input(17);
output(0, 153) <= input(18);
output(0, 154) <= input(19);
output(0, 155) <= input(20);
output(0, 156) <= input(21);
output(0, 157) <= input(22);
output(0, 158) <= input(23);
output(0, 159) <= input(24);
output(0, 160) <= input(10);
output(0, 161) <= input(11);
output(0, 162) <= input(12);
output(0, 163) <= input(13);
output(0, 164) <= input(14);
output(0, 165) <= input(15);
output(0, 166) <= input(16);
output(0, 167) <= input(17);
output(0, 168) <= input(18);
output(0, 169) <= input(19);
output(0, 170) <= input(20);
output(0, 171) <= input(21);
output(0, 172) <= input(22);
output(0, 173) <= input(23);
output(0, 174) <= input(24);
output(0, 175) <= input(25);
output(0, 176) <= input(11);
output(0, 177) <= input(12);
output(0, 178) <= input(13);
output(0, 179) <= input(14);
output(0, 180) <= input(15);
output(0, 181) <= input(16);
output(0, 182) <= input(17);
output(0, 183) <= input(18);
output(0, 184) <= input(19);
output(0, 185) <= input(20);
output(0, 186) <= input(21);
output(0, 187) <= input(22);
output(0, 188) <= input(23);
output(0, 189) <= input(24);
output(0, 190) <= input(25);
output(0, 191) <= input(26);
output(0, 192) <= input(12);
output(0, 193) <= input(13);
output(0, 194) <= input(14);
output(0, 195) <= input(15);
output(0, 196) <= input(16);
output(0, 197) <= input(17);
output(0, 198) <= input(18);
output(0, 199) <= input(19);
output(0, 200) <= input(20);
output(0, 201) <= input(21);
output(0, 202) <= input(22);
output(0, 203) <= input(23);
output(0, 204) <= input(24);
output(0, 205) <= input(25);
output(0, 206) <= input(26);
output(0, 207) <= input(27);
output(0, 208) <= input(13);
output(0, 209) <= input(14);
output(0, 210) <= input(15);
output(0, 211) <= input(16);
output(0, 212) <= input(17);
output(0, 213) <= input(18);
output(0, 214) <= input(19);
output(0, 215) <= input(20);
output(0, 216) <= input(21);
output(0, 217) <= input(22);
output(0, 218) <= input(23);
output(0, 219) <= input(24);
output(0, 220) <= input(25);
output(0, 221) <= input(26);
output(0, 222) <= input(27);
output(0, 223) <= input(28);
output(0, 224) <= input(14);
output(0, 225) <= input(15);
output(0, 226) <= input(16);
output(0, 227) <= input(17);
output(0, 228) <= input(18);
output(0, 229) <= input(19);
output(0, 230) <= input(20);
output(0, 231) <= input(21);
output(0, 232) <= input(22);
output(0, 233) <= input(23);
output(0, 234) <= input(24);
output(0, 235) <= input(25);
output(0, 236) <= input(26);
output(0, 237) <= input(27);
output(0, 238) <= input(28);
output(0, 239) <= input(29);
output(0, 240) <= input(15);
output(0, 241) <= input(16);
output(0, 242) <= input(17);
output(0, 243) <= input(18);
output(0, 244) <= input(19);
output(0, 245) <= input(20);
output(0, 246) <= input(21);
output(0, 247) <= input(22);
output(0, 248) <= input(23);
output(0, 249) <= input(24);
output(0, 250) <= input(25);
output(0, 251) <= input(26);
output(0, 252) <= input(27);
output(0, 253) <= input(28);
output(0, 254) <= input(29);
output(0, 255) <= input(30);
output(1, 0) <= input(31);
output(1, 1) <= input(32);
output(1, 2) <= input(0);
output(1, 3) <= input(1);
output(1, 4) <= input(2);
output(1, 5) <= input(3);
output(1, 6) <= input(4);
output(1, 7) <= input(5);
output(1, 8) <= input(6);
output(1, 9) <= input(7);
output(1, 10) <= input(8);
output(1, 11) <= input(9);
output(1, 12) <= input(10);
output(1, 13) <= input(11);
output(1, 14) <= input(12);
output(1, 15) <= input(13);
output(1, 16) <= input(32);
output(1, 17) <= input(0);
output(1, 18) <= input(1);
output(1, 19) <= input(2);
output(1, 20) <= input(3);
output(1, 21) <= input(4);
output(1, 22) <= input(5);
output(1, 23) <= input(6);
output(1, 24) <= input(7);
output(1, 25) <= input(8);
output(1, 26) <= input(9);
output(1, 27) <= input(10);
output(1, 28) <= input(11);
output(1, 29) <= input(12);
output(1, 30) <= input(13);
output(1, 31) <= input(14);
output(1, 32) <= input(0);
output(1, 33) <= input(1);
output(1, 34) <= input(2);
output(1, 35) <= input(3);
output(1, 36) <= input(4);
output(1, 37) <= input(5);
output(1, 38) <= input(6);
output(1, 39) <= input(7);
output(1, 40) <= input(8);
output(1, 41) <= input(9);
output(1, 42) <= input(10);
output(1, 43) <= input(11);
output(1, 44) <= input(12);
output(1, 45) <= input(13);
output(1, 46) <= input(14);
output(1, 47) <= input(15);
output(1, 48) <= input(1);
output(1, 49) <= input(2);
output(1, 50) <= input(3);
output(1, 51) <= input(4);
output(1, 52) <= input(5);
output(1, 53) <= input(6);
output(1, 54) <= input(7);
output(1, 55) <= input(8);
output(1, 56) <= input(9);
output(1, 57) <= input(10);
output(1, 58) <= input(11);
output(1, 59) <= input(12);
output(1, 60) <= input(13);
output(1, 61) <= input(14);
output(1, 62) <= input(15);
output(1, 63) <= input(16);
output(1, 64) <= input(2);
output(1, 65) <= input(3);
output(1, 66) <= input(4);
output(1, 67) <= input(5);
output(1, 68) <= input(6);
output(1, 69) <= input(7);
output(1, 70) <= input(8);
output(1, 71) <= input(9);
output(1, 72) <= input(10);
output(1, 73) <= input(11);
output(1, 74) <= input(12);
output(1, 75) <= input(13);
output(1, 76) <= input(14);
output(1, 77) <= input(15);
output(1, 78) <= input(16);
output(1, 79) <= input(17);
output(1, 80) <= input(33);
output(1, 81) <= input(34);
output(1, 82) <= input(35);
output(1, 83) <= input(36);
output(1, 84) <= input(37);
output(1, 85) <= input(38);
output(1, 86) <= input(39);
output(1, 87) <= input(40);
output(1, 88) <= input(41);
output(1, 89) <= input(42);
output(1, 90) <= input(43);
output(1, 91) <= input(44);
output(1, 92) <= input(45);
output(1, 93) <= input(46);
output(1, 94) <= input(47);
output(1, 95) <= input(48);
output(1, 96) <= input(34);
output(1, 97) <= input(35);
output(1, 98) <= input(36);
output(1, 99) <= input(37);
output(1, 100) <= input(38);
output(1, 101) <= input(39);
output(1, 102) <= input(40);
output(1, 103) <= input(41);
output(1, 104) <= input(42);
output(1, 105) <= input(43);
output(1, 106) <= input(44);
output(1, 107) <= input(45);
output(1, 108) <= input(46);
output(1, 109) <= input(47);
output(1, 110) <= input(48);
output(1, 111) <= input(49);
output(1, 112) <= input(35);
output(1, 113) <= input(36);
output(1, 114) <= input(37);
output(1, 115) <= input(38);
output(1, 116) <= input(39);
output(1, 117) <= input(40);
output(1, 118) <= input(41);
output(1, 119) <= input(42);
output(1, 120) <= input(43);
output(1, 121) <= input(44);
output(1, 122) <= input(45);
output(1, 123) <= input(46);
output(1, 124) <= input(47);
output(1, 125) <= input(48);
output(1, 126) <= input(49);
output(1, 127) <= input(50);
output(1, 128) <= input(36);
output(1, 129) <= input(37);
output(1, 130) <= input(38);
output(1, 131) <= input(39);
output(1, 132) <= input(40);
output(1, 133) <= input(41);
output(1, 134) <= input(42);
output(1, 135) <= input(43);
output(1, 136) <= input(44);
output(1, 137) <= input(45);
output(1, 138) <= input(46);
output(1, 139) <= input(47);
output(1, 140) <= input(48);
output(1, 141) <= input(49);
output(1, 142) <= input(50);
output(1, 143) <= input(51);
output(1, 144) <= input(37);
output(1, 145) <= input(38);
output(1, 146) <= input(39);
output(1, 147) <= input(40);
output(1, 148) <= input(41);
output(1, 149) <= input(42);
output(1, 150) <= input(43);
output(1, 151) <= input(44);
output(1, 152) <= input(45);
output(1, 153) <= input(46);
output(1, 154) <= input(47);
output(1, 155) <= input(48);
output(1, 156) <= input(49);
output(1, 157) <= input(50);
output(1, 158) <= input(51);
output(1, 159) <= input(52);
output(1, 160) <= input(7);
output(1, 161) <= input(8);
output(1, 162) <= input(9);
output(1, 163) <= input(10);
output(1, 164) <= input(11);
output(1, 165) <= input(12);
output(1, 166) <= input(13);
output(1, 167) <= input(14);
output(1, 168) <= input(15);
output(1, 169) <= input(16);
output(1, 170) <= input(17);
output(1, 171) <= input(18);
output(1, 172) <= input(19);
output(1, 173) <= input(20);
output(1, 174) <= input(21);
output(1, 175) <= input(22);
output(1, 176) <= input(8);
output(1, 177) <= input(9);
output(1, 178) <= input(10);
output(1, 179) <= input(11);
output(1, 180) <= input(12);
output(1, 181) <= input(13);
output(1, 182) <= input(14);
output(1, 183) <= input(15);
output(1, 184) <= input(16);
output(1, 185) <= input(17);
output(1, 186) <= input(18);
output(1, 187) <= input(19);
output(1, 188) <= input(20);
output(1, 189) <= input(21);
output(1, 190) <= input(22);
output(1, 191) <= input(23);
output(1, 192) <= input(9);
output(1, 193) <= input(10);
output(1, 194) <= input(11);
output(1, 195) <= input(12);
output(1, 196) <= input(13);
output(1, 197) <= input(14);
output(1, 198) <= input(15);
output(1, 199) <= input(16);
output(1, 200) <= input(17);
output(1, 201) <= input(18);
output(1, 202) <= input(19);
output(1, 203) <= input(20);
output(1, 204) <= input(21);
output(1, 205) <= input(22);
output(1, 206) <= input(23);
output(1, 207) <= input(24);
output(1, 208) <= input(10);
output(1, 209) <= input(11);
output(1, 210) <= input(12);
output(1, 211) <= input(13);
output(1, 212) <= input(14);
output(1, 213) <= input(15);
output(1, 214) <= input(16);
output(1, 215) <= input(17);
output(1, 216) <= input(18);
output(1, 217) <= input(19);
output(1, 218) <= input(20);
output(1, 219) <= input(21);
output(1, 220) <= input(22);
output(1, 221) <= input(23);
output(1, 222) <= input(24);
output(1, 223) <= input(25);
output(1, 224) <= input(11);
output(1, 225) <= input(12);
output(1, 226) <= input(13);
output(1, 227) <= input(14);
output(1, 228) <= input(15);
output(1, 229) <= input(16);
output(1, 230) <= input(17);
output(1, 231) <= input(18);
output(1, 232) <= input(19);
output(1, 233) <= input(20);
output(1, 234) <= input(21);
output(1, 235) <= input(22);
output(1, 236) <= input(23);
output(1, 237) <= input(24);
output(1, 238) <= input(25);
output(1, 239) <= input(26);
output(1, 240) <= input(12);
output(1, 241) <= input(13);
output(1, 242) <= input(14);
output(1, 243) <= input(15);
output(1, 244) <= input(16);
output(1, 245) <= input(17);
output(1, 246) <= input(18);
output(1, 247) <= input(19);
output(1, 248) <= input(20);
output(1, 249) <= input(21);
output(1, 250) <= input(22);
output(1, 251) <= input(23);
output(1, 252) <= input(24);
output(1, 253) <= input(25);
output(1, 254) <= input(26);
output(1, 255) <= input(27);
output(2, 0) <= input(53);
output(2, 1) <= input(54);
output(2, 2) <= input(55);
output(2, 3) <= input(56);
output(2, 4) <= input(57);
output(2, 5) <= input(58);
output(2, 6) <= input(33);
output(2, 7) <= input(34);
output(2, 8) <= input(35);
output(2, 9) <= input(36);
output(2, 10) <= input(37);
output(2, 11) <= input(38);
output(2, 12) <= input(39);
output(2, 13) <= input(40);
output(2, 14) <= input(41);
output(2, 15) <= input(42);
output(2, 16) <= input(54);
output(2, 17) <= input(55);
output(2, 18) <= input(56);
output(2, 19) <= input(57);
output(2, 20) <= input(58);
output(2, 21) <= input(33);
output(2, 22) <= input(34);
output(2, 23) <= input(35);
output(2, 24) <= input(36);
output(2, 25) <= input(37);
output(2, 26) <= input(38);
output(2, 27) <= input(39);
output(2, 28) <= input(40);
output(2, 29) <= input(41);
output(2, 30) <= input(42);
output(2, 31) <= input(43);
output(2, 32) <= input(31);
output(2, 33) <= input(32);
output(2, 34) <= input(0);
output(2, 35) <= input(1);
output(2, 36) <= input(2);
output(2, 37) <= input(3);
output(2, 38) <= input(4);
output(2, 39) <= input(5);
output(2, 40) <= input(6);
output(2, 41) <= input(7);
output(2, 42) <= input(8);
output(2, 43) <= input(9);
output(2, 44) <= input(10);
output(2, 45) <= input(11);
output(2, 46) <= input(12);
output(2, 47) <= input(13);
output(2, 48) <= input(32);
output(2, 49) <= input(0);
output(2, 50) <= input(1);
output(2, 51) <= input(2);
output(2, 52) <= input(3);
output(2, 53) <= input(4);
output(2, 54) <= input(5);
output(2, 55) <= input(6);
output(2, 56) <= input(7);
output(2, 57) <= input(8);
output(2, 58) <= input(9);
output(2, 59) <= input(10);
output(2, 60) <= input(11);
output(2, 61) <= input(12);
output(2, 62) <= input(13);
output(2, 63) <= input(14);
output(2, 64) <= input(0);
output(2, 65) <= input(1);
output(2, 66) <= input(2);
output(2, 67) <= input(3);
output(2, 68) <= input(4);
output(2, 69) <= input(5);
output(2, 70) <= input(6);
output(2, 71) <= input(7);
output(2, 72) <= input(8);
output(2, 73) <= input(9);
output(2, 74) <= input(10);
output(2, 75) <= input(11);
output(2, 76) <= input(12);
output(2, 77) <= input(13);
output(2, 78) <= input(14);
output(2, 79) <= input(15);
output(2, 80) <= input(57);
output(2, 81) <= input(58);
output(2, 82) <= input(33);
output(2, 83) <= input(34);
output(2, 84) <= input(35);
output(2, 85) <= input(36);
output(2, 86) <= input(37);
output(2, 87) <= input(38);
output(2, 88) <= input(39);
output(2, 89) <= input(40);
output(2, 90) <= input(41);
output(2, 91) <= input(42);
output(2, 92) <= input(43);
output(2, 93) <= input(44);
output(2, 94) <= input(45);
output(2, 95) <= input(46);
output(2, 96) <= input(58);
output(2, 97) <= input(33);
output(2, 98) <= input(34);
output(2, 99) <= input(35);
output(2, 100) <= input(36);
output(2, 101) <= input(37);
output(2, 102) <= input(38);
output(2, 103) <= input(39);
output(2, 104) <= input(40);
output(2, 105) <= input(41);
output(2, 106) <= input(42);
output(2, 107) <= input(43);
output(2, 108) <= input(44);
output(2, 109) <= input(45);
output(2, 110) <= input(46);
output(2, 111) <= input(47);
output(2, 112) <= input(33);
output(2, 113) <= input(34);
output(2, 114) <= input(35);
output(2, 115) <= input(36);
output(2, 116) <= input(37);
output(2, 117) <= input(38);
output(2, 118) <= input(39);
output(2, 119) <= input(40);
output(2, 120) <= input(41);
output(2, 121) <= input(42);
output(2, 122) <= input(43);
output(2, 123) <= input(44);
output(2, 124) <= input(45);
output(2, 125) <= input(46);
output(2, 126) <= input(47);
output(2, 127) <= input(48);
output(2, 128) <= input(3);
output(2, 129) <= input(4);
output(2, 130) <= input(5);
output(2, 131) <= input(6);
output(2, 132) <= input(7);
output(2, 133) <= input(8);
output(2, 134) <= input(9);
output(2, 135) <= input(10);
output(2, 136) <= input(11);
output(2, 137) <= input(12);
output(2, 138) <= input(13);
output(2, 139) <= input(14);
output(2, 140) <= input(15);
output(2, 141) <= input(16);
output(2, 142) <= input(17);
output(2, 143) <= input(18);
output(2, 144) <= input(4);
output(2, 145) <= input(5);
output(2, 146) <= input(6);
output(2, 147) <= input(7);
output(2, 148) <= input(8);
output(2, 149) <= input(9);
output(2, 150) <= input(10);
output(2, 151) <= input(11);
output(2, 152) <= input(12);
output(2, 153) <= input(13);
output(2, 154) <= input(14);
output(2, 155) <= input(15);
output(2, 156) <= input(16);
output(2, 157) <= input(17);
output(2, 158) <= input(18);
output(2, 159) <= input(19);
output(2, 160) <= input(35);
output(2, 161) <= input(36);
output(2, 162) <= input(37);
output(2, 163) <= input(38);
output(2, 164) <= input(39);
output(2, 165) <= input(40);
output(2, 166) <= input(41);
output(2, 167) <= input(42);
output(2, 168) <= input(43);
output(2, 169) <= input(44);
output(2, 170) <= input(45);
output(2, 171) <= input(46);
output(2, 172) <= input(47);
output(2, 173) <= input(48);
output(2, 174) <= input(49);
output(2, 175) <= input(50);
output(2, 176) <= input(36);
output(2, 177) <= input(37);
output(2, 178) <= input(38);
output(2, 179) <= input(39);
output(2, 180) <= input(40);
output(2, 181) <= input(41);
output(2, 182) <= input(42);
output(2, 183) <= input(43);
output(2, 184) <= input(44);
output(2, 185) <= input(45);
output(2, 186) <= input(46);
output(2, 187) <= input(47);
output(2, 188) <= input(48);
output(2, 189) <= input(49);
output(2, 190) <= input(50);
output(2, 191) <= input(51);
output(2, 192) <= input(37);
output(2, 193) <= input(38);
output(2, 194) <= input(39);
output(2, 195) <= input(40);
output(2, 196) <= input(41);
output(2, 197) <= input(42);
output(2, 198) <= input(43);
output(2, 199) <= input(44);
output(2, 200) <= input(45);
output(2, 201) <= input(46);
output(2, 202) <= input(47);
output(2, 203) <= input(48);
output(2, 204) <= input(49);
output(2, 205) <= input(50);
output(2, 206) <= input(51);
output(2, 207) <= input(52);
output(2, 208) <= input(7);
output(2, 209) <= input(8);
output(2, 210) <= input(9);
output(2, 211) <= input(10);
output(2, 212) <= input(11);
output(2, 213) <= input(12);
output(2, 214) <= input(13);
output(2, 215) <= input(14);
output(2, 216) <= input(15);
output(2, 217) <= input(16);
output(2, 218) <= input(17);
output(2, 219) <= input(18);
output(2, 220) <= input(19);
output(2, 221) <= input(20);
output(2, 222) <= input(21);
output(2, 223) <= input(22);
output(2, 224) <= input(8);
output(2, 225) <= input(9);
output(2, 226) <= input(10);
output(2, 227) <= input(11);
output(2, 228) <= input(12);
output(2, 229) <= input(13);
output(2, 230) <= input(14);
output(2, 231) <= input(15);
output(2, 232) <= input(16);
output(2, 233) <= input(17);
output(2, 234) <= input(18);
output(2, 235) <= input(19);
output(2, 236) <= input(20);
output(2, 237) <= input(21);
output(2, 238) <= input(22);
output(2, 239) <= input(23);
output(2, 240) <= input(9);
output(2, 241) <= input(10);
output(2, 242) <= input(11);
output(2, 243) <= input(12);
output(2, 244) <= input(13);
output(2, 245) <= input(14);
output(2, 246) <= input(15);
output(2, 247) <= input(16);
output(2, 248) <= input(17);
output(2, 249) <= input(18);
output(2, 250) <= input(19);
output(2, 251) <= input(20);
output(2, 252) <= input(21);
output(2, 253) <= input(22);
output(2, 254) <= input(23);
output(2, 255) <= input(24);
output(3, 0) <= input(59);
output(3, 1) <= input(60);
output(3, 2) <= input(61);
output(3, 3) <= input(31);
output(3, 4) <= input(32);
output(3, 5) <= input(0);
output(3, 6) <= input(1);
output(3, 7) <= input(2);
output(3, 8) <= input(3);
output(3, 9) <= input(4);
output(3, 10) <= input(5);
output(3, 11) <= input(6);
output(3, 12) <= input(7);
output(3, 13) <= input(8);
output(3, 14) <= input(9);
output(3, 15) <= input(10);
output(3, 16) <= input(62);
output(3, 17) <= input(53);
output(3, 18) <= input(54);
output(3, 19) <= input(55);
output(3, 20) <= input(56);
output(3, 21) <= input(57);
output(3, 22) <= input(58);
output(3, 23) <= input(33);
output(3, 24) <= input(34);
output(3, 25) <= input(35);
output(3, 26) <= input(36);
output(3, 27) <= input(37);
output(3, 28) <= input(38);
output(3, 29) <= input(39);
output(3, 30) <= input(40);
output(3, 31) <= input(41);
output(3, 32) <= input(53);
output(3, 33) <= input(54);
output(3, 34) <= input(55);
output(3, 35) <= input(56);
output(3, 36) <= input(57);
output(3, 37) <= input(58);
output(3, 38) <= input(33);
output(3, 39) <= input(34);
output(3, 40) <= input(35);
output(3, 41) <= input(36);
output(3, 42) <= input(37);
output(3, 43) <= input(38);
output(3, 44) <= input(39);
output(3, 45) <= input(40);
output(3, 46) <= input(41);
output(3, 47) <= input(42);
output(3, 48) <= input(61);
output(3, 49) <= input(31);
output(3, 50) <= input(32);
output(3, 51) <= input(0);
output(3, 52) <= input(1);
output(3, 53) <= input(2);
output(3, 54) <= input(3);
output(3, 55) <= input(4);
output(3, 56) <= input(5);
output(3, 57) <= input(6);
output(3, 58) <= input(7);
output(3, 59) <= input(8);
output(3, 60) <= input(9);
output(3, 61) <= input(10);
output(3, 62) <= input(11);
output(3, 63) <= input(12);
output(3, 64) <= input(31);
output(3, 65) <= input(32);
output(3, 66) <= input(0);
output(3, 67) <= input(1);
output(3, 68) <= input(2);
output(3, 69) <= input(3);
output(3, 70) <= input(4);
output(3, 71) <= input(5);
output(3, 72) <= input(6);
output(3, 73) <= input(7);
output(3, 74) <= input(8);
output(3, 75) <= input(9);
output(3, 76) <= input(10);
output(3, 77) <= input(11);
output(3, 78) <= input(12);
output(3, 79) <= input(13);
output(3, 80) <= input(55);
output(3, 81) <= input(56);
output(3, 82) <= input(57);
output(3, 83) <= input(58);
output(3, 84) <= input(33);
output(3, 85) <= input(34);
output(3, 86) <= input(35);
output(3, 87) <= input(36);
output(3, 88) <= input(37);
output(3, 89) <= input(38);
output(3, 90) <= input(39);
output(3, 91) <= input(40);
output(3, 92) <= input(41);
output(3, 93) <= input(42);
output(3, 94) <= input(43);
output(3, 95) <= input(44);
output(3, 96) <= input(56);
output(3, 97) <= input(57);
output(3, 98) <= input(58);
output(3, 99) <= input(33);
output(3, 100) <= input(34);
output(3, 101) <= input(35);
output(3, 102) <= input(36);
output(3, 103) <= input(37);
output(3, 104) <= input(38);
output(3, 105) <= input(39);
output(3, 106) <= input(40);
output(3, 107) <= input(41);
output(3, 108) <= input(42);
output(3, 109) <= input(43);
output(3, 110) <= input(44);
output(3, 111) <= input(45);
output(3, 112) <= input(0);
output(3, 113) <= input(1);
output(3, 114) <= input(2);
output(3, 115) <= input(3);
output(3, 116) <= input(4);
output(3, 117) <= input(5);
output(3, 118) <= input(6);
output(3, 119) <= input(7);
output(3, 120) <= input(8);
output(3, 121) <= input(9);
output(3, 122) <= input(10);
output(3, 123) <= input(11);
output(3, 124) <= input(12);
output(3, 125) <= input(13);
output(3, 126) <= input(14);
output(3, 127) <= input(15);
output(3, 128) <= input(57);
output(3, 129) <= input(58);
output(3, 130) <= input(33);
output(3, 131) <= input(34);
output(3, 132) <= input(35);
output(3, 133) <= input(36);
output(3, 134) <= input(37);
output(3, 135) <= input(38);
output(3, 136) <= input(39);
output(3, 137) <= input(40);
output(3, 138) <= input(41);
output(3, 139) <= input(42);
output(3, 140) <= input(43);
output(3, 141) <= input(44);
output(3, 142) <= input(45);
output(3, 143) <= input(46);
output(3, 144) <= input(58);
output(3, 145) <= input(33);
output(3, 146) <= input(34);
output(3, 147) <= input(35);
output(3, 148) <= input(36);
output(3, 149) <= input(37);
output(3, 150) <= input(38);
output(3, 151) <= input(39);
output(3, 152) <= input(40);
output(3, 153) <= input(41);
output(3, 154) <= input(42);
output(3, 155) <= input(43);
output(3, 156) <= input(44);
output(3, 157) <= input(45);
output(3, 158) <= input(46);
output(3, 159) <= input(47);
output(3, 160) <= input(2);
output(3, 161) <= input(3);
output(3, 162) <= input(4);
output(3, 163) <= input(5);
output(3, 164) <= input(6);
output(3, 165) <= input(7);
output(3, 166) <= input(8);
output(3, 167) <= input(9);
output(3, 168) <= input(10);
output(3, 169) <= input(11);
output(3, 170) <= input(12);
output(3, 171) <= input(13);
output(3, 172) <= input(14);
output(3, 173) <= input(15);
output(3, 174) <= input(16);
output(3, 175) <= input(17);
output(3, 176) <= input(3);
output(3, 177) <= input(4);
output(3, 178) <= input(5);
output(3, 179) <= input(6);
output(3, 180) <= input(7);
output(3, 181) <= input(8);
output(3, 182) <= input(9);
output(3, 183) <= input(10);
output(3, 184) <= input(11);
output(3, 185) <= input(12);
output(3, 186) <= input(13);
output(3, 187) <= input(14);
output(3, 188) <= input(15);
output(3, 189) <= input(16);
output(3, 190) <= input(17);
output(3, 191) <= input(18);
output(3, 192) <= input(34);
output(3, 193) <= input(35);
output(3, 194) <= input(36);
output(3, 195) <= input(37);
output(3, 196) <= input(38);
output(3, 197) <= input(39);
output(3, 198) <= input(40);
output(3, 199) <= input(41);
output(3, 200) <= input(42);
output(3, 201) <= input(43);
output(3, 202) <= input(44);
output(3, 203) <= input(45);
output(3, 204) <= input(46);
output(3, 205) <= input(47);
output(3, 206) <= input(48);
output(3, 207) <= input(49);
output(3, 208) <= input(35);
output(3, 209) <= input(36);
output(3, 210) <= input(37);
output(3, 211) <= input(38);
output(3, 212) <= input(39);
output(3, 213) <= input(40);
output(3, 214) <= input(41);
output(3, 215) <= input(42);
output(3, 216) <= input(43);
output(3, 217) <= input(44);
output(3, 218) <= input(45);
output(3, 219) <= input(46);
output(3, 220) <= input(47);
output(3, 221) <= input(48);
output(3, 222) <= input(49);
output(3, 223) <= input(50);
output(3, 224) <= input(5);
output(3, 225) <= input(6);
output(3, 226) <= input(7);
output(3, 227) <= input(8);
output(3, 228) <= input(9);
output(3, 229) <= input(10);
output(3, 230) <= input(11);
output(3, 231) <= input(12);
output(3, 232) <= input(13);
output(3, 233) <= input(14);
output(3, 234) <= input(15);
output(3, 235) <= input(16);
output(3, 236) <= input(17);
output(3, 237) <= input(18);
output(3, 238) <= input(19);
output(3, 239) <= input(20);
output(3, 240) <= input(6);
output(3, 241) <= input(7);
output(3, 242) <= input(8);
output(3, 243) <= input(9);
output(3, 244) <= input(10);
output(3, 245) <= input(11);
output(3, 246) <= input(12);
output(3, 247) <= input(13);
output(3, 248) <= input(14);
output(3, 249) <= input(15);
output(3, 250) <= input(16);
output(3, 251) <= input(17);
output(3, 252) <= input(18);
output(3, 253) <= input(19);
output(3, 254) <= input(20);
output(3, 255) <= input(21);
output(4, 0) <= input(63);
output(4, 1) <= input(64);
output(4, 2) <= input(62);
output(4, 3) <= input(53);
output(4, 4) <= input(54);
output(4, 5) <= input(55);
output(4, 6) <= input(56);
output(4, 7) <= input(57);
output(4, 8) <= input(58);
output(4, 9) <= input(33);
output(4, 10) <= input(34);
output(4, 11) <= input(35);
output(4, 12) <= input(36);
output(4, 13) <= input(37);
output(4, 14) <= input(38);
output(4, 15) <= input(39);
output(4, 16) <= input(65);
output(4, 17) <= input(59);
output(4, 18) <= input(60);
output(4, 19) <= input(61);
output(4, 20) <= input(31);
output(4, 21) <= input(32);
output(4, 22) <= input(0);
output(4, 23) <= input(1);
output(4, 24) <= input(2);
output(4, 25) <= input(3);
output(4, 26) <= input(4);
output(4, 27) <= input(5);
output(4, 28) <= input(6);
output(4, 29) <= input(7);
output(4, 30) <= input(8);
output(4, 31) <= input(9);
output(4, 32) <= input(64);
output(4, 33) <= input(62);
output(4, 34) <= input(53);
output(4, 35) <= input(54);
output(4, 36) <= input(55);
output(4, 37) <= input(56);
output(4, 38) <= input(57);
output(4, 39) <= input(58);
output(4, 40) <= input(33);
output(4, 41) <= input(34);
output(4, 42) <= input(35);
output(4, 43) <= input(36);
output(4, 44) <= input(37);
output(4, 45) <= input(38);
output(4, 46) <= input(39);
output(4, 47) <= input(40);
output(4, 48) <= input(62);
output(4, 49) <= input(53);
output(4, 50) <= input(54);
output(4, 51) <= input(55);
output(4, 52) <= input(56);
output(4, 53) <= input(57);
output(4, 54) <= input(58);
output(4, 55) <= input(33);
output(4, 56) <= input(34);
output(4, 57) <= input(35);
output(4, 58) <= input(36);
output(4, 59) <= input(37);
output(4, 60) <= input(38);
output(4, 61) <= input(39);
output(4, 62) <= input(40);
output(4, 63) <= input(41);
output(4, 64) <= input(60);
output(4, 65) <= input(61);
output(4, 66) <= input(31);
output(4, 67) <= input(32);
output(4, 68) <= input(0);
output(4, 69) <= input(1);
output(4, 70) <= input(2);
output(4, 71) <= input(3);
output(4, 72) <= input(4);
output(4, 73) <= input(5);
output(4, 74) <= input(6);
output(4, 75) <= input(7);
output(4, 76) <= input(8);
output(4, 77) <= input(9);
output(4, 78) <= input(10);
output(4, 79) <= input(11);
output(4, 80) <= input(53);
output(4, 81) <= input(54);
output(4, 82) <= input(55);
output(4, 83) <= input(56);
output(4, 84) <= input(57);
output(4, 85) <= input(58);
output(4, 86) <= input(33);
output(4, 87) <= input(34);
output(4, 88) <= input(35);
output(4, 89) <= input(36);
output(4, 90) <= input(37);
output(4, 91) <= input(38);
output(4, 92) <= input(39);
output(4, 93) <= input(40);
output(4, 94) <= input(41);
output(4, 95) <= input(42);
output(4, 96) <= input(61);
output(4, 97) <= input(31);
output(4, 98) <= input(32);
output(4, 99) <= input(0);
output(4, 100) <= input(1);
output(4, 101) <= input(2);
output(4, 102) <= input(3);
output(4, 103) <= input(4);
output(4, 104) <= input(5);
output(4, 105) <= input(6);
output(4, 106) <= input(7);
output(4, 107) <= input(8);
output(4, 108) <= input(9);
output(4, 109) <= input(10);
output(4, 110) <= input(11);
output(4, 111) <= input(12);
output(4, 112) <= input(31);
output(4, 113) <= input(32);
output(4, 114) <= input(0);
output(4, 115) <= input(1);
output(4, 116) <= input(2);
output(4, 117) <= input(3);
output(4, 118) <= input(4);
output(4, 119) <= input(5);
output(4, 120) <= input(6);
output(4, 121) <= input(7);
output(4, 122) <= input(8);
output(4, 123) <= input(9);
output(4, 124) <= input(10);
output(4, 125) <= input(11);
output(4, 126) <= input(12);
output(4, 127) <= input(13);
output(4, 128) <= input(55);
output(4, 129) <= input(56);
output(4, 130) <= input(57);
output(4, 131) <= input(58);
output(4, 132) <= input(33);
output(4, 133) <= input(34);
output(4, 134) <= input(35);
output(4, 135) <= input(36);
output(4, 136) <= input(37);
output(4, 137) <= input(38);
output(4, 138) <= input(39);
output(4, 139) <= input(40);
output(4, 140) <= input(41);
output(4, 141) <= input(42);
output(4, 142) <= input(43);
output(4, 143) <= input(44);
output(4, 144) <= input(32);
output(4, 145) <= input(0);
output(4, 146) <= input(1);
output(4, 147) <= input(2);
output(4, 148) <= input(3);
output(4, 149) <= input(4);
output(4, 150) <= input(5);
output(4, 151) <= input(6);
output(4, 152) <= input(7);
output(4, 153) <= input(8);
output(4, 154) <= input(9);
output(4, 155) <= input(10);
output(4, 156) <= input(11);
output(4, 157) <= input(12);
output(4, 158) <= input(13);
output(4, 159) <= input(14);
output(4, 160) <= input(56);
output(4, 161) <= input(57);
output(4, 162) <= input(58);
output(4, 163) <= input(33);
output(4, 164) <= input(34);
output(4, 165) <= input(35);
output(4, 166) <= input(36);
output(4, 167) <= input(37);
output(4, 168) <= input(38);
output(4, 169) <= input(39);
output(4, 170) <= input(40);
output(4, 171) <= input(41);
output(4, 172) <= input(42);
output(4, 173) <= input(43);
output(4, 174) <= input(44);
output(4, 175) <= input(45);
output(4, 176) <= input(57);
output(4, 177) <= input(58);
output(4, 178) <= input(33);
output(4, 179) <= input(34);
output(4, 180) <= input(35);
output(4, 181) <= input(36);
output(4, 182) <= input(37);
output(4, 183) <= input(38);
output(4, 184) <= input(39);
output(4, 185) <= input(40);
output(4, 186) <= input(41);
output(4, 187) <= input(42);
output(4, 188) <= input(43);
output(4, 189) <= input(44);
output(4, 190) <= input(45);
output(4, 191) <= input(46);
output(4, 192) <= input(1);
output(4, 193) <= input(2);
output(4, 194) <= input(3);
output(4, 195) <= input(4);
output(4, 196) <= input(5);
output(4, 197) <= input(6);
output(4, 198) <= input(7);
output(4, 199) <= input(8);
output(4, 200) <= input(9);
output(4, 201) <= input(10);
output(4, 202) <= input(11);
output(4, 203) <= input(12);
output(4, 204) <= input(13);
output(4, 205) <= input(14);
output(4, 206) <= input(15);
output(4, 207) <= input(16);
output(4, 208) <= input(58);
output(4, 209) <= input(33);
output(4, 210) <= input(34);
output(4, 211) <= input(35);
output(4, 212) <= input(36);
output(4, 213) <= input(37);
output(4, 214) <= input(38);
output(4, 215) <= input(39);
output(4, 216) <= input(40);
output(4, 217) <= input(41);
output(4, 218) <= input(42);
output(4, 219) <= input(43);
output(4, 220) <= input(44);
output(4, 221) <= input(45);
output(4, 222) <= input(46);
output(4, 223) <= input(47);
output(4, 224) <= input(2);
output(4, 225) <= input(3);
output(4, 226) <= input(4);
output(4, 227) <= input(5);
output(4, 228) <= input(6);
output(4, 229) <= input(7);
output(4, 230) <= input(8);
output(4, 231) <= input(9);
output(4, 232) <= input(10);
output(4, 233) <= input(11);
output(4, 234) <= input(12);
output(4, 235) <= input(13);
output(4, 236) <= input(14);
output(4, 237) <= input(15);
output(4, 238) <= input(16);
output(4, 239) <= input(17);
output(4, 240) <= input(3);
output(4, 241) <= input(4);
output(4, 242) <= input(5);
output(4, 243) <= input(6);
output(4, 244) <= input(7);
output(4, 245) <= input(8);
output(4, 246) <= input(9);
output(4, 247) <= input(10);
output(4, 248) <= input(11);
output(4, 249) <= input(12);
output(4, 250) <= input(13);
output(4, 251) <= input(14);
output(4, 252) <= input(15);
output(4, 253) <= input(16);
output(4, 254) <= input(17);
output(4, 255) <= input(18);
output(5, 0) <= input(66);
output(5, 1) <= input(63);
output(5, 2) <= input(64);
output(5, 3) <= input(62);
output(5, 4) <= input(53);
output(5, 5) <= input(54);
output(5, 6) <= input(55);
output(5, 7) <= input(56);
output(5, 8) <= input(57);
output(5, 9) <= input(58);
output(5, 10) <= input(33);
output(5, 11) <= input(34);
output(5, 12) <= input(35);
output(5, 13) <= input(36);
output(5, 14) <= input(37);
output(5, 15) <= input(38);
output(5, 16) <= input(67);
output(5, 17) <= input(65);
output(5, 18) <= input(59);
output(5, 19) <= input(60);
output(5, 20) <= input(61);
output(5, 21) <= input(31);
output(5, 22) <= input(32);
output(5, 23) <= input(0);
output(5, 24) <= input(1);
output(5, 25) <= input(2);
output(5, 26) <= input(3);
output(5, 27) <= input(4);
output(5, 28) <= input(5);
output(5, 29) <= input(6);
output(5, 30) <= input(7);
output(5, 31) <= input(8);
output(5, 32) <= input(63);
output(5, 33) <= input(64);
output(5, 34) <= input(62);
output(5, 35) <= input(53);
output(5, 36) <= input(54);
output(5, 37) <= input(55);
output(5, 38) <= input(56);
output(5, 39) <= input(57);
output(5, 40) <= input(58);
output(5, 41) <= input(33);
output(5, 42) <= input(34);
output(5, 43) <= input(35);
output(5, 44) <= input(36);
output(5, 45) <= input(37);
output(5, 46) <= input(38);
output(5, 47) <= input(39);
output(5, 48) <= input(65);
output(5, 49) <= input(59);
output(5, 50) <= input(60);
output(5, 51) <= input(61);
output(5, 52) <= input(31);
output(5, 53) <= input(32);
output(5, 54) <= input(0);
output(5, 55) <= input(1);
output(5, 56) <= input(2);
output(5, 57) <= input(3);
output(5, 58) <= input(4);
output(5, 59) <= input(5);
output(5, 60) <= input(6);
output(5, 61) <= input(7);
output(5, 62) <= input(8);
output(5, 63) <= input(9);
output(5, 64) <= input(64);
output(5, 65) <= input(62);
output(5, 66) <= input(53);
output(5, 67) <= input(54);
output(5, 68) <= input(55);
output(5, 69) <= input(56);
output(5, 70) <= input(57);
output(5, 71) <= input(58);
output(5, 72) <= input(33);
output(5, 73) <= input(34);
output(5, 74) <= input(35);
output(5, 75) <= input(36);
output(5, 76) <= input(37);
output(5, 77) <= input(38);
output(5, 78) <= input(39);
output(5, 79) <= input(40);
output(5, 80) <= input(59);
output(5, 81) <= input(60);
output(5, 82) <= input(61);
output(5, 83) <= input(31);
output(5, 84) <= input(32);
output(5, 85) <= input(0);
output(5, 86) <= input(1);
output(5, 87) <= input(2);
output(5, 88) <= input(3);
output(5, 89) <= input(4);
output(5, 90) <= input(5);
output(5, 91) <= input(6);
output(5, 92) <= input(7);
output(5, 93) <= input(8);
output(5, 94) <= input(9);
output(5, 95) <= input(10);
output(5, 96) <= input(62);
output(5, 97) <= input(53);
output(5, 98) <= input(54);
output(5, 99) <= input(55);
output(5, 100) <= input(56);
output(5, 101) <= input(57);
output(5, 102) <= input(58);
output(5, 103) <= input(33);
output(5, 104) <= input(34);
output(5, 105) <= input(35);
output(5, 106) <= input(36);
output(5, 107) <= input(37);
output(5, 108) <= input(38);
output(5, 109) <= input(39);
output(5, 110) <= input(40);
output(5, 111) <= input(41);
output(5, 112) <= input(53);
output(5, 113) <= input(54);
output(5, 114) <= input(55);
output(5, 115) <= input(56);
output(5, 116) <= input(57);
output(5, 117) <= input(58);
output(5, 118) <= input(33);
output(5, 119) <= input(34);
output(5, 120) <= input(35);
output(5, 121) <= input(36);
output(5, 122) <= input(37);
output(5, 123) <= input(38);
output(5, 124) <= input(39);
output(5, 125) <= input(40);
output(5, 126) <= input(41);
output(5, 127) <= input(42);
output(5, 128) <= input(61);
output(5, 129) <= input(31);
output(5, 130) <= input(32);
output(5, 131) <= input(0);
output(5, 132) <= input(1);
output(5, 133) <= input(2);
output(5, 134) <= input(3);
output(5, 135) <= input(4);
output(5, 136) <= input(5);
output(5, 137) <= input(6);
output(5, 138) <= input(7);
output(5, 139) <= input(8);
output(5, 140) <= input(9);
output(5, 141) <= input(10);
output(5, 142) <= input(11);
output(5, 143) <= input(12);
output(5, 144) <= input(54);
output(5, 145) <= input(55);
output(5, 146) <= input(56);
output(5, 147) <= input(57);
output(5, 148) <= input(58);
output(5, 149) <= input(33);
output(5, 150) <= input(34);
output(5, 151) <= input(35);
output(5, 152) <= input(36);
output(5, 153) <= input(37);
output(5, 154) <= input(38);
output(5, 155) <= input(39);
output(5, 156) <= input(40);
output(5, 157) <= input(41);
output(5, 158) <= input(42);
output(5, 159) <= input(43);
output(5, 160) <= input(31);
output(5, 161) <= input(32);
output(5, 162) <= input(0);
output(5, 163) <= input(1);
output(5, 164) <= input(2);
output(5, 165) <= input(3);
output(5, 166) <= input(4);
output(5, 167) <= input(5);
output(5, 168) <= input(6);
output(5, 169) <= input(7);
output(5, 170) <= input(8);
output(5, 171) <= input(9);
output(5, 172) <= input(10);
output(5, 173) <= input(11);
output(5, 174) <= input(12);
output(5, 175) <= input(13);
output(5, 176) <= input(55);
output(5, 177) <= input(56);
output(5, 178) <= input(57);
output(5, 179) <= input(58);
output(5, 180) <= input(33);
output(5, 181) <= input(34);
output(5, 182) <= input(35);
output(5, 183) <= input(36);
output(5, 184) <= input(37);
output(5, 185) <= input(38);
output(5, 186) <= input(39);
output(5, 187) <= input(40);
output(5, 188) <= input(41);
output(5, 189) <= input(42);
output(5, 190) <= input(43);
output(5, 191) <= input(44);
output(5, 192) <= input(32);
output(5, 193) <= input(0);
output(5, 194) <= input(1);
output(5, 195) <= input(2);
output(5, 196) <= input(3);
output(5, 197) <= input(4);
output(5, 198) <= input(5);
output(5, 199) <= input(6);
output(5, 200) <= input(7);
output(5, 201) <= input(8);
output(5, 202) <= input(9);
output(5, 203) <= input(10);
output(5, 204) <= input(11);
output(5, 205) <= input(12);
output(5, 206) <= input(13);
output(5, 207) <= input(14);
output(5, 208) <= input(56);
output(5, 209) <= input(57);
output(5, 210) <= input(58);
output(5, 211) <= input(33);
output(5, 212) <= input(34);
output(5, 213) <= input(35);
output(5, 214) <= input(36);
output(5, 215) <= input(37);
output(5, 216) <= input(38);
output(5, 217) <= input(39);
output(5, 218) <= input(40);
output(5, 219) <= input(41);
output(5, 220) <= input(42);
output(5, 221) <= input(43);
output(5, 222) <= input(44);
output(5, 223) <= input(45);
output(5, 224) <= input(0);
output(5, 225) <= input(1);
output(5, 226) <= input(2);
output(5, 227) <= input(3);
output(5, 228) <= input(4);
output(5, 229) <= input(5);
output(5, 230) <= input(6);
output(5, 231) <= input(7);
output(5, 232) <= input(8);
output(5, 233) <= input(9);
output(5, 234) <= input(10);
output(5, 235) <= input(11);
output(5, 236) <= input(12);
output(5, 237) <= input(13);
output(5, 238) <= input(14);
output(5, 239) <= input(15);
output(5, 240) <= input(1);
output(5, 241) <= input(2);
output(5, 242) <= input(3);
output(5, 243) <= input(4);
output(5, 244) <= input(5);
output(5, 245) <= input(6);
output(5, 246) <= input(7);
output(5, 247) <= input(8);
output(5, 248) <= input(9);
output(5, 249) <= input(10);
output(5, 250) <= input(11);
output(5, 251) <= input(12);
output(5, 252) <= input(13);
output(5, 253) <= input(14);
output(5, 254) <= input(15);
output(5, 255) <= input(16);
when "0001" =>
output(0, 0) <= input(0);
output(0, 1) <= input(1);
output(0, 2) <= input(2);
output(0, 3) <= input(3);
output(0, 4) <= input(4);
output(0, 5) <= input(5);
output(0, 6) <= input(6);
output(0, 7) <= input(7);
output(0, 8) <= input(8);
output(0, 9) <= input(9);
output(0, 10) <= input(10);
output(0, 11) <= input(11);
output(0, 12) <= input(12);
output(0, 13) <= input(13);
output(0, 14) <= input(14);
output(0, 15) <= input(15);
output(0, 16) <= input(16);
output(0, 17) <= input(17);
output(0, 18) <= input(18);
output(0, 19) <= input(19);
output(0, 20) <= input(20);
output(0, 21) <= input(21);
output(0, 22) <= input(22);
output(0, 23) <= input(23);
output(0, 24) <= input(24);
output(0, 25) <= input(25);
output(0, 26) <= input(26);
output(0, 27) <= input(27);
output(0, 28) <= input(28);
output(0, 29) <= input(29);
output(0, 30) <= input(30);
output(0, 31) <= input(31);
output(0, 32) <= input(1);
output(0, 33) <= input(2);
output(0, 34) <= input(3);
output(0, 35) <= input(4);
output(0, 36) <= input(5);
output(0, 37) <= input(6);
output(0, 38) <= input(7);
output(0, 39) <= input(8);
output(0, 40) <= input(9);
output(0, 41) <= input(10);
output(0, 42) <= input(11);
output(0, 43) <= input(12);
output(0, 44) <= input(13);
output(0, 45) <= input(14);
output(0, 46) <= input(15);
output(0, 47) <= input(32);
output(0, 48) <= input(17);
output(0, 49) <= input(18);
output(0, 50) <= input(19);
output(0, 51) <= input(20);
output(0, 52) <= input(21);
output(0, 53) <= input(22);
output(0, 54) <= input(23);
output(0, 55) <= input(24);
output(0, 56) <= input(25);
output(0, 57) <= input(26);
output(0, 58) <= input(27);
output(0, 59) <= input(28);
output(0, 60) <= input(29);
output(0, 61) <= input(30);
output(0, 62) <= input(31);
output(0, 63) <= input(33);
output(0, 64) <= input(2);
output(0, 65) <= input(3);
output(0, 66) <= input(4);
output(0, 67) <= input(5);
output(0, 68) <= input(6);
output(0, 69) <= input(7);
output(0, 70) <= input(8);
output(0, 71) <= input(9);
output(0, 72) <= input(10);
output(0, 73) <= input(11);
output(0, 74) <= input(12);
output(0, 75) <= input(13);
output(0, 76) <= input(14);
output(0, 77) <= input(15);
output(0, 78) <= input(32);
output(0, 79) <= input(34);
output(0, 80) <= input(18);
output(0, 81) <= input(19);
output(0, 82) <= input(20);
output(0, 83) <= input(21);
output(0, 84) <= input(22);
output(0, 85) <= input(23);
output(0, 86) <= input(24);
output(0, 87) <= input(25);
output(0, 88) <= input(26);
output(0, 89) <= input(27);
output(0, 90) <= input(28);
output(0, 91) <= input(29);
output(0, 92) <= input(30);
output(0, 93) <= input(31);
output(0, 94) <= input(33);
output(0, 95) <= input(35);
output(0, 96) <= input(3);
output(0, 97) <= input(4);
output(0, 98) <= input(5);
output(0, 99) <= input(6);
output(0, 100) <= input(7);
output(0, 101) <= input(8);
output(0, 102) <= input(9);
output(0, 103) <= input(10);
output(0, 104) <= input(11);
output(0, 105) <= input(12);
output(0, 106) <= input(13);
output(0, 107) <= input(14);
output(0, 108) <= input(15);
output(0, 109) <= input(32);
output(0, 110) <= input(34);
output(0, 111) <= input(36);
output(0, 112) <= input(19);
output(0, 113) <= input(20);
output(0, 114) <= input(21);
output(0, 115) <= input(22);
output(0, 116) <= input(23);
output(0, 117) <= input(24);
output(0, 118) <= input(25);
output(0, 119) <= input(26);
output(0, 120) <= input(27);
output(0, 121) <= input(28);
output(0, 122) <= input(29);
output(0, 123) <= input(30);
output(0, 124) <= input(31);
output(0, 125) <= input(33);
output(0, 126) <= input(35);
output(0, 127) <= input(37);
output(0, 128) <= input(4);
output(0, 129) <= input(5);
output(0, 130) <= input(6);
output(0, 131) <= input(7);
output(0, 132) <= input(8);
output(0, 133) <= input(9);
output(0, 134) <= input(10);
output(0, 135) <= input(11);
output(0, 136) <= input(12);
output(0, 137) <= input(13);
output(0, 138) <= input(14);
output(0, 139) <= input(15);
output(0, 140) <= input(32);
output(0, 141) <= input(34);
output(0, 142) <= input(36);
output(0, 143) <= input(38);
output(0, 144) <= input(20);
output(0, 145) <= input(21);
output(0, 146) <= input(22);
output(0, 147) <= input(23);
output(0, 148) <= input(24);
output(0, 149) <= input(25);
output(0, 150) <= input(26);
output(0, 151) <= input(27);
output(0, 152) <= input(28);
output(0, 153) <= input(29);
output(0, 154) <= input(30);
output(0, 155) <= input(31);
output(0, 156) <= input(33);
output(0, 157) <= input(35);
output(0, 158) <= input(37);
output(0, 159) <= input(39);
output(0, 160) <= input(5);
output(0, 161) <= input(6);
output(0, 162) <= input(7);
output(0, 163) <= input(8);
output(0, 164) <= input(9);
output(0, 165) <= input(10);
output(0, 166) <= input(11);
output(0, 167) <= input(12);
output(0, 168) <= input(13);
output(0, 169) <= input(14);
output(0, 170) <= input(15);
output(0, 171) <= input(32);
output(0, 172) <= input(34);
output(0, 173) <= input(36);
output(0, 174) <= input(38);
output(0, 175) <= input(40);
output(0, 176) <= input(21);
output(0, 177) <= input(22);
output(0, 178) <= input(23);
output(0, 179) <= input(24);
output(0, 180) <= input(25);
output(0, 181) <= input(26);
output(0, 182) <= input(27);
output(0, 183) <= input(28);
output(0, 184) <= input(29);
output(0, 185) <= input(30);
output(0, 186) <= input(31);
output(0, 187) <= input(33);
output(0, 188) <= input(35);
output(0, 189) <= input(37);
output(0, 190) <= input(39);
output(0, 191) <= input(41);
output(0, 192) <= input(6);
output(0, 193) <= input(7);
output(0, 194) <= input(8);
output(0, 195) <= input(9);
output(0, 196) <= input(10);
output(0, 197) <= input(11);
output(0, 198) <= input(12);
output(0, 199) <= input(13);
output(0, 200) <= input(14);
output(0, 201) <= input(15);
output(0, 202) <= input(32);
output(0, 203) <= input(34);
output(0, 204) <= input(36);
output(0, 205) <= input(38);
output(0, 206) <= input(40);
output(0, 207) <= input(42);
output(0, 208) <= input(22);
output(0, 209) <= input(23);
output(0, 210) <= input(24);
output(0, 211) <= input(25);
output(0, 212) <= input(26);
output(0, 213) <= input(27);
output(0, 214) <= input(28);
output(0, 215) <= input(29);
output(0, 216) <= input(30);
output(0, 217) <= input(31);
output(0, 218) <= input(33);
output(0, 219) <= input(35);
output(0, 220) <= input(37);
output(0, 221) <= input(39);
output(0, 222) <= input(41);
output(0, 223) <= input(43);
output(0, 224) <= input(7);
output(0, 225) <= input(8);
output(0, 226) <= input(9);
output(0, 227) <= input(10);
output(0, 228) <= input(11);
output(0, 229) <= input(12);
output(0, 230) <= input(13);
output(0, 231) <= input(14);
output(0, 232) <= input(15);
output(0, 233) <= input(32);
output(0, 234) <= input(34);
output(0, 235) <= input(36);
output(0, 236) <= input(38);
output(0, 237) <= input(40);
output(0, 238) <= input(42);
output(0, 239) <= input(44);
output(0, 240) <= input(23);
output(0, 241) <= input(24);
output(0, 242) <= input(25);
output(0, 243) <= input(26);
output(0, 244) <= input(27);
output(0, 245) <= input(28);
output(0, 246) <= input(29);
output(0, 247) <= input(30);
output(0, 248) <= input(31);
output(0, 249) <= input(33);
output(0, 250) <= input(35);
output(0, 251) <= input(37);
output(0, 252) <= input(39);
output(0, 253) <= input(41);
output(0, 254) <= input(43);
output(0, 255) <= input(45);
output(1, 0) <= input(46);
output(1, 1) <= input(47);
output(1, 2) <= input(16);
output(1, 3) <= input(17);
output(1, 4) <= input(18);
output(1, 5) <= input(19);
output(1, 6) <= input(20);
output(1, 7) <= input(21);
output(1, 8) <= input(22);
output(1, 9) <= input(23);
output(1, 10) <= input(24);
output(1, 11) <= input(25);
output(1, 12) <= input(26);
output(1, 13) <= input(27);
output(1, 14) <= input(28);
output(1, 15) <= input(29);
output(1, 16) <= input(48);
output(1, 17) <= input(0);
output(1, 18) <= input(1);
output(1, 19) <= input(2);
output(1, 20) <= input(3);
output(1, 21) <= input(4);
output(1, 22) <= input(5);
output(1, 23) <= input(6);
output(1, 24) <= input(7);
output(1, 25) <= input(8);
output(1, 26) <= input(9);
output(1, 27) <= input(10);
output(1, 28) <= input(11);
output(1, 29) <= input(12);
output(1, 30) <= input(13);
output(1, 31) <= input(14);
output(1, 32) <= input(47);
output(1, 33) <= input(16);
output(1, 34) <= input(17);
output(1, 35) <= input(18);
output(1, 36) <= input(19);
output(1, 37) <= input(20);
output(1, 38) <= input(21);
output(1, 39) <= input(22);
output(1, 40) <= input(23);
output(1, 41) <= input(24);
output(1, 42) <= input(25);
output(1, 43) <= input(26);
output(1, 44) <= input(27);
output(1, 45) <= input(28);
output(1, 46) <= input(29);
output(1, 47) <= input(30);
output(1, 48) <= input(0);
output(1, 49) <= input(1);
output(1, 50) <= input(2);
output(1, 51) <= input(3);
output(1, 52) <= input(4);
output(1, 53) <= input(5);
output(1, 54) <= input(6);
output(1, 55) <= input(7);
output(1, 56) <= input(8);
output(1, 57) <= input(9);
output(1, 58) <= input(10);
output(1, 59) <= input(11);
output(1, 60) <= input(12);
output(1, 61) <= input(13);
output(1, 62) <= input(14);
output(1, 63) <= input(15);
output(1, 64) <= input(16);
output(1, 65) <= input(17);
output(1, 66) <= input(18);
output(1, 67) <= input(19);
output(1, 68) <= input(20);
output(1, 69) <= input(21);
output(1, 70) <= input(22);
output(1, 71) <= input(23);
output(1, 72) <= input(24);
output(1, 73) <= input(25);
output(1, 74) <= input(26);
output(1, 75) <= input(27);
output(1, 76) <= input(28);
output(1, 77) <= input(29);
output(1, 78) <= input(30);
output(1, 79) <= input(31);
output(1, 80) <= input(1);
output(1, 81) <= input(2);
output(1, 82) <= input(3);
output(1, 83) <= input(4);
output(1, 84) <= input(5);
output(1, 85) <= input(6);
output(1, 86) <= input(7);
output(1, 87) <= input(8);
output(1, 88) <= input(9);
output(1, 89) <= input(10);
output(1, 90) <= input(11);
output(1, 91) <= input(12);
output(1, 92) <= input(13);
output(1, 93) <= input(14);
output(1, 94) <= input(15);
output(1, 95) <= input(32);
output(1, 96) <= input(17);
output(1, 97) <= input(18);
output(1, 98) <= input(19);
output(1, 99) <= input(20);
output(1, 100) <= input(21);
output(1, 101) <= input(22);
output(1, 102) <= input(23);
output(1, 103) <= input(24);
output(1, 104) <= input(25);
output(1, 105) <= input(26);
output(1, 106) <= input(27);
output(1, 107) <= input(28);
output(1, 108) <= input(29);
output(1, 109) <= input(30);
output(1, 110) <= input(31);
output(1, 111) <= input(33);
output(1, 112) <= input(2);
output(1, 113) <= input(3);
output(1, 114) <= input(4);
output(1, 115) <= input(5);
output(1, 116) <= input(6);
output(1, 117) <= input(7);
output(1, 118) <= input(8);
output(1, 119) <= input(9);
output(1, 120) <= input(10);
output(1, 121) <= input(11);
output(1, 122) <= input(12);
output(1, 123) <= input(13);
output(1, 124) <= input(14);
output(1, 125) <= input(15);
output(1, 126) <= input(32);
output(1, 127) <= input(34);
output(1, 128) <= input(2);
output(1, 129) <= input(3);
output(1, 130) <= input(4);
output(1, 131) <= input(5);
output(1, 132) <= input(6);
output(1, 133) <= input(7);
output(1, 134) <= input(8);
output(1, 135) <= input(9);
output(1, 136) <= input(10);
output(1, 137) <= input(11);
output(1, 138) <= input(12);
output(1, 139) <= input(13);
output(1, 140) <= input(14);
output(1, 141) <= input(15);
output(1, 142) <= input(32);
output(1, 143) <= input(34);
output(1, 144) <= input(18);
output(1, 145) <= input(19);
output(1, 146) <= input(20);
output(1, 147) <= input(21);
output(1, 148) <= input(22);
output(1, 149) <= input(23);
output(1, 150) <= input(24);
output(1, 151) <= input(25);
output(1, 152) <= input(26);
output(1, 153) <= input(27);
output(1, 154) <= input(28);
output(1, 155) <= input(29);
output(1, 156) <= input(30);
output(1, 157) <= input(31);
output(1, 158) <= input(33);
output(1, 159) <= input(35);
output(1, 160) <= input(3);
output(1, 161) <= input(4);
output(1, 162) <= input(5);
output(1, 163) <= input(6);
output(1, 164) <= input(7);
output(1, 165) <= input(8);
output(1, 166) <= input(9);
output(1, 167) <= input(10);
output(1, 168) <= input(11);
output(1, 169) <= input(12);
output(1, 170) <= input(13);
output(1, 171) <= input(14);
output(1, 172) <= input(15);
output(1, 173) <= input(32);
output(1, 174) <= input(34);
output(1, 175) <= input(36);
output(1, 176) <= input(19);
output(1, 177) <= input(20);
output(1, 178) <= input(21);
output(1, 179) <= input(22);
output(1, 180) <= input(23);
output(1, 181) <= input(24);
output(1, 182) <= input(25);
output(1, 183) <= input(26);
output(1, 184) <= input(27);
output(1, 185) <= input(28);
output(1, 186) <= input(29);
output(1, 187) <= input(30);
output(1, 188) <= input(31);
output(1, 189) <= input(33);
output(1, 190) <= input(35);
output(1, 191) <= input(37);
output(1, 192) <= input(4);
output(1, 193) <= input(5);
output(1, 194) <= input(6);
output(1, 195) <= input(7);
output(1, 196) <= input(8);
output(1, 197) <= input(9);
output(1, 198) <= input(10);
output(1, 199) <= input(11);
output(1, 200) <= input(12);
output(1, 201) <= input(13);
output(1, 202) <= input(14);
output(1, 203) <= input(15);
output(1, 204) <= input(32);
output(1, 205) <= input(34);
output(1, 206) <= input(36);
output(1, 207) <= input(38);
output(1, 208) <= input(20);
output(1, 209) <= input(21);
output(1, 210) <= input(22);
output(1, 211) <= input(23);
output(1, 212) <= input(24);
output(1, 213) <= input(25);
output(1, 214) <= input(26);
output(1, 215) <= input(27);
output(1, 216) <= input(28);
output(1, 217) <= input(29);
output(1, 218) <= input(30);
output(1, 219) <= input(31);
output(1, 220) <= input(33);
output(1, 221) <= input(35);
output(1, 222) <= input(37);
output(1, 223) <= input(39);
output(1, 224) <= input(5);
output(1, 225) <= input(6);
output(1, 226) <= input(7);
output(1, 227) <= input(8);
output(1, 228) <= input(9);
output(1, 229) <= input(10);
output(1, 230) <= input(11);
output(1, 231) <= input(12);
output(1, 232) <= input(13);
output(1, 233) <= input(14);
output(1, 234) <= input(15);
output(1, 235) <= input(32);
output(1, 236) <= input(34);
output(1, 237) <= input(36);
output(1, 238) <= input(38);
output(1, 239) <= input(40);
output(1, 240) <= input(21);
output(1, 241) <= input(22);
output(1, 242) <= input(23);
output(1, 243) <= input(24);
output(1, 244) <= input(25);
output(1, 245) <= input(26);
output(1, 246) <= input(27);
output(1, 247) <= input(28);
output(1, 248) <= input(29);
output(1, 249) <= input(30);
output(1, 250) <= input(31);
output(1, 251) <= input(33);
output(1, 252) <= input(35);
output(1, 253) <= input(37);
output(1, 254) <= input(39);
output(1, 255) <= input(41);
output(2, 0) <= input(49);
output(2, 1) <= input(46);
output(2, 2) <= input(47);
output(2, 3) <= input(16);
output(2, 4) <= input(17);
output(2, 5) <= input(18);
output(2, 6) <= input(19);
output(2, 7) <= input(20);
output(2, 8) <= input(21);
output(2, 9) <= input(22);
output(2, 10) <= input(23);
output(2, 11) <= input(24);
output(2, 12) <= input(25);
output(2, 13) <= input(26);
output(2, 14) <= input(27);
output(2, 15) <= input(28);
output(2, 16) <= input(50);
output(2, 17) <= input(48);
output(2, 18) <= input(0);
output(2, 19) <= input(1);
output(2, 20) <= input(2);
output(2, 21) <= input(3);
output(2, 22) <= input(4);
output(2, 23) <= input(5);
output(2, 24) <= input(6);
output(2, 25) <= input(7);
output(2, 26) <= input(8);
output(2, 27) <= input(9);
output(2, 28) <= input(10);
output(2, 29) <= input(11);
output(2, 30) <= input(12);
output(2, 31) <= input(13);
output(2, 32) <= input(46);
output(2, 33) <= input(47);
output(2, 34) <= input(16);
output(2, 35) <= input(17);
output(2, 36) <= input(18);
output(2, 37) <= input(19);
output(2, 38) <= input(20);
output(2, 39) <= input(21);
output(2, 40) <= input(22);
output(2, 41) <= input(23);
output(2, 42) <= input(24);
output(2, 43) <= input(25);
output(2, 44) <= input(26);
output(2, 45) <= input(27);
output(2, 46) <= input(28);
output(2, 47) <= input(29);
output(2, 48) <= input(48);
output(2, 49) <= input(0);
output(2, 50) <= input(1);
output(2, 51) <= input(2);
output(2, 52) <= input(3);
output(2, 53) <= input(4);
output(2, 54) <= input(5);
output(2, 55) <= input(6);
output(2, 56) <= input(7);
output(2, 57) <= input(8);
output(2, 58) <= input(9);
output(2, 59) <= input(10);
output(2, 60) <= input(11);
output(2, 61) <= input(12);
output(2, 62) <= input(13);
output(2, 63) <= input(14);
output(2, 64) <= input(48);
output(2, 65) <= input(0);
output(2, 66) <= input(1);
output(2, 67) <= input(2);
output(2, 68) <= input(3);
output(2, 69) <= input(4);
output(2, 70) <= input(5);
output(2, 71) <= input(6);
output(2, 72) <= input(7);
output(2, 73) <= input(8);
output(2, 74) <= input(9);
output(2, 75) <= input(10);
output(2, 76) <= input(11);
output(2, 77) <= input(12);
output(2, 78) <= input(13);
output(2, 79) <= input(14);
output(2, 80) <= input(47);
output(2, 81) <= input(16);
output(2, 82) <= input(17);
output(2, 83) <= input(18);
output(2, 84) <= input(19);
output(2, 85) <= input(20);
output(2, 86) <= input(21);
output(2, 87) <= input(22);
output(2, 88) <= input(23);
output(2, 89) <= input(24);
output(2, 90) <= input(25);
output(2, 91) <= input(26);
output(2, 92) <= input(27);
output(2, 93) <= input(28);
output(2, 94) <= input(29);
output(2, 95) <= input(30);
output(2, 96) <= input(0);
output(2, 97) <= input(1);
output(2, 98) <= input(2);
output(2, 99) <= input(3);
output(2, 100) <= input(4);
output(2, 101) <= input(5);
output(2, 102) <= input(6);
output(2, 103) <= input(7);
output(2, 104) <= input(8);
output(2, 105) <= input(9);
output(2, 106) <= input(10);
output(2, 107) <= input(11);
output(2, 108) <= input(12);
output(2, 109) <= input(13);
output(2, 110) <= input(14);
output(2, 111) <= input(15);
output(2, 112) <= input(16);
output(2, 113) <= input(17);
output(2, 114) <= input(18);
output(2, 115) <= input(19);
output(2, 116) <= input(20);
output(2, 117) <= input(21);
output(2, 118) <= input(22);
output(2, 119) <= input(23);
output(2, 120) <= input(24);
output(2, 121) <= input(25);
output(2, 122) <= input(26);
output(2, 123) <= input(27);
output(2, 124) <= input(28);
output(2, 125) <= input(29);
output(2, 126) <= input(30);
output(2, 127) <= input(31);
output(2, 128) <= input(16);
output(2, 129) <= input(17);
output(2, 130) <= input(18);
output(2, 131) <= input(19);
output(2, 132) <= input(20);
output(2, 133) <= input(21);
output(2, 134) <= input(22);
output(2, 135) <= input(23);
output(2, 136) <= input(24);
output(2, 137) <= input(25);
output(2, 138) <= input(26);
output(2, 139) <= input(27);
output(2, 140) <= input(28);
output(2, 141) <= input(29);
output(2, 142) <= input(30);
output(2, 143) <= input(31);
output(2, 144) <= input(1);
output(2, 145) <= input(2);
output(2, 146) <= input(3);
output(2, 147) <= input(4);
output(2, 148) <= input(5);
output(2, 149) <= input(6);
output(2, 150) <= input(7);
output(2, 151) <= input(8);
output(2, 152) <= input(9);
output(2, 153) <= input(10);
output(2, 154) <= input(11);
output(2, 155) <= input(12);
output(2, 156) <= input(13);
output(2, 157) <= input(14);
output(2, 158) <= input(15);
output(2, 159) <= input(32);
output(2, 160) <= input(17);
output(2, 161) <= input(18);
output(2, 162) <= input(19);
output(2, 163) <= input(20);
output(2, 164) <= input(21);
output(2, 165) <= input(22);
output(2, 166) <= input(23);
output(2, 167) <= input(24);
output(2, 168) <= input(25);
output(2, 169) <= input(26);
output(2, 170) <= input(27);
output(2, 171) <= input(28);
output(2, 172) <= input(29);
output(2, 173) <= input(30);
output(2, 174) <= input(31);
output(2, 175) <= input(33);
output(2, 176) <= input(2);
output(2, 177) <= input(3);
output(2, 178) <= input(4);
output(2, 179) <= input(5);
output(2, 180) <= input(6);
output(2, 181) <= input(7);
output(2, 182) <= input(8);
output(2, 183) <= input(9);
output(2, 184) <= input(10);
output(2, 185) <= input(11);
output(2, 186) <= input(12);
output(2, 187) <= input(13);
output(2, 188) <= input(14);
output(2, 189) <= input(15);
output(2, 190) <= input(32);
output(2, 191) <= input(34);
output(2, 192) <= input(2);
output(2, 193) <= input(3);
output(2, 194) <= input(4);
output(2, 195) <= input(5);
output(2, 196) <= input(6);
output(2, 197) <= input(7);
output(2, 198) <= input(8);
output(2, 199) <= input(9);
output(2, 200) <= input(10);
output(2, 201) <= input(11);
output(2, 202) <= input(12);
output(2, 203) <= input(13);
output(2, 204) <= input(14);
output(2, 205) <= input(15);
output(2, 206) <= input(32);
output(2, 207) <= input(34);
output(2, 208) <= input(18);
output(2, 209) <= input(19);
output(2, 210) <= input(20);
output(2, 211) <= input(21);
output(2, 212) <= input(22);
output(2, 213) <= input(23);
output(2, 214) <= input(24);
output(2, 215) <= input(25);
output(2, 216) <= input(26);
output(2, 217) <= input(27);
output(2, 218) <= input(28);
output(2, 219) <= input(29);
output(2, 220) <= input(30);
output(2, 221) <= input(31);
output(2, 222) <= input(33);
output(2, 223) <= input(35);
output(2, 224) <= input(3);
output(2, 225) <= input(4);
output(2, 226) <= input(5);
output(2, 227) <= input(6);
output(2, 228) <= input(7);
output(2, 229) <= input(8);
output(2, 230) <= input(9);
output(2, 231) <= input(10);
output(2, 232) <= input(11);
output(2, 233) <= input(12);
output(2, 234) <= input(13);
output(2, 235) <= input(14);
output(2, 236) <= input(15);
output(2, 237) <= input(32);
output(2, 238) <= input(34);
output(2, 239) <= input(36);
output(2, 240) <= input(19);
output(2, 241) <= input(20);
output(2, 242) <= input(21);
output(2, 243) <= input(22);
output(2, 244) <= input(23);
output(2, 245) <= input(24);
output(2, 246) <= input(25);
output(2, 247) <= input(26);
output(2, 248) <= input(27);
output(2, 249) <= input(28);
output(2, 250) <= input(29);
output(2, 251) <= input(30);
output(2, 252) <= input(31);
output(2, 253) <= input(33);
output(2, 254) <= input(35);
output(2, 255) <= input(37);
output(3, 0) <= input(51);
output(3, 1) <= input(49);
output(3, 2) <= input(46);
output(3, 3) <= input(47);
output(3, 4) <= input(16);
output(3, 5) <= input(17);
output(3, 6) <= input(18);
output(3, 7) <= input(19);
output(3, 8) <= input(20);
output(3, 9) <= input(21);
output(3, 10) <= input(22);
output(3, 11) <= input(23);
output(3, 12) <= input(24);
output(3, 13) <= input(25);
output(3, 14) <= input(26);
output(3, 15) <= input(27);
output(3, 16) <= input(52);
output(3, 17) <= input(50);
output(3, 18) <= input(48);
output(3, 19) <= input(0);
output(3, 20) <= input(1);
output(3, 21) <= input(2);
output(3, 22) <= input(3);
output(3, 23) <= input(4);
output(3, 24) <= input(5);
output(3, 25) <= input(6);
output(3, 26) <= input(7);
output(3, 27) <= input(8);
output(3, 28) <= input(9);
output(3, 29) <= input(10);
output(3, 30) <= input(11);
output(3, 31) <= input(12);
output(3, 32) <= input(52);
output(3, 33) <= input(50);
output(3, 34) <= input(48);
output(3, 35) <= input(0);
output(3, 36) <= input(1);
output(3, 37) <= input(2);
output(3, 38) <= input(3);
output(3, 39) <= input(4);
output(3, 40) <= input(5);
output(3, 41) <= input(6);
output(3, 42) <= input(7);
output(3, 43) <= input(8);
output(3, 44) <= input(9);
output(3, 45) <= input(10);
output(3, 46) <= input(11);
output(3, 47) <= input(12);
output(3, 48) <= input(49);
output(3, 49) <= input(46);
output(3, 50) <= input(47);
output(3, 51) <= input(16);
output(3, 52) <= input(17);
output(3, 53) <= input(18);
output(3, 54) <= input(19);
output(3, 55) <= input(20);
output(3, 56) <= input(21);
output(3, 57) <= input(22);
output(3, 58) <= input(23);
output(3, 59) <= input(24);
output(3, 60) <= input(25);
output(3, 61) <= input(26);
output(3, 62) <= input(27);
output(3, 63) <= input(28);
output(3, 64) <= input(50);
output(3, 65) <= input(48);
output(3, 66) <= input(0);
output(3, 67) <= input(1);
output(3, 68) <= input(2);
output(3, 69) <= input(3);
output(3, 70) <= input(4);
output(3, 71) <= input(5);
output(3, 72) <= input(6);
output(3, 73) <= input(7);
output(3, 74) <= input(8);
output(3, 75) <= input(9);
output(3, 76) <= input(10);
output(3, 77) <= input(11);
output(3, 78) <= input(12);
output(3, 79) <= input(13);
output(3, 80) <= input(50);
output(3, 81) <= input(48);
output(3, 82) <= input(0);
output(3, 83) <= input(1);
output(3, 84) <= input(2);
output(3, 85) <= input(3);
output(3, 86) <= input(4);
output(3, 87) <= input(5);
output(3, 88) <= input(6);
output(3, 89) <= input(7);
output(3, 90) <= input(8);
output(3, 91) <= input(9);
output(3, 92) <= input(10);
output(3, 93) <= input(11);
output(3, 94) <= input(12);
output(3, 95) <= input(13);
output(3, 96) <= input(46);
output(3, 97) <= input(47);
output(3, 98) <= input(16);
output(3, 99) <= input(17);
output(3, 100) <= input(18);
output(3, 101) <= input(19);
output(3, 102) <= input(20);
output(3, 103) <= input(21);
output(3, 104) <= input(22);
output(3, 105) <= input(23);
output(3, 106) <= input(24);
output(3, 107) <= input(25);
output(3, 108) <= input(26);
output(3, 109) <= input(27);
output(3, 110) <= input(28);
output(3, 111) <= input(29);
output(3, 112) <= input(48);
output(3, 113) <= input(0);
output(3, 114) <= input(1);
output(3, 115) <= input(2);
output(3, 116) <= input(3);
output(3, 117) <= input(4);
output(3, 118) <= input(5);
output(3, 119) <= input(6);
output(3, 120) <= input(7);
output(3, 121) <= input(8);
output(3, 122) <= input(9);
output(3, 123) <= input(10);
output(3, 124) <= input(11);
output(3, 125) <= input(12);
output(3, 126) <= input(13);
output(3, 127) <= input(14);
output(3, 128) <= input(48);
output(3, 129) <= input(0);
output(3, 130) <= input(1);
output(3, 131) <= input(2);
output(3, 132) <= input(3);
output(3, 133) <= input(4);
output(3, 134) <= input(5);
output(3, 135) <= input(6);
output(3, 136) <= input(7);
output(3, 137) <= input(8);
output(3, 138) <= input(9);
output(3, 139) <= input(10);
output(3, 140) <= input(11);
output(3, 141) <= input(12);
output(3, 142) <= input(13);
output(3, 143) <= input(14);
output(3, 144) <= input(47);
output(3, 145) <= input(16);
output(3, 146) <= input(17);
output(3, 147) <= input(18);
output(3, 148) <= input(19);
output(3, 149) <= input(20);
output(3, 150) <= input(21);
output(3, 151) <= input(22);
output(3, 152) <= input(23);
output(3, 153) <= input(24);
output(3, 154) <= input(25);
output(3, 155) <= input(26);
output(3, 156) <= input(27);
output(3, 157) <= input(28);
output(3, 158) <= input(29);
output(3, 159) <= input(30);
output(3, 160) <= input(47);
output(3, 161) <= input(16);
output(3, 162) <= input(17);
output(3, 163) <= input(18);
output(3, 164) <= input(19);
output(3, 165) <= input(20);
output(3, 166) <= input(21);
output(3, 167) <= input(22);
output(3, 168) <= input(23);
output(3, 169) <= input(24);
output(3, 170) <= input(25);
output(3, 171) <= input(26);
output(3, 172) <= input(27);
output(3, 173) <= input(28);
output(3, 174) <= input(29);
output(3, 175) <= input(30);
output(3, 176) <= input(0);
output(3, 177) <= input(1);
output(3, 178) <= input(2);
output(3, 179) <= input(3);
output(3, 180) <= input(4);
output(3, 181) <= input(5);
output(3, 182) <= input(6);
output(3, 183) <= input(7);
output(3, 184) <= input(8);
output(3, 185) <= input(9);
output(3, 186) <= input(10);
output(3, 187) <= input(11);
output(3, 188) <= input(12);
output(3, 189) <= input(13);
output(3, 190) <= input(14);
output(3, 191) <= input(15);
output(3, 192) <= input(16);
output(3, 193) <= input(17);
output(3, 194) <= input(18);
output(3, 195) <= input(19);
output(3, 196) <= input(20);
output(3, 197) <= input(21);
output(3, 198) <= input(22);
output(3, 199) <= input(23);
output(3, 200) <= input(24);
output(3, 201) <= input(25);
output(3, 202) <= input(26);
output(3, 203) <= input(27);
output(3, 204) <= input(28);
output(3, 205) <= input(29);
output(3, 206) <= input(30);
output(3, 207) <= input(31);
output(3, 208) <= input(16);
output(3, 209) <= input(17);
output(3, 210) <= input(18);
output(3, 211) <= input(19);
output(3, 212) <= input(20);
output(3, 213) <= input(21);
output(3, 214) <= input(22);
output(3, 215) <= input(23);
output(3, 216) <= input(24);
output(3, 217) <= input(25);
output(3, 218) <= input(26);
output(3, 219) <= input(27);
output(3, 220) <= input(28);
output(3, 221) <= input(29);
output(3, 222) <= input(30);
output(3, 223) <= input(31);
output(3, 224) <= input(1);
output(3, 225) <= input(2);
output(3, 226) <= input(3);
output(3, 227) <= input(4);
output(3, 228) <= input(5);
output(3, 229) <= input(6);
output(3, 230) <= input(7);
output(3, 231) <= input(8);
output(3, 232) <= input(9);
output(3, 233) <= input(10);
output(3, 234) <= input(11);
output(3, 235) <= input(12);
output(3, 236) <= input(13);
output(3, 237) <= input(14);
output(3, 238) <= input(15);
output(3, 239) <= input(32);
output(3, 240) <= input(17);
output(3, 241) <= input(18);
output(3, 242) <= input(19);
output(3, 243) <= input(20);
output(3, 244) <= input(21);
output(3, 245) <= input(22);
output(3, 246) <= input(23);
output(3, 247) <= input(24);
output(3, 248) <= input(25);
output(3, 249) <= input(26);
output(3, 250) <= input(27);
output(3, 251) <= input(28);
output(3, 252) <= input(29);
output(3, 253) <= input(30);
output(3, 254) <= input(31);
output(3, 255) <= input(33);
output(4, 0) <= input(53);
output(4, 1) <= input(51);
output(4, 2) <= input(49);
output(4, 3) <= input(46);
output(4, 4) <= input(47);
output(4, 5) <= input(16);
output(4, 6) <= input(17);
output(4, 7) <= input(18);
output(4, 8) <= input(19);
output(4, 9) <= input(20);
output(4, 10) <= input(21);
output(4, 11) <= input(22);
output(4, 12) <= input(23);
output(4, 13) <= input(24);
output(4, 14) <= input(25);
output(4, 15) <= input(26);
output(4, 16) <= input(54);
output(4, 17) <= input(52);
output(4, 18) <= input(50);
output(4, 19) <= input(48);
output(4, 20) <= input(0);
output(4, 21) <= input(1);
output(4, 22) <= input(2);
output(4, 23) <= input(3);
output(4, 24) <= input(4);
output(4, 25) <= input(5);
output(4, 26) <= input(6);
output(4, 27) <= input(7);
output(4, 28) <= input(8);
output(4, 29) <= input(9);
output(4, 30) <= input(10);
output(4, 31) <= input(11);
output(4, 32) <= input(54);
output(4, 33) <= input(52);
output(4, 34) <= input(50);
output(4, 35) <= input(48);
output(4, 36) <= input(0);
output(4, 37) <= input(1);
output(4, 38) <= input(2);
output(4, 39) <= input(3);
output(4, 40) <= input(4);
output(4, 41) <= input(5);
output(4, 42) <= input(6);
output(4, 43) <= input(7);
output(4, 44) <= input(8);
output(4, 45) <= input(9);
output(4, 46) <= input(10);
output(4, 47) <= input(11);
output(4, 48) <= input(51);
output(4, 49) <= input(49);
output(4, 50) <= input(46);
output(4, 51) <= input(47);
output(4, 52) <= input(16);
output(4, 53) <= input(17);
output(4, 54) <= input(18);
output(4, 55) <= input(19);
output(4, 56) <= input(20);
output(4, 57) <= input(21);
output(4, 58) <= input(22);
output(4, 59) <= input(23);
output(4, 60) <= input(24);
output(4, 61) <= input(25);
output(4, 62) <= input(26);
output(4, 63) <= input(27);
output(4, 64) <= input(51);
output(4, 65) <= input(49);
output(4, 66) <= input(46);
output(4, 67) <= input(47);
output(4, 68) <= input(16);
output(4, 69) <= input(17);
output(4, 70) <= input(18);
output(4, 71) <= input(19);
output(4, 72) <= input(20);
output(4, 73) <= input(21);
output(4, 74) <= input(22);
output(4, 75) <= input(23);
output(4, 76) <= input(24);
output(4, 77) <= input(25);
output(4, 78) <= input(26);
output(4, 79) <= input(27);
output(4, 80) <= input(52);
output(4, 81) <= input(50);
output(4, 82) <= input(48);
output(4, 83) <= input(0);
output(4, 84) <= input(1);
output(4, 85) <= input(2);
output(4, 86) <= input(3);
output(4, 87) <= input(4);
output(4, 88) <= input(5);
output(4, 89) <= input(6);
output(4, 90) <= input(7);
output(4, 91) <= input(8);
output(4, 92) <= input(9);
output(4, 93) <= input(10);
output(4, 94) <= input(11);
output(4, 95) <= input(12);
output(4, 96) <= input(52);
output(4, 97) <= input(50);
output(4, 98) <= input(48);
output(4, 99) <= input(0);
output(4, 100) <= input(1);
output(4, 101) <= input(2);
output(4, 102) <= input(3);
output(4, 103) <= input(4);
output(4, 104) <= input(5);
output(4, 105) <= input(6);
output(4, 106) <= input(7);
output(4, 107) <= input(8);
output(4, 108) <= input(9);
output(4, 109) <= input(10);
output(4, 110) <= input(11);
output(4, 111) <= input(12);
output(4, 112) <= input(49);
output(4, 113) <= input(46);
output(4, 114) <= input(47);
output(4, 115) <= input(16);
output(4, 116) <= input(17);
output(4, 117) <= input(18);
output(4, 118) <= input(19);
output(4, 119) <= input(20);
output(4, 120) <= input(21);
output(4, 121) <= input(22);
output(4, 122) <= input(23);
output(4, 123) <= input(24);
output(4, 124) <= input(25);
output(4, 125) <= input(26);
output(4, 126) <= input(27);
output(4, 127) <= input(28);
output(4, 128) <= input(49);
output(4, 129) <= input(46);
output(4, 130) <= input(47);
output(4, 131) <= input(16);
output(4, 132) <= input(17);
output(4, 133) <= input(18);
output(4, 134) <= input(19);
output(4, 135) <= input(20);
output(4, 136) <= input(21);
output(4, 137) <= input(22);
output(4, 138) <= input(23);
output(4, 139) <= input(24);
output(4, 140) <= input(25);
output(4, 141) <= input(26);
output(4, 142) <= input(27);
output(4, 143) <= input(28);
output(4, 144) <= input(50);
output(4, 145) <= input(48);
output(4, 146) <= input(0);
output(4, 147) <= input(1);
output(4, 148) <= input(2);
output(4, 149) <= input(3);
output(4, 150) <= input(4);
output(4, 151) <= input(5);
output(4, 152) <= input(6);
output(4, 153) <= input(7);
output(4, 154) <= input(8);
output(4, 155) <= input(9);
output(4, 156) <= input(10);
output(4, 157) <= input(11);
output(4, 158) <= input(12);
output(4, 159) <= input(13);
output(4, 160) <= input(50);
output(4, 161) <= input(48);
output(4, 162) <= input(0);
output(4, 163) <= input(1);
output(4, 164) <= input(2);
output(4, 165) <= input(3);
output(4, 166) <= input(4);
output(4, 167) <= input(5);
output(4, 168) <= input(6);
output(4, 169) <= input(7);
output(4, 170) <= input(8);
output(4, 171) <= input(9);
output(4, 172) <= input(10);
output(4, 173) <= input(11);
output(4, 174) <= input(12);
output(4, 175) <= input(13);
output(4, 176) <= input(46);
output(4, 177) <= input(47);
output(4, 178) <= input(16);
output(4, 179) <= input(17);
output(4, 180) <= input(18);
output(4, 181) <= input(19);
output(4, 182) <= input(20);
output(4, 183) <= input(21);
output(4, 184) <= input(22);
output(4, 185) <= input(23);
output(4, 186) <= input(24);
output(4, 187) <= input(25);
output(4, 188) <= input(26);
output(4, 189) <= input(27);
output(4, 190) <= input(28);
output(4, 191) <= input(29);
output(4, 192) <= input(46);
output(4, 193) <= input(47);
output(4, 194) <= input(16);
output(4, 195) <= input(17);
output(4, 196) <= input(18);
output(4, 197) <= input(19);
output(4, 198) <= input(20);
output(4, 199) <= input(21);
output(4, 200) <= input(22);
output(4, 201) <= input(23);
output(4, 202) <= input(24);
output(4, 203) <= input(25);
output(4, 204) <= input(26);
output(4, 205) <= input(27);
output(4, 206) <= input(28);
output(4, 207) <= input(29);
output(4, 208) <= input(48);
output(4, 209) <= input(0);
output(4, 210) <= input(1);
output(4, 211) <= input(2);
output(4, 212) <= input(3);
output(4, 213) <= input(4);
output(4, 214) <= input(5);
output(4, 215) <= input(6);
output(4, 216) <= input(7);
output(4, 217) <= input(8);
output(4, 218) <= input(9);
output(4, 219) <= input(10);
output(4, 220) <= input(11);
output(4, 221) <= input(12);
output(4, 222) <= input(13);
output(4, 223) <= input(14);
output(4, 224) <= input(48);
output(4, 225) <= input(0);
output(4, 226) <= input(1);
output(4, 227) <= input(2);
output(4, 228) <= input(3);
output(4, 229) <= input(4);
output(4, 230) <= input(5);
output(4, 231) <= input(6);
output(4, 232) <= input(7);
output(4, 233) <= input(8);
output(4, 234) <= input(9);
output(4, 235) <= input(10);
output(4, 236) <= input(11);
output(4, 237) <= input(12);
output(4, 238) <= input(13);
output(4, 239) <= input(14);
output(4, 240) <= input(47);
output(4, 241) <= input(16);
output(4, 242) <= input(17);
output(4, 243) <= input(18);
output(4, 244) <= input(19);
output(4, 245) <= input(20);
output(4, 246) <= input(21);
output(4, 247) <= input(22);
output(4, 248) <= input(23);
output(4, 249) <= input(24);
output(4, 250) <= input(25);
output(4, 251) <= input(26);
output(4, 252) <= input(27);
output(4, 253) <= input(28);
output(4, 254) <= input(29);
output(4, 255) <= input(30);
output(5, 0) <= input(55);
output(5, 1) <= input(53);
output(5, 2) <= input(51);
output(5, 3) <= input(49);
output(5, 4) <= input(46);
output(5, 5) <= input(47);
output(5, 6) <= input(16);
output(5, 7) <= input(17);
output(5, 8) <= input(18);
output(5, 9) <= input(19);
output(5, 10) <= input(20);
output(5, 11) <= input(21);
output(5, 12) <= input(22);
output(5, 13) <= input(23);
output(5, 14) <= input(24);
output(5, 15) <= input(25);
output(5, 16) <= input(55);
output(5, 17) <= input(53);
output(5, 18) <= input(51);
output(5, 19) <= input(49);
output(5, 20) <= input(46);
output(5, 21) <= input(47);
output(5, 22) <= input(16);
output(5, 23) <= input(17);
output(5, 24) <= input(18);
output(5, 25) <= input(19);
output(5, 26) <= input(20);
output(5, 27) <= input(21);
output(5, 28) <= input(22);
output(5, 29) <= input(23);
output(5, 30) <= input(24);
output(5, 31) <= input(25);
output(5, 32) <= input(56);
output(5, 33) <= input(54);
output(5, 34) <= input(52);
output(5, 35) <= input(50);
output(5, 36) <= input(48);
output(5, 37) <= input(0);
output(5, 38) <= input(1);
output(5, 39) <= input(2);
output(5, 40) <= input(3);
output(5, 41) <= input(4);
output(5, 42) <= input(5);
output(5, 43) <= input(6);
output(5, 44) <= input(7);
output(5, 45) <= input(8);
output(5, 46) <= input(9);
output(5, 47) <= input(10);
output(5, 48) <= input(56);
output(5, 49) <= input(54);
output(5, 50) <= input(52);
output(5, 51) <= input(50);
output(5, 52) <= input(48);
output(5, 53) <= input(0);
output(5, 54) <= input(1);
output(5, 55) <= input(2);
output(5, 56) <= input(3);
output(5, 57) <= input(4);
output(5, 58) <= input(5);
output(5, 59) <= input(6);
output(5, 60) <= input(7);
output(5, 61) <= input(8);
output(5, 62) <= input(9);
output(5, 63) <= input(10);
output(5, 64) <= input(56);
output(5, 65) <= input(54);
output(5, 66) <= input(52);
output(5, 67) <= input(50);
output(5, 68) <= input(48);
output(5, 69) <= input(0);
output(5, 70) <= input(1);
output(5, 71) <= input(2);
output(5, 72) <= input(3);
output(5, 73) <= input(4);
output(5, 74) <= input(5);
output(5, 75) <= input(6);
output(5, 76) <= input(7);
output(5, 77) <= input(8);
output(5, 78) <= input(9);
output(5, 79) <= input(10);
output(5, 80) <= input(53);
output(5, 81) <= input(51);
output(5, 82) <= input(49);
output(5, 83) <= input(46);
output(5, 84) <= input(47);
output(5, 85) <= input(16);
output(5, 86) <= input(17);
output(5, 87) <= input(18);
output(5, 88) <= input(19);
output(5, 89) <= input(20);
output(5, 90) <= input(21);
output(5, 91) <= input(22);
output(5, 92) <= input(23);
output(5, 93) <= input(24);
output(5, 94) <= input(25);
output(5, 95) <= input(26);
output(5, 96) <= input(53);
output(5, 97) <= input(51);
output(5, 98) <= input(49);
output(5, 99) <= input(46);
output(5, 100) <= input(47);
output(5, 101) <= input(16);
output(5, 102) <= input(17);
output(5, 103) <= input(18);
output(5, 104) <= input(19);
output(5, 105) <= input(20);
output(5, 106) <= input(21);
output(5, 107) <= input(22);
output(5, 108) <= input(23);
output(5, 109) <= input(24);
output(5, 110) <= input(25);
output(5, 111) <= input(26);
output(5, 112) <= input(54);
output(5, 113) <= input(52);
output(5, 114) <= input(50);
output(5, 115) <= input(48);
output(5, 116) <= input(0);
output(5, 117) <= input(1);
output(5, 118) <= input(2);
output(5, 119) <= input(3);
output(5, 120) <= input(4);
output(5, 121) <= input(5);
output(5, 122) <= input(6);
output(5, 123) <= input(7);
output(5, 124) <= input(8);
output(5, 125) <= input(9);
output(5, 126) <= input(10);
output(5, 127) <= input(11);
output(5, 128) <= input(54);
output(5, 129) <= input(52);
output(5, 130) <= input(50);
output(5, 131) <= input(48);
output(5, 132) <= input(0);
output(5, 133) <= input(1);
output(5, 134) <= input(2);
output(5, 135) <= input(3);
output(5, 136) <= input(4);
output(5, 137) <= input(5);
output(5, 138) <= input(6);
output(5, 139) <= input(7);
output(5, 140) <= input(8);
output(5, 141) <= input(9);
output(5, 142) <= input(10);
output(5, 143) <= input(11);
output(5, 144) <= input(54);
output(5, 145) <= input(52);
output(5, 146) <= input(50);
output(5, 147) <= input(48);
output(5, 148) <= input(0);
output(5, 149) <= input(1);
output(5, 150) <= input(2);
output(5, 151) <= input(3);
output(5, 152) <= input(4);
output(5, 153) <= input(5);
output(5, 154) <= input(6);
output(5, 155) <= input(7);
output(5, 156) <= input(8);
output(5, 157) <= input(9);
output(5, 158) <= input(10);
output(5, 159) <= input(11);
output(5, 160) <= input(51);
output(5, 161) <= input(49);
output(5, 162) <= input(46);
output(5, 163) <= input(47);
output(5, 164) <= input(16);
output(5, 165) <= input(17);
output(5, 166) <= input(18);
output(5, 167) <= input(19);
output(5, 168) <= input(20);
output(5, 169) <= input(21);
output(5, 170) <= input(22);
output(5, 171) <= input(23);
output(5, 172) <= input(24);
output(5, 173) <= input(25);
output(5, 174) <= input(26);
output(5, 175) <= input(27);
output(5, 176) <= input(51);
output(5, 177) <= input(49);
output(5, 178) <= input(46);
output(5, 179) <= input(47);
output(5, 180) <= input(16);
output(5, 181) <= input(17);
output(5, 182) <= input(18);
output(5, 183) <= input(19);
output(5, 184) <= input(20);
output(5, 185) <= input(21);
output(5, 186) <= input(22);
output(5, 187) <= input(23);
output(5, 188) <= input(24);
output(5, 189) <= input(25);
output(5, 190) <= input(26);
output(5, 191) <= input(27);
output(5, 192) <= input(51);
output(5, 193) <= input(49);
output(5, 194) <= input(46);
output(5, 195) <= input(47);
output(5, 196) <= input(16);
output(5, 197) <= input(17);
output(5, 198) <= input(18);
output(5, 199) <= input(19);
output(5, 200) <= input(20);
output(5, 201) <= input(21);
output(5, 202) <= input(22);
output(5, 203) <= input(23);
output(5, 204) <= input(24);
output(5, 205) <= input(25);
output(5, 206) <= input(26);
output(5, 207) <= input(27);
output(5, 208) <= input(52);
output(5, 209) <= input(50);
output(5, 210) <= input(48);
output(5, 211) <= input(0);
output(5, 212) <= input(1);
output(5, 213) <= input(2);
output(5, 214) <= input(3);
output(5, 215) <= input(4);
output(5, 216) <= input(5);
output(5, 217) <= input(6);
output(5, 218) <= input(7);
output(5, 219) <= input(8);
output(5, 220) <= input(9);
output(5, 221) <= input(10);
output(5, 222) <= input(11);
output(5, 223) <= input(12);
output(5, 224) <= input(52);
output(5, 225) <= input(50);
output(5, 226) <= input(48);
output(5, 227) <= input(0);
output(5, 228) <= input(1);
output(5, 229) <= input(2);
output(5, 230) <= input(3);
output(5, 231) <= input(4);
output(5, 232) <= input(5);
output(5, 233) <= input(6);
output(5, 234) <= input(7);
output(5, 235) <= input(8);
output(5, 236) <= input(9);
output(5, 237) <= input(10);
output(5, 238) <= input(11);
output(5, 239) <= input(12);
output(5, 240) <= input(49);
output(5, 241) <= input(46);
output(5, 242) <= input(47);
output(5, 243) <= input(16);
output(5, 244) <= input(17);
output(5, 245) <= input(18);
output(5, 246) <= input(19);
output(5, 247) <= input(20);
output(5, 248) <= input(21);
output(5, 249) <= input(22);
output(5, 250) <= input(23);
output(5, 251) <= input(24);
output(5, 252) <= input(25);
output(5, 253) <= input(26);
output(5, 254) <= input(27);
output(5, 255) <= input(28);
when "0010" =>
output(0, 0) <= input(0);
output(0, 1) <= input(1);
output(0, 2) <= input(2);
output(0, 3) <= input(3);
output(0, 4) <= input(4);
output(0, 5) <= input(5);
output(0, 6) <= input(6);
output(0, 7) <= input(7);
output(0, 8) <= input(8);
output(0, 9) <= input(9);
output(0, 10) <= input(10);
output(0, 11) <= input(11);
output(0, 12) <= input(12);
output(0, 13) <= input(13);
output(0, 14) <= input(14);
output(0, 15) <= input(15);
output(0, 16) <= input(0);
output(0, 17) <= input(1);
output(0, 18) <= input(2);
output(0, 19) <= input(3);
output(0, 20) <= input(4);
output(0, 21) <= input(5);
output(0, 22) <= input(6);
output(0, 23) <= input(7);
output(0, 24) <= input(8);
output(0, 25) <= input(9);
output(0, 26) <= input(10);
output(0, 27) <= input(11);
output(0, 28) <= input(12);
output(0, 29) <= input(13);
output(0, 30) <= input(14);
output(0, 31) <= input(15);
output(0, 32) <= input(0);
output(0, 33) <= input(1);
output(0, 34) <= input(2);
output(0, 35) <= input(3);
output(0, 36) <= input(4);
output(0, 37) <= input(5);
output(0, 38) <= input(6);
output(0, 39) <= input(7);
output(0, 40) <= input(8);
output(0, 41) <= input(9);
output(0, 42) <= input(10);
output(0, 43) <= input(11);
output(0, 44) <= input(12);
output(0, 45) <= input(13);
output(0, 46) <= input(14);
output(0, 47) <= input(15);
output(0, 48) <= input(16);
output(0, 49) <= input(17);
output(0, 50) <= input(18);
output(0, 51) <= input(19);
output(0, 52) <= input(20);
output(0, 53) <= input(21);
output(0, 54) <= input(22);
output(0, 55) <= input(23);
output(0, 56) <= input(24);
output(0, 57) <= input(25);
output(0, 58) <= input(26);
output(0, 59) <= input(27);
output(0, 60) <= input(28);
output(0, 61) <= input(29);
output(0, 62) <= input(30);
output(0, 63) <= input(31);
output(0, 64) <= input(16);
output(0, 65) <= input(17);
output(0, 66) <= input(18);
output(0, 67) <= input(19);
output(0, 68) <= input(20);
output(0, 69) <= input(21);
output(0, 70) <= input(22);
output(0, 71) <= input(23);
output(0, 72) <= input(24);
output(0, 73) <= input(25);
output(0, 74) <= input(26);
output(0, 75) <= input(27);
output(0, 76) <= input(28);
output(0, 77) <= input(29);
output(0, 78) <= input(30);
output(0, 79) <= input(31);
output(0, 80) <= input(16);
output(0, 81) <= input(17);
output(0, 82) <= input(18);
output(0, 83) <= input(19);
output(0, 84) <= input(20);
output(0, 85) <= input(21);
output(0, 86) <= input(22);
output(0, 87) <= input(23);
output(0, 88) <= input(24);
output(0, 89) <= input(25);
output(0, 90) <= input(26);
output(0, 91) <= input(27);
output(0, 92) <= input(28);
output(0, 93) <= input(29);
output(0, 94) <= input(30);
output(0, 95) <= input(31);
output(0, 96) <= input(16);
output(0, 97) <= input(17);
output(0, 98) <= input(18);
output(0, 99) <= input(19);
output(0, 100) <= input(20);
output(0, 101) <= input(21);
output(0, 102) <= input(22);
output(0, 103) <= input(23);
output(0, 104) <= input(24);
output(0, 105) <= input(25);
output(0, 106) <= input(26);
output(0, 107) <= input(27);
output(0, 108) <= input(28);
output(0, 109) <= input(29);
output(0, 110) <= input(30);
output(0, 111) <= input(31);
output(0, 112) <= input(1);
output(0, 113) <= input(2);
output(0, 114) <= input(3);
output(0, 115) <= input(4);
output(0, 116) <= input(5);
output(0, 117) <= input(6);
output(0, 118) <= input(7);
output(0, 119) <= input(8);
output(0, 120) <= input(9);
output(0, 121) <= input(10);
output(0, 122) <= input(11);
output(0, 123) <= input(12);
output(0, 124) <= input(13);
output(0, 125) <= input(14);
output(0, 126) <= input(15);
output(0, 127) <= input(32);
output(0, 128) <= input(1);
output(0, 129) <= input(2);
output(0, 130) <= input(3);
output(0, 131) <= input(4);
output(0, 132) <= input(5);
output(0, 133) <= input(6);
output(0, 134) <= input(7);
output(0, 135) <= input(8);
output(0, 136) <= input(9);
output(0, 137) <= input(10);
output(0, 138) <= input(11);
output(0, 139) <= input(12);
output(0, 140) <= input(13);
output(0, 141) <= input(14);
output(0, 142) <= input(15);
output(0, 143) <= input(32);
output(0, 144) <= input(1);
output(0, 145) <= input(2);
output(0, 146) <= input(3);
output(0, 147) <= input(4);
output(0, 148) <= input(5);
output(0, 149) <= input(6);
output(0, 150) <= input(7);
output(0, 151) <= input(8);
output(0, 152) <= input(9);
output(0, 153) <= input(10);
output(0, 154) <= input(11);
output(0, 155) <= input(12);
output(0, 156) <= input(13);
output(0, 157) <= input(14);
output(0, 158) <= input(15);
output(0, 159) <= input(32);
output(0, 160) <= input(1);
output(0, 161) <= input(2);
output(0, 162) <= input(3);
output(0, 163) <= input(4);
output(0, 164) <= input(5);
output(0, 165) <= input(6);
output(0, 166) <= input(7);
output(0, 167) <= input(8);
output(0, 168) <= input(9);
output(0, 169) <= input(10);
output(0, 170) <= input(11);
output(0, 171) <= input(12);
output(0, 172) <= input(13);
output(0, 173) <= input(14);
output(0, 174) <= input(15);
output(0, 175) <= input(32);
output(0, 176) <= input(17);
output(0, 177) <= input(18);
output(0, 178) <= input(19);
output(0, 179) <= input(20);
output(0, 180) <= input(21);
output(0, 181) <= input(22);
output(0, 182) <= input(23);
output(0, 183) <= input(24);
output(0, 184) <= input(25);
output(0, 185) <= input(26);
output(0, 186) <= input(27);
output(0, 187) <= input(28);
output(0, 188) <= input(29);
output(0, 189) <= input(30);
output(0, 190) <= input(31);
output(0, 191) <= input(33);
output(0, 192) <= input(17);
output(0, 193) <= input(18);
output(0, 194) <= input(19);
output(0, 195) <= input(20);
output(0, 196) <= input(21);
output(0, 197) <= input(22);
output(0, 198) <= input(23);
output(0, 199) <= input(24);
output(0, 200) <= input(25);
output(0, 201) <= input(26);
output(0, 202) <= input(27);
output(0, 203) <= input(28);
output(0, 204) <= input(29);
output(0, 205) <= input(30);
output(0, 206) <= input(31);
output(0, 207) <= input(33);
output(0, 208) <= input(17);
output(0, 209) <= input(18);
output(0, 210) <= input(19);
output(0, 211) <= input(20);
output(0, 212) <= input(21);
output(0, 213) <= input(22);
output(0, 214) <= input(23);
output(0, 215) <= input(24);
output(0, 216) <= input(25);
output(0, 217) <= input(26);
output(0, 218) <= input(27);
output(0, 219) <= input(28);
output(0, 220) <= input(29);
output(0, 221) <= input(30);
output(0, 222) <= input(31);
output(0, 223) <= input(33);
output(0, 224) <= input(17);
output(0, 225) <= input(18);
output(0, 226) <= input(19);
output(0, 227) <= input(20);
output(0, 228) <= input(21);
output(0, 229) <= input(22);
output(0, 230) <= input(23);
output(0, 231) <= input(24);
output(0, 232) <= input(25);
output(0, 233) <= input(26);
output(0, 234) <= input(27);
output(0, 235) <= input(28);
output(0, 236) <= input(29);
output(0, 237) <= input(30);
output(0, 238) <= input(31);
output(0, 239) <= input(33);
output(0, 240) <= input(2);
output(0, 241) <= input(3);
output(0, 242) <= input(4);
output(0, 243) <= input(5);
output(0, 244) <= input(6);
output(0, 245) <= input(7);
output(0, 246) <= input(8);
output(0, 247) <= input(9);
output(0, 248) <= input(10);
output(0, 249) <= input(11);
output(0, 250) <= input(12);
output(0, 251) <= input(13);
output(0, 252) <= input(14);
output(0, 253) <= input(15);
output(0, 254) <= input(32);
output(0, 255) <= input(34);
output(1, 0) <= input(35);
output(1, 1) <= input(16);
output(1, 2) <= input(17);
output(1, 3) <= input(18);
output(1, 4) <= input(19);
output(1, 5) <= input(20);
output(1, 6) <= input(21);
output(1, 7) <= input(22);
output(1, 8) <= input(23);
output(1, 9) <= input(24);
output(1, 10) <= input(25);
output(1, 11) <= input(26);
output(1, 12) <= input(27);
output(1, 13) <= input(28);
output(1, 14) <= input(29);
output(1, 15) <= input(30);
output(1, 16) <= input(35);
output(1, 17) <= input(16);
output(1, 18) <= input(17);
output(1, 19) <= input(18);
output(1, 20) <= input(19);
output(1, 21) <= input(20);
output(1, 22) <= input(21);
output(1, 23) <= input(22);
output(1, 24) <= input(23);
output(1, 25) <= input(24);
output(1, 26) <= input(25);
output(1, 27) <= input(26);
output(1, 28) <= input(27);
output(1, 29) <= input(28);
output(1, 30) <= input(29);
output(1, 31) <= input(30);
output(1, 32) <= input(35);
output(1, 33) <= input(16);
output(1, 34) <= input(17);
output(1, 35) <= input(18);
output(1, 36) <= input(19);
output(1, 37) <= input(20);
output(1, 38) <= input(21);
output(1, 39) <= input(22);
output(1, 40) <= input(23);
output(1, 41) <= input(24);
output(1, 42) <= input(25);
output(1, 43) <= input(26);
output(1, 44) <= input(27);
output(1, 45) <= input(28);
output(1, 46) <= input(29);
output(1, 47) <= input(30);
output(1, 48) <= input(35);
output(1, 49) <= input(16);
output(1, 50) <= input(17);
output(1, 51) <= input(18);
output(1, 52) <= input(19);
output(1, 53) <= input(20);
output(1, 54) <= input(21);
output(1, 55) <= input(22);
output(1, 56) <= input(23);
output(1, 57) <= input(24);
output(1, 58) <= input(25);
output(1, 59) <= input(26);
output(1, 60) <= input(27);
output(1, 61) <= input(28);
output(1, 62) <= input(29);
output(1, 63) <= input(30);
output(1, 64) <= input(35);
output(1, 65) <= input(16);
output(1, 66) <= input(17);
output(1, 67) <= input(18);
output(1, 68) <= input(19);
output(1, 69) <= input(20);
output(1, 70) <= input(21);
output(1, 71) <= input(22);
output(1, 72) <= input(23);
output(1, 73) <= input(24);
output(1, 74) <= input(25);
output(1, 75) <= input(26);
output(1, 76) <= input(27);
output(1, 77) <= input(28);
output(1, 78) <= input(29);
output(1, 79) <= input(30);
output(1, 80) <= input(0);
output(1, 81) <= input(1);
output(1, 82) <= input(2);
output(1, 83) <= input(3);
output(1, 84) <= input(4);
output(1, 85) <= input(5);
output(1, 86) <= input(6);
output(1, 87) <= input(7);
output(1, 88) <= input(8);
output(1, 89) <= input(9);
output(1, 90) <= input(10);
output(1, 91) <= input(11);
output(1, 92) <= input(12);
output(1, 93) <= input(13);
output(1, 94) <= input(14);
output(1, 95) <= input(15);
output(1, 96) <= input(0);
output(1, 97) <= input(1);
output(1, 98) <= input(2);
output(1, 99) <= input(3);
output(1, 100) <= input(4);
output(1, 101) <= input(5);
output(1, 102) <= input(6);
output(1, 103) <= input(7);
output(1, 104) <= input(8);
output(1, 105) <= input(9);
output(1, 106) <= input(10);
output(1, 107) <= input(11);
output(1, 108) <= input(12);
output(1, 109) <= input(13);
output(1, 110) <= input(14);
output(1, 111) <= input(15);
output(1, 112) <= input(0);
output(1, 113) <= input(1);
output(1, 114) <= input(2);
output(1, 115) <= input(3);
output(1, 116) <= input(4);
output(1, 117) <= input(5);
output(1, 118) <= input(6);
output(1, 119) <= input(7);
output(1, 120) <= input(8);
output(1, 121) <= input(9);
output(1, 122) <= input(10);
output(1, 123) <= input(11);
output(1, 124) <= input(12);
output(1, 125) <= input(13);
output(1, 126) <= input(14);
output(1, 127) <= input(15);
output(1, 128) <= input(0);
output(1, 129) <= input(1);
output(1, 130) <= input(2);
output(1, 131) <= input(3);
output(1, 132) <= input(4);
output(1, 133) <= input(5);
output(1, 134) <= input(6);
output(1, 135) <= input(7);
output(1, 136) <= input(8);
output(1, 137) <= input(9);
output(1, 138) <= input(10);
output(1, 139) <= input(11);
output(1, 140) <= input(12);
output(1, 141) <= input(13);
output(1, 142) <= input(14);
output(1, 143) <= input(15);
output(1, 144) <= input(0);
output(1, 145) <= input(1);
output(1, 146) <= input(2);
output(1, 147) <= input(3);
output(1, 148) <= input(4);
output(1, 149) <= input(5);
output(1, 150) <= input(6);
output(1, 151) <= input(7);
output(1, 152) <= input(8);
output(1, 153) <= input(9);
output(1, 154) <= input(10);
output(1, 155) <= input(11);
output(1, 156) <= input(12);
output(1, 157) <= input(13);
output(1, 158) <= input(14);
output(1, 159) <= input(15);
output(1, 160) <= input(16);
output(1, 161) <= input(17);
output(1, 162) <= input(18);
output(1, 163) <= input(19);
output(1, 164) <= input(20);
output(1, 165) <= input(21);
output(1, 166) <= input(22);
output(1, 167) <= input(23);
output(1, 168) <= input(24);
output(1, 169) <= input(25);
output(1, 170) <= input(26);
output(1, 171) <= input(27);
output(1, 172) <= input(28);
output(1, 173) <= input(29);
output(1, 174) <= input(30);
output(1, 175) <= input(31);
output(1, 176) <= input(16);
output(1, 177) <= input(17);
output(1, 178) <= input(18);
output(1, 179) <= input(19);
output(1, 180) <= input(20);
output(1, 181) <= input(21);
output(1, 182) <= input(22);
output(1, 183) <= input(23);
output(1, 184) <= input(24);
output(1, 185) <= input(25);
output(1, 186) <= input(26);
output(1, 187) <= input(27);
output(1, 188) <= input(28);
output(1, 189) <= input(29);
output(1, 190) <= input(30);
output(1, 191) <= input(31);
output(1, 192) <= input(16);
output(1, 193) <= input(17);
output(1, 194) <= input(18);
output(1, 195) <= input(19);
output(1, 196) <= input(20);
output(1, 197) <= input(21);
output(1, 198) <= input(22);
output(1, 199) <= input(23);
output(1, 200) <= input(24);
output(1, 201) <= input(25);
output(1, 202) <= input(26);
output(1, 203) <= input(27);
output(1, 204) <= input(28);
output(1, 205) <= input(29);
output(1, 206) <= input(30);
output(1, 207) <= input(31);
output(1, 208) <= input(16);
output(1, 209) <= input(17);
output(1, 210) <= input(18);
output(1, 211) <= input(19);
output(1, 212) <= input(20);
output(1, 213) <= input(21);
output(1, 214) <= input(22);
output(1, 215) <= input(23);
output(1, 216) <= input(24);
output(1, 217) <= input(25);
output(1, 218) <= input(26);
output(1, 219) <= input(27);
output(1, 220) <= input(28);
output(1, 221) <= input(29);
output(1, 222) <= input(30);
output(1, 223) <= input(31);
output(1, 224) <= input(16);
output(1, 225) <= input(17);
output(1, 226) <= input(18);
output(1, 227) <= input(19);
output(1, 228) <= input(20);
output(1, 229) <= input(21);
output(1, 230) <= input(22);
output(1, 231) <= input(23);
output(1, 232) <= input(24);
output(1, 233) <= input(25);
output(1, 234) <= input(26);
output(1, 235) <= input(27);
output(1, 236) <= input(28);
output(1, 237) <= input(29);
output(1, 238) <= input(30);
output(1, 239) <= input(31);
output(1, 240) <= input(1);
output(1, 241) <= input(2);
output(1, 242) <= input(3);
output(1, 243) <= input(4);
output(1, 244) <= input(5);
output(1, 245) <= input(6);
output(1, 246) <= input(7);
output(1, 247) <= input(8);
output(1, 248) <= input(9);
output(1, 249) <= input(10);
output(1, 250) <= input(11);
output(1, 251) <= input(12);
output(1, 252) <= input(13);
output(1, 253) <= input(14);
output(1, 254) <= input(15);
output(1, 255) <= input(32);
output(2, 0) <= input(36);
output(2, 1) <= input(0);
output(2, 2) <= input(1);
output(2, 3) <= input(2);
output(2, 4) <= input(3);
output(2, 5) <= input(4);
output(2, 6) <= input(5);
output(2, 7) <= input(6);
output(2, 8) <= input(7);
output(2, 9) <= input(8);
output(2, 10) <= input(9);
output(2, 11) <= input(10);
output(2, 12) <= input(11);
output(2, 13) <= input(12);
output(2, 14) <= input(13);
output(2, 15) <= input(14);
output(2, 16) <= input(36);
output(2, 17) <= input(0);
output(2, 18) <= input(1);
output(2, 19) <= input(2);
output(2, 20) <= input(3);
output(2, 21) <= input(4);
output(2, 22) <= input(5);
output(2, 23) <= input(6);
output(2, 24) <= input(7);
output(2, 25) <= input(8);
output(2, 26) <= input(9);
output(2, 27) <= input(10);
output(2, 28) <= input(11);
output(2, 29) <= input(12);
output(2, 30) <= input(13);
output(2, 31) <= input(14);
output(2, 32) <= input(36);
output(2, 33) <= input(0);
output(2, 34) <= input(1);
output(2, 35) <= input(2);
output(2, 36) <= input(3);
output(2, 37) <= input(4);
output(2, 38) <= input(5);
output(2, 39) <= input(6);
output(2, 40) <= input(7);
output(2, 41) <= input(8);
output(2, 42) <= input(9);
output(2, 43) <= input(10);
output(2, 44) <= input(11);
output(2, 45) <= input(12);
output(2, 46) <= input(13);
output(2, 47) <= input(14);
output(2, 48) <= input(36);
output(2, 49) <= input(0);
output(2, 50) <= input(1);
output(2, 51) <= input(2);
output(2, 52) <= input(3);
output(2, 53) <= input(4);
output(2, 54) <= input(5);
output(2, 55) <= input(6);
output(2, 56) <= input(7);
output(2, 57) <= input(8);
output(2, 58) <= input(9);
output(2, 59) <= input(10);
output(2, 60) <= input(11);
output(2, 61) <= input(12);
output(2, 62) <= input(13);
output(2, 63) <= input(14);
output(2, 64) <= input(36);
output(2, 65) <= input(0);
output(2, 66) <= input(1);
output(2, 67) <= input(2);
output(2, 68) <= input(3);
output(2, 69) <= input(4);
output(2, 70) <= input(5);
output(2, 71) <= input(6);
output(2, 72) <= input(7);
output(2, 73) <= input(8);
output(2, 74) <= input(9);
output(2, 75) <= input(10);
output(2, 76) <= input(11);
output(2, 77) <= input(12);
output(2, 78) <= input(13);
output(2, 79) <= input(14);
output(2, 80) <= input(36);
output(2, 81) <= input(0);
output(2, 82) <= input(1);
output(2, 83) <= input(2);
output(2, 84) <= input(3);
output(2, 85) <= input(4);
output(2, 86) <= input(5);
output(2, 87) <= input(6);
output(2, 88) <= input(7);
output(2, 89) <= input(8);
output(2, 90) <= input(9);
output(2, 91) <= input(10);
output(2, 92) <= input(11);
output(2, 93) <= input(12);
output(2, 94) <= input(13);
output(2, 95) <= input(14);
output(2, 96) <= input(36);
output(2, 97) <= input(0);
output(2, 98) <= input(1);
output(2, 99) <= input(2);
output(2, 100) <= input(3);
output(2, 101) <= input(4);
output(2, 102) <= input(5);
output(2, 103) <= input(6);
output(2, 104) <= input(7);
output(2, 105) <= input(8);
output(2, 106) <= input(9);
output(2, 107) <= input(10);
output(2, 108) <= input(11);
output(2, 109) <= input(12);
output(2, 110) <= input(13);
output(2, 111) <= input(14);
output(2, 112) <= input(35);
output(2, 113) <= input(16);
output(2, 114) <= input(17);
output(2, 115) <= input(18);
output(2, 116) <= input(19);
output(2, 117) <= input(20);
output(2, 118) <= input(21);
output(2, 119) <= input(22);
output(2, 120) <= input(23);
output(2, 121) <= input(24);
output(2, 122) <= input(25);
output(2, 123) <= input(26);
output(2, 124) <= input(27);
output(2, 125) <= input(28);
output(2, 126) <= input(29);
output(2, 127) <= input(30);
output(2, 128) <= input(35);
output(2, 129) <= input(16);
output(2, 130) <= input(17);
output(2, 131) <= input(18);
output(2, 132) <= input(19);
output(2, 133) <= input(20);
output(2, 134) <= input(21);
output(2, 135) <= input(22);
output(2, 136) <= input(23);
output(2, 137) <= input(24);
output(2, 138) <= input(25);
output(2, 139) <= input(26);
output(2, 140) <= input(27);
output(2, 141) <= input(28);
output(2, 142) <= input(29);
output(2, 143) <= input(30);
output(2, 144) <= input(35);
output(2, 145) <= input(16);
output(2, 146) <= input(17);
output(2, 147) <= input(18);
output(2, 148) <= input(19);
output(2, 149) <= input(20);
output(2, 150) <= input(21);
output(2, 151) <= input(22);
output(2, 152) <= input(23);
output(2, 153) <= input(24);
output(2, 154) <= input(25);
output(2, 155) <= input(26);
output(2, 156) <= input(27);
output(2, 157) <= input(28);
output(2, 158) <= input(29);
output(2, 159) <= input(30);
output(2, 160) <= input(35);
output(2, 161) <= input(16);
output(2, 162) <= input(17);
output(2, 163) <= input(18);
output(2, 164) <= input(19);
output(2, 165) <= input(20);
output(2, 166) <= input(21);
output(2, 167) <= input(22);
output(2, 168) <= input(23);
output(2, 169) <= input(24);
output(2, 170) <= input(25);
output(2, 171) <= input(26);
output(2, 172) <= input(27);
output(2, 173) <= input(28);
output(2, 174) <= input(29);
output(2, 175) <= input(30);
output(2, 176) <= input(35);
output(2, 177) <= input(16);
output(2, 178) <= input(17);
output(2, 179) <= input(18);
output(2, 180) <= input(19);
output(2, 181) <= input(20);
output(2, 182) <= input(21);
output(2, 183) <= input(22);
output(2, 184) <= input(23);
output(2, 185) <= input(24);
output(2, 186) <= input(25);
output(2, 187) <= input(26);
output(2, 188) <= input(27);
output(2, 189) <= input(28);
output(2, 190) <= input(29);
output(2, 191) <= input(30);
output(2, 192) <= input(35);
output(2, 193) <= input(16);
output(2, 194) <= input(17);
output(2, 195) <= input(18);
output(2, 196) <= input(19);
output(2, 197) <= input(20);
output(2, 198) <= input(21);
output(2, 199) <= input(22);
output(2, 200) <= input(23);
output(2, 201) <= input(24);
output(2, 202) <= input(25);
output(2, 203) <= input(26);
output(2, 204) <= input(27);
output(2, 205) <= input(28);
output(2, 206) <= input(29);
output(2, 207) <= input(30);
output(2, 208) <= input(35);
output(2, 209) <= input(16);
output(2, 210) <= input(17);
output(2, 211) <= input(18);
output(2, 212) <= input(19);
output(2, 213) <= input(20);
output(2, 214) <= input(21);
output(2, 215) <= input(22);
output(2, 216) <= input(23);
output(2, 217) <= input(24);
output(2, 218) <= input(25);
output(2, 219) <= input(26);
output(2, 220) <= input(27);
output(2, 221) <= input(28);
output(2, 222) <= input(29);
output(2, 223) <= input(30);
output(2, 224) <= input(35);
output(2, 225) <= input(16);
output(2, 226) <= input(17);
output(2, 227) <= input(18);
output(2, 228) <= input(19);
output(2, 229) <= input(20);
output(2, 230) <= input(21);
output(2, 231) <= input(22);
output(2, 232) <= input(23);
output(2, 233) <= input(24);
output(2, 234) <= input(25);
output(2, 235) <= input(26);
output(2, 236) <= input(27);
output(2, 237) <= input(28);
output(2, 238) <= input(29);
output(2, 239) <= input(30);
output(2, 240) <= input(0);
output(2, 241) <= input(1);
output(2, 242) <= input(2);
output(2, 243) <= input(3);
output(2, 244) <= input(4);
output(2, 245) <= input(5);
output(2, 246) <= input(6);
output(2, 247) <= input(7);
output(2, 248) <= input(8);
output(2, 249) <= input(9);
output(2, 250) <= input(10);
output(2, 251) <= input(11);
output(2, 252) <= input(12);
output(2, 253) <= input(13);
output(2, 254) <= input(14);
output(2, 255) <= input(15);
output(3, 0) <= input(37);
output(3, 1) <= input(35);
output(3, 2) <= input(16);
output(3, 3) <= input(17);
output(3, 4) <= input(18);
output(3, 5) <= input(19);
output(3, 6) <= input(20);
output(3, 7) <= input(21);
output(3, 8) <= input(22);
output(3, 9) <= input(23);
output(3, 10) <= input(24);
output(3, 11) <= input(25);
output(3, 12) <= input(26);
output(3, 13) <= input(27);
output(3, 14) <= input(28);
output(3, 15) <= input(29);
output(3, 16) <= input(37);
output(3, 17) <= input(35);
output(3, 18) <= input(16);
output(3, 19) <= input(17);
output(3, 20) <= input(18);
output(3, 21) <= input(19);
output(3, 22) <= input(20);
output(3, 23) <= input(21);
output(3, 24) <= input(22);
output(3, 25) <= input(23);
output(3, 26) <= input(24);
output(3, 27) <= input(25);
output(3, 28) <= input(26);
output(3, 29) <= input(27);
output(3, 30) <= input(28);
output(3, 31) <= input(29);
output(3, 32) <= input(37);
output(3, 33) <= input(35);
output(3, 34) <= input(16);
output(3, 35) <= input(17);
output(3, 36) <= input(18);
output(3, 37) <= input(19);
output(3, 38) <= input(20);
output(3, 39) <= input(21);
output(3, 40) <= input(22);
output(3, 41) <= input(23);
output(3, 42) <= input(24);
output(3, 43) <= input(25);
output(3, 44) <= input(26);
output(3, 45) <= input(27);
output(3, 46) <= input(28);
output(3, 47) <= input(29);
output(3, 48) <= input(37);
output(3, 49) <= input(35);
output(3, 50) <= input(16);
output(3, 51) <= input(17);
output(3, 52) <= input(18);
output(3, 53) <= input(19);
output(3, 54) <= input(20);
output(3, 55) <= input(21);
output(3, 56) <= input(22);
output(3, 57) <= input(23);
output(3, 58) <= input(24);
output(3, 59) <= input(25);
output(3, 60) <= input(26);
output(3, 61) <= input(27);
output(3, 62) <= input(28);
output(3, 63) <= input(29);
output(3, 64) <= input(37);
output(3, 65) <= input(35);
output(3, 66) <= input(16);
output(3, 67) <= input(17);
output(3, 68) <= input(18);
output(3, 69) <= input(19);
output(3, 70) <= input(20);
output(3, 71) <= input(21);
output(3, 72) <= input(22);
output(3, 73) <= input(23);
output(3, 74) <= input(24);
output(3, 75) <= input(25);
output(3, 76) <= input(26);
output(3, 77) <= input(27);
output(3, 78) <= input(28);
output(3, 79) <= input(29);
output(3, 80) <= input(37);
output(3, 81) <= input(35);
output(3, 82) <= input(16);
output(3, 83) <= input(17);
output(3, 84) <= input(18);
output(3, 85) <= input(19);
output(3, 86) <= input(20);
output(3, 87) <= input(21);
output(3, 88) <= input(22);
output(3, 89) <= input(23);
output(3, 90) <= input(24);
output(3, 91) <= input(25);
output(3, 92) <= input(26);
output(3, 93) <= input(27);
output(3, 94) <= input(28);
output(3, 95) <= input(29);
output(3, 96) <= input(37);
output(3, 97) <= input(35);
output(3, 98) <= input(16);
output(3, 99) <= input(17);
output(3, 100) <= input(18);
output(3, 101) <= input(19);
output(3, 102) <= input(20);
output(3, 103) <= input(21);
output(3, 104) <= input(22);
output(3, 105) <= input(23);
output(3, 106) <= input(24);
output(3, 107) <= input(25);
output(3, 108) <= input(26);
output(3, 109) <= input(27);
output(3, 110) <= input(28);
output(3, 111) <= input(29);
output(3, 112) <= input(37);
output(3, 113) <= input(35);
output(3, 114) <= input(16);
output(3, 115) <= input(17);
output(3, 116) <= input(18);
output(3, 117) <= input(19);
output(3, 118) <= input(20);
output(3, 119) <= input(21);
output(3, 120) <= input(22);
output(3, 121) <= input(23);
output(3, 122) <= input(24);
output(3, 123) <= input(25);
output(3, 124) <= input(26);
output(3, 125) <= input(27);
output(3, 126) <= input(28);
output(3, 127) <= input(29);
output(3, 128) <= input(37);
output(3, 129) <= input(35);
output(3, 130) <= input(16);
output(3, 131) <= input(17);
output(3, 132) <= input(18);
output(3, 133) <= input(19);
output(3, 134) <= input(20);
output(3, 135) <= input(21);
output(3, 136) <= input(22);
output(3, 137) <= input(23);
output(3, 138) <= input(24);
output(3, 139) <= input(25);
output(3, 140) <= input(26);
output(3, 141) <= input(27);
output(3, 142) <= input(28);
output(3, 143) <= input(29);
output(3, 144) <= input(37);
output(3, 145) <= input(35);
output(3, 146) <= input(16);
output(3, 147) <= input(17);
output(3, 148) <= input(18);
output(3, 149) <= input(19);
output(3, 150) <= input(20);
output(3, 151) <= input(21);
output(3, 152) <= input(22);
output(3, 153) <= input(23);
output(3, 154) <= input(24);
output(3, 155) <= input(25);
output(3, 156) <= input(26);
output(3, 157) <= input(27);
output(3, 158) <= input(28);
output(3, 159) <= input(29);
output(3, 160) <= input(37);
output(3, 161) <= input(35);
output(3, 162) <= input(16);
output(3, 163) <= input(17);
output(3, 164) <= input(18);
output(3, 165) <= input(19);
output(3, 166) <= input(20);
output(3, 167) <= input(21);
output(3, 168) <= input(22);
output(3, 169) <= input(23);
output(3, 170) <= input(24);
output(3, 171) <= input(25);
output(3, 172) <= input(26);
output(3, 173) <= input(27);
output(3, 174) <= input(28);
output(3, 175) <= input(29);
output(3, 176) <= input(37);
output(3, 177) <= input(35);
output(3, 178) <= input(16);
output(3, 179) <= input(17);
output(3, 180) <= input(18);
output(3, 181) <= input(19);
output(3, 182) <= input(20);
output(3, 183) <= input(21);
output(3, 184) <= input(22);
output(3, 185) <= input(23);
output(3, 186) <= input(24);
output(3, 187) <= input(25);
output(3, 188) <= input(26);
output(3, 189) <= input(27);
output(3, 190) <= input(28);
output(3, 191) <= input(29);
output(3, 192) <= input(37);
output(3, 193) <= input(35);
output(3, 194) <= input(16);
output(3, 195) <= input(17);
output(3, 196) <= input(18);
output(3, 197) <= input(19);
output(3, 198) <= input(20);
output(3, 199) <= input(21);
output(3, 200) <= input(22);
output(3, 201) <= input(23);
output(3, 202) <= input(24);
output(3, 203) <= input(25);
output(3, 204) <= input(26);
output(3, 205) <= input(27);
output(3, 206) <= input(28);
output(3, 207) <= input(29);
output(3, 208) <= input(37);
output(3, 209) <= input(35);
output(3, 210) <= input(16);
output(3, 211) <= input(17);
output(3, 212) <= input(18);
output(3, 213) <= input(19);
output(3, 214) <= input(20);
output(3, 215) <= input(21);
output(3, 216) <= input(22);
output(3, 217) <= input(23);
output(3, 218) <= input(24);
output(3, 219) <= input(25);
output(3, 220) <= input(26);
output(3, 221) <= input(27);
output(3, 222) <= input(28);
output(3, 223) <= input(29);
output(3, 224) <= input(37);
output(3, 225) <= input(35);
output(3, 226) <= input(16);
output(3, 227) <= input(17);
output(3, 228) <= input(18);
output(3, 229) <= input(19);
output(3, 230) <= input(20);
output(3, 231) <= input(21);
output(3, 232) <= input(22);
output(3, 233) <= input(23);
output(3, 234) <= input(24);
output(3, 235) <= input(25);
output(3, 236) <= input(26);
output(3, 237) <= input(27);
output(3, 238) <= input(28);
output(3, 239) <= input(29);
output(3, 240) <= input(36);
output(3, 241) <= input(0);
output(3, 242) <= input(1);
output(3, 243) <= input(2);
output(3, 244) <= input(3);
output(3, 245) <= input(4);
output(3, 246) <= input(5);
output(3, 247) <= input(6);
output(3, 248) <= input(7);
output(3, 249) <= input(8);
output(3, 250) <= input(9);
output(3, 251) <= input(10);
output(3, 252) <= input(11);
output(3, 253) <= input(12);
output(3, 254) <= input(13);
output(3, 255) <= input(14);
output(4, 0) <= input(38);
output(4, 1) <= input(36);
output(4, 2) <= input(0);
output(4, 3) <= input(1);
output(4, 4) <= input(2);
output(4, 5) <= input(3);
output(4, 6) <= input(4);
output(4, 7) <= input(5);
output(4, 8) <= input(6);
output(4, 9) <= input(7);
output(4, 10) <= input(8);
output(4, 11) <= input(9);
output(4, 12) <= input(10);
output(4, 13) <= input(11);
output(4, 14) <= input(12);
output(4, 15) <= input(13);
output(4, 16) <= input(38);
output(4, 17) <= input(36);
output(4, 18) <= input(0);
output(4, 19) <= input(1);
output(4, 20) <= input(2);
output(4, 21) <= input(3);
output(4, 22) <= input(4);
output(4, 23) <= input(5);
output(4, 24) <= input(6);
output(4, 25) <= input(7);
output(4, 26) <= input(8);
output(4, 27) <= input(9);
output(4, 28) <= input(10);
output(4, 29) <= input(11);
output(4, 30) <= input(12);
output(4, 31) <= input(13);
output(4, 32) <= input(38);
output(4, 33) <= input(36);
output(4, 34) <= input(0);
output(4, 35) <= input(1);
output(4, 36) <= input(2);
output(4, 37) <= input(3);
output(4, 38) <= input(4);
output(4, 39) <= input(5);
output(4, 40) <= input(6);
output(4, 41) <= input(7);
output(4, 42) <= input(8);
output(4, 43) <= input(9);
output(4, 44) <= input(10);
output(4, 45) <= input(11);
output(4, 46) <= input(12);
output(4, 47) <= input(13);
output(4, 48) <= input(38);
output(4, 49) <= input(36);
output(4, 50) <= input(0);
output(4, 51) <= input(1);
output(4, 52) <= input(2);
output(4, 53) <= input(3);
output(4, 54) <= input(4);
output(4, 55) <= input(5);
output(4, 56) <= input(6);
output(4, 57) <= input(7);
output(4, 58) <= input(8);
output(4, 59) <= input(9);
output(4, 60) <= input(10);
output(4, 61) <= input(11);
output(4, 62) <= input(12);
output(4, 63) <= input(13);
output(4, 64) <= input(38);
output(4, 65) <= input(36);
output(4, 66) <= input(0);
output(4, 67) <= input(1);
output(4, 68) <= input(2);
output(4, 69) <= input(3);
output(4, 70) <= input(4);
output(4, 71) <= input(5);
output(4, 72) <= input(6);
output(4, 73) <= input(7);
output(4, 74) <= input(8);
output(4, 75) <= input(9);
output(4, 76) <= input(10);
output(4, 77) <= input(11);
output(4, 78) <= input(12);
output(4, 79) <= input(13);
output(4, 80) <= input(38);
output(4, 81) <= input(36);
output(4, 82) <= input(0);
output(4, 83) <= input(1);
output(4, 84) <= input(2);
output(4, 85) <= input(3);
output(4, 86) <= input(4);
output(4, 87) <= input(5);
output(4, 88) <= input(6);
output(4, 89) <= input(7);
output(4, 90) <= input(8);
output(4, 91) <= input(9);
output(4, 92) <= input(10);
output(4, 93) <= input(11);
output(4, 94) <= input(12);
output(4, 95) <= input(13);
output(4, 96) <= input(38);
output(4, 97) <= input(36);
output(4, 98) <= input(0);
output(4, 99) <= input(1);
output(4, 100) <= input(2);
output(4, 101) <= input(3);
output(4, 102) <= input(4);
output(4, 103) <= input(5);
output(4, 104) <= input(6);
output(4, 105) <= input(7);
output(4, 106) <= input(8);
output(4, 107) <= input(9);
output(4, 108) <= input(10);
output(4, 109) <= input(11);
output(4, 110) <= input(12);
output(4, 111) <= input(13);
output(4, 112) <= input(38);
output(4, 113) <= input(36);
output(4, 114) <= input(0);
output(4, 115) <= input(1);
output(4, 116) <= input(2);
output(4, 117) <= input(3);
output(4, 118) <= input(4);
output(4, 119) <= input(5);
output(4, 120) <= input(6);
output(4, 121) <= input(7);
output(4, 122) <= input(8);
output(4, 123) <= input(9);
output(4, 124) <= input(10);
output(4, 125) <= input(11);
output(4, 126) <= input(12);
output(4, 127) <= input(13);
output(4, 128) <= input(38);
output(4, 129) <= input(36);
output(4, 130) <= input(0);
output(4, 131) <= input(1);
output(4, 132) <= input(2);
output(4, 133) <= input(3);
output(4, 134) <= input(4);
output(4, 135) <= input(5);
output(4, 136) <= input(6);
output(4, 137) <= input(7);
output(4, 138) <= input(8);
output(4, 139) <= input(9);
output(4, 140) <= input(10);
output(4, 141) <= input(11);
output(4, 142) <= input(12);
output(4, 143) <= input(13);
output(4, 144) <= input(38);
output(4, 145) <= input(36);
output(4, 146) <= input(0);
output(4, 147) <= input(1);
output(4, 148) <= input(2);
output(4, 149) <= input(3);
output(4, 150) <= input(4);
output(4, 151) <= input(5);
output(4, 152) <= input(6);
output(4, 153) <= input(7);
output(4, 154) <= input(8);
output(4, 155) <= input(9);
output(4, 156) <= input(10);
output(4, 157) <= input(11);
output(4, 158) <= input(12);
output(4, 159) <= input(13);
output(4, 160) <= input(38);
output(4, 161) <= input(36);
output(4, 162) <= input(0);
output(4, 163) <= input(1);
output(4, 164) <= input(2);
output(4, 165) <= input(3);
output(4, 166) <= input(4);
output(4, 167) <= input(5);
output(4, 168) <= input(6);
output(4, 169) <= input(7);
output(4, 170) <= input(8);
output(4, 171) <= input(9);
output(4, 172) <= input(10);
output(4, 173) <= input(11);
output(4, 174) <= input(12);
output(4, 175) <= input(13);
output(4, 176) <= input(38);
output(4, 177) <= input(36);
output(4, 178) <= input(0);
output(4, 179) <= input(1);
output(4, 180) <= input(2);
output(4, 181) <= input(3);
output(4, 182) <= input(4);
output(4, 183) <= input(5);
output(4, 184) <= input(6);
output(4, 185) <= input(7);
output(4, 186) <= input(8);
output(4, 187) <= input(9);
output(4, 188) <= input(10);
output(4, 189) <= input(11);
output(4, 190) <= input(12);
output(4, 191) <= input(13);
output(4, 192) <= input(38);
output(4, 193) <= input(36);
output(4, 194) <= input(0);
output(4, 195) <= input(1);
output(4, 196) <= input(2);
output(4, 197) <= input(3);
output(4, 198) <= input(4);
output(4, 199) <= input(5);
output(4, 200) <= input(6);
output(4, 201) <= input(7);
output(4, 202) <= input(8);
output(4, 203) <= input(9);
output(4, 204) <= input(10);
output(4, 205) <= input(11);
output(4, 206) <= input(12);
output(4, 207) <= input(13);
output(4, 208) <= input(38);
output(4, 209) <= input(36);
output(4, 210) <= input(0);
output(4, 211) <= input(1);
output(4, 212) <= input(2);
output(4, 213) <= input(3);
output(4, 214) <= input(4);
output(4, 215) <= input(5);
output(4, 216) <= input(6);
output(4, 217) <= input(7);
output(4, 218) <= input(8);
output(4, 219) <= input(9);
output(4, 220) <= input(10);
output(4, 221) <= input(11);
output(4, 222) <= input(12);
output(4, 223) <= input(13);
output(4, 224) <= input(38);
output(4, 225) <= input(36);
output(4, 226) <= input(0);
output(4, 227) <= input(1);
output(4, 228) <= input(2);
output(4, 229) <= input(3);
output(4, 230) <= input(4);
output(4, 231) <= input(5);
output(4, 232) <= input(6);
output(4, 233) <= input(7);
output(4, 234) <= input(8);
output(4, 235) <= input(9);
output(4, 236) <= input(10);
output(4, 237) <= input(11);
output(4, 238) <= input(12);
output(4, 239) <= input(13);
output(4, 240) <= input(38);
output(4, 241) <= input(36);
output(4, 242) <= input(0);
output(4, 243) <= input(1);
output(4, 244) <= input(2);
output(4, 245) <= input(3);
output(4, 246) <= input(4);
output(4, 247) <= input(5);
output(4, 248) <= input(6);
output(4, 249) <= input(7);
output(4, 250) <= input(8);
output(4, 251) <= input(9);
output(4, 252) <= input(10);
output(4, 253) <= input(11);
output(4, 254) <= input(12);
output(4, 255) <= input(13);
output(5, 0) <= input(39);
output(5, 1) <= input(38);
output(5, 2) <= input(36);
output(5, 3) <= input(0);
output(5, 4) <= input(1);
output(5, 5) <= input(2);
output(5, 6) <= input(3);
output(5, 7) <= input(4);
output(5, 8) <= input(5);
output(5, 9) <= input(6);
output(5, 10) <= input(7);
output(5, 11) <= input(8);
output(5, 12) <= input(9);
output(5, 13) <= input(10);
output(5, 14) <= input(11);
output(5, 15) <= input(12);
output(5, 16) <= input(39);
output(5, 17) <= input(38);
output(5, 18) <= input(36);
output(5, 19) <= input(0);
output(5, 20) <= input(1);
output(5, 21) <= input(2);
output(5, 22) <= input(3);
output(5, 23) <= input(4);
output(5, 24) <= input(5);
output(5, 25) <= input(6);
output(5, 26) <= input(7);
output(5, 27) <= input(8);
output(5, 28) <= input(9);
output(5, 29) <= input(10);
output(5, 30) <= input(11);
output(5, 31) <= input(12);
output(5, 32) <= input(39);
output(5, 33) <= input(38);
output(5, 34) <= input(36);
output(5, 35) <= input(0);
output(5, 36) <= input(1);
output(5, 37) <= input(2);
output(5, 38) <= input(3);
output(5, 39) <= input(4);
output(5, 40) <= input(5);
output(5, 41) <= input(6);
output(5, 42) <= input(7);
output(5, 43) <= input(8);
output(5, 44) <= input(9);
output(5, 45) <= input(10);
output(5, 46) <= input(11);
output(5, 47) <= input(12);
output(5, 48) <= input(39);
output(5, 49) <= input(38);
output(5, 50) <= input(36);
output(5, 51) <= input(0);
output(5, 52) <= input(1);
output(5, 53) <= input(2);
output(5, 54) <= input(3);
output(5, 55) <= input(4);
output(5, 56) <= input(5);
output(5, 57) <= input(6);
output(5, 58) <= input(7);
output(5, 59) <= input(8);
output(5, 60) <= input(9);
output(5, 61) <= input(10);
output(5, 62) <= input(11);
output(5, 63) <= input(12);
output(5, 64) <= input(39);
output(5, 65) <= input(38);
output(5, 66) <= input(36);
output(5, 67) <= input(0);
output(5, 68) <= input(1);
output(5, 69) <= input(2);
output(5, 70) <= input(3);
output(5, 71) <= input(4);
output(5, 72) <= input(5);
output(5, 73) <= input(6);
output(5, 74) <= input(7);
output(5, 75) <= input(8);
output(5, 76) <= input(9);
output(5, 77) <= input(10);
output(5, 78) <= input(11);
output(5, 79) <= input(12);
output(5, 80) <= input(39);
output(5, 81) <= input(38);
output(5, 82) <= input(36);
output(5, 83) <= input(0);
output(5, 84) <= input(1);
output(5, 85) <= input(2);
output(5, 86) <= input(3);
output(5, 87) <= input(4);
output(5, 88) <= input(5);
output(5, 89) <= input(6);
output(5, 90) <= input(7);
output(5, 91) <= input(8);
output(5, 92) <= input(9);
output(5, 93) <= input(10);
output(5, 94) <= input(11);
output(5, 95) <= input(12);
output(5, 96) <= input(39);
output(5, 97) <= input(38);
output(5, 98) <= input(36);
output(5, 99) <= input(0);
output(5, 100) <= input(1);
output(5, 101) <= input(2);
output(5, 102) <= input(3);
output(5, 103) <= input(4);
output(5, 104) <= input(5);
output(5, 105) <= input(6);
output(5, 106) <= input(7);
output(5, 107) <= input(8);
output(5, 108) <= input(9);
output(5, 109) <= input(10);
output(5, 110) <= input(11);
output(5, 111) <= input(12);
output(5, 112) <= input(39);
output(5, 113) <= input(38);
output(5, 114) <= input(36);
output(5, 115) <= input(0);
output(5, 116) <= input(1);
output(5, 117) <= input(2);
output(5, 118) <= input(3);
output(5, 119) <= input(4);
output(5, 120) <= input(5);
output(5, 121) <= input(6);
output(5, 122) <= input(7);
output(5, 123) <= input(8);
output(5, 124) <= input(9);
output(5, 125) <= input(10);
output(5, 126) <= input(11);
output(5, 127) <= input(12);
output(5, 128) <= input(39);
output(5, 129) <= input(38);
output(5, 130) <= input(36);
output(5, 131) <= input(0);
output(5, 132) <= input(1);
output(5, 133) <= input(2);
output(5, 134) <= input(3);
output(5, 135) <= input(4);
output(5, 136) <= input(5);
output(5, 137) <= input(6);
output(5, 138) <= input(7);
output(5, 139) <= input(8);
output(5, 140) <= input(9);
output(5, 141) <= input(10);
output(5, 142) <= input(11);
output(5, 143) <= input(12);
output(5, 144) <= input(39);
output(5, 145) <= input(38);
output(5, 146) <= input(36);
output(5, 147) <= input(0);
output(5, 148) <= input(1);
output(5, 149) <= input(2);
output(5, 150) <= input(3);
output(5, 151) <= input(4);
output(5, 152) <= input(5);
output(5, 153) <= input(6);
output(5, 154) <= input(7);
output(5, 155) <= input(8);
output(5, 156) <= input(9);
output(5, 157) <= input(10);
output(5, 158) <= input(11);
output(5, 159) <= input(12);
output(5, 160) <= input(39);
output(5, 161) <= input(38);
output(5, 162) <= input(36);
output(5, 163) <= input(0);
output(5, 164) <= input(1);
output(5, 165) <= input(2);
output(5, 166) <= input(3);
output(5, 167) <= input(4);
output(5, 168) <= input(5);
output(5, 169) <= input(6);
output(5, 170) <= input(7);
output(5, 171) <= input(8);
output(5, 172) <= input(9);
output(5, 173) <= input(10);
output(5, 174) <= input(11);
output(5, 175) <= input(12);
output(5, 176) <= input(39);
output(5, 177) <= input(38);
output(5, 178) <= input(36);
output(5, 179) <= input(0);
output(5, 180) <= input(1);
output(5, 181) <= input(2);
output(5, 182) <= input(3);
output(5, 183) <= input(4);
output(5, 184) <= input(5);
output(5, 185) <= input(6);
output(5, 186) <= input(7);
output(5, 187) <= input(8);
output(5, 188) <= input(9);
output(5, 189) <= input(10);
output(5, 190) <= input(11);
output(5, 191) <= input(12);
output(5, 192) <= input(39);
output(5, 193) <= input(38);
output(5, 194) <= input(36);
output(5, 195) <= input(0);
output(5, 196) <= input(1);
output(5, 197) <= input(2);
output(5, 198) <= input(3);
output(5, 199) <= input(4);
output(5, 200) <= input(5);
output(5, 201) <= input(6);
output(5, 202) <= input(7);
output(5, 203) <= input(8);
output(5, 204) <= input(9);
output(5, 205) <= input(10);
output(5, 206) <= input(11);
output(5, 207) <= input(12);
output(5, 208) <= input(39);
output(5, 209) <= input(38);
output(5, 210) <= input(36);
output(5, 211) <= input(0);
output(5, 212) <= input(1);
output(5, 213) <= input(2);
output(5, 214) <= input(3);
output(5, 215) <= input(4);
output(5, 216) <= input(5);
output(5, 217) <= input(6);
output(5, 218) <= input(7);
output(5, 219) <= input(8);
output(5, 220) <= input(9);
output(5, 221) <= input(10);
output(5, 222) <= input(11);
output(5, 223) <= input(12);
output(5, 224) <= input(39);
output(5, 225) <= input(38);
output(5, 226) <= input(36);
output(5, 227) <= input(0);
output(5, 228) <= input(1);
output(5, 229) <= input(2);
output(5, 230) <= input(3);
output(5, 231) <= input(4);
output(5, 232) <= input(5);
output(5, 233) <= input(6);
output(5, 234) <= input(7);
output(5, 235) <= input(8);
output(5, 236) <= input(9);
output(5, 237) <= input(10);
output(5, 238) <= input(11);
output(5, 239) <= input(12);
output(5, 240) <= input(39);
output(5, 241) <= input(38);
output(5, 242) <= input(36);
output(5, 243) <= input(0);
output(5, 244) <= input(1);
output(5, 245) <= input(2);
output(5, 246) <= input(3);
output(5, 247) <= input(4);
output(5, 248) <= input(5);
output(5, 249) <= input(6);
output(5, 250) <= input(7);
output(5, 251) <= input(8);
output(5, 252) <= input(9);
output(5, 253) <= input(10);
output(5, 254) <= input(11);
output(5, 255) <= input(12);
output(6, 0) <= input(40);
output(6, 1) <= input(41);
output(6, 2) <= input(37);
output(6, 3) <= input(35);
output(6, 4) <= input(16);
output(6, 5) <= input(17);
output(6, 6) <= input(18);
output(6, 7) <= input(19);
output(6, 8) <= input(20);
output(6, 9) <= input(21);
output(6, 10) <= input(22);
output(6, 11) <= input(23);
output(6, 12) <= input(24);
output(6, 13) <= input(25);
output(6, 14) <= input(26);
output(6, 15) <= input(27);
output(6, 16) <= input(40);
output(6, 17) <= input(41);
output(6, 18) <= input(37);
output(6, 19) <= input(35);
output(6, 20) <= input(16);
output(6, 21) <= input(17);
output(6, 22) <= input(18);
output(6, 23) <= input(19);
output(6, 24) <= input(20);
output(6, 25) <= input(21);
output(6, 26) <= input(22);
output(6, 27) <= input(23);
output(6, 28) <= input(24);
output(6, 29) <= input(25);
output(6, 30) <= input(26);
output(6, 31) <= input(27);
output(6, 32) <= input(40);
output(6, 33) <= input(41);
output(6, 34) <= input(37);
output(6, 35) <= input(35);
output(6, 36) <= input(16);
output(6, 37) <= input(17);
output(6, 38) <= input(18);
output(6, 39) <= input(19);
output(6, 40) <= input(20);
output(6, 41) <= input(21);
output(6, 42) <= input(22);
output(6, 43) <= input(23);
output(6, 44) <= input(24);
output(6, 45) <= input(25);
output(6, 46) <= input(26);
output(6, 47) <= input(27);
output(6, 48) <= input(40);
output(6, 49) <= input(41);
output(6, 50) <= input(37);
output(6, 51) <= input(35);
output(6, 52) <= input(16);
output(6, 53) <= input(17);
output(6, 54) <= input(18);
output(6, 55) <= input(19);
output(6, 56) <= input(20);
output(6, 57) <= input(21);
output(6, 58) <= input(22);
output(6, 59) <= input(23);
output(6, 60) <= input(24);
output(6, 61) <= input(25);
output(6, 62) <= input(26);
output(6, 63) <= input(27);
output(6, 64) <= input(40);
output(6, 65) <= input(41);
output(6, 66) <= input(37);
output(6, 67) <= input(35);
output(6, 68) <= input(16);
output(6, 69) <= input(17);
output(6, 70) <= input(18);
output(6, 71) <= input(19);
output(6, 72) <= input(20);
output(6, 73) <= input(21);
output(6, 74) <= input(22);
output(6, 75) <= input(23);
output(6, 76) <= input(24);
output(6, 77) <= input(25);
output(6, 78) <= input(26);
output(6, 79) <= input(27);
output(6, 80) <= input(40);
output(6, 81) <= input(41);
output(6, 82) <= input(37);
output(6, 83) <= input(35);
output(6, 84) <= input(16);
output(6, 85) <= input(17);
output(6, 86) <= input(18);
output(6, 87) <= input(19);
output(6, 88) <= input(20);
output(6, 89) <= input(21);
output(6, 90) <= input(22);
output(6, 91) <= input(23);
output(6, 92) <= input(24);
output(6, 93) <= input(25);
output(6, 94) <= input(26);
output(6, 95) <= input(27);
output(6, 96) <= input(40);
output(6, 97) <= input(41);
output(6, 98) <= input(37);
output(6, 99) <= input(35);
output(6, 100) <= input(16);
output(6, 101) <= input(17);
output(6, 102) <= input(18);
output(6, 103) <= input(19);
output(6, 104) <= input(20);
output(6, 105) <= input(21);
output(6, 106) <= input(22);
output(6, 107) <= input(23);
output(6, 108) <= input(24);
output(6, 109) <= input(25);
output(6, 110) <= input(26);
output(6, 111) <= input(27);
output(6, 112) <= input(40);
output(6, 113) <= input(41);
output(6, 114) <= input(37);
output(6, 115) <= input(35);
output(6, 116) <= input(16);
output(6, 117) <= input(17);
output(6, 118) <= input(18);
output(6, 119) <= input(19);
output(6, 120) <= input(20);
output(6, 121) <= input(21);
output(6, 122) <= input(22);
output(6, 123) <= input(23);
output(6, 124) <= input(24);
output(6, 125) <= input(25);
output(6, 126) <= input(26);
output(6, 127) <= input(27);
output(6, 128) <= input(42);
output(6, 129) <= input(43);
output(6, 130) <= input(38);
output(6, 131) <= input(36);
output(6, 132) <= input(0);
output(6, 133) <= input(1);
output(6, 134) <= input(2);
output(6, 135) <= input(3);
output(6, 136) <= input(4);
output(6, 137) <= input(5);
output(6, 138) <= input(6);
output(6, 139) <= input(7);
output(6, 140) <= input(8);
output(6, 141) <= input(9);
output(6, 142) <= input(10);
output(6, 143) <= input(11);
output(6, 144) <= input(42);
output(6, 145) <= input(43);
output(6, 146) <= input(38);
output(6, 147) <= input(36);
output(6, 148) <= input(0);
output(6, 149) <= input(1);
output(6, 150) <= input(2);
output(6, 151) <= input(3);
output(6, 152) <= input(4);
output(6, 153) <= input(5);
output(6, 154) <= input(6);
output(6, 155) <= input(7);
output(6, 156) <= input(8);
output(6, 157) <= input(9);
output(6, 158) <= input(10);
output(6, 159) <= input(11);
output(6, 160) <= input(42);
output(6, 161) <= input(43);
output(6, 162) <= input(38);
output(6, 163) <= input(36);
output(6, 164) <= input(0);
output(6, 165) <= input(1);
output(6, 166) <= input(2);
output(6, 167) <= input(3);
output(6, 168) <= input(4);
output(6, 169) <= input(5);
output(6, 170) <= input(6);
output(6, 171) <= input(7);
output(6, 172) <= input(8);
output(6, 173) <= input(9);
output(6, 174) <= input(10);
output(6, 175) <= input(11);
output(6, 176) <= input(42);
output(6, 177) <= input(43);
output(6, 178) <= input(38);
output(6, 179) <= input(36);
output(6, 180) <= input(0);
output(6, 181) <= input(1);
output(6, 182) <= input(2);
output(6, 183) <= input(3);
output(6, 184) <= input(4);
output(6, 185) <= input(5);
output(6, 186) <= input(6);
output(6, 187) <= input(7);
output(6, 188) <= input(8);
output(6, 189) <= input(9);
output(6, 190) <= input(10);
output(6, 191) <= input(11);
output(6, 192) <= input(42);
output(6, 193) <= input(43);
output(6, 194) <= input(38);
output(6, 195) <= input(36);
output(6, 196) <= input(0);
output(6, 197) <= input(1);
output(6, 198) <= input(2);
output(6, 199) <= input(3);
output(6, 200) <= input(4);
output(6, 201) <= input(5);
output(6, 202) <= input(6);
output(6, 203) <= input(7);
output(6, 204) <= input(8);
output(6, 205) <= input(9);
output(6, 206) <= input(10);
output(6, 207) <= input(11);
output(6, 208) <= input(42);
output(6, 209) <= input(43);
output(6, 210) <= input(38);
output(6, 211) <= input(36);
output(6, 212) <= input(0);
output(6, 213) <= input(1);
output(6, 214) <= input(2);
output(6, 215) <= input(3);
output(6, 216) <= input(4);
output(6, 217) <= input(5);
output(6, 218) <= input(6);
output(6, 219) <= input(7);
output(6, 220) <= input(8);
output(6, 221) <= input(9);
output(6, 222) <= input(10);
output(6, 223) <= input(11);
output(6, 224) <= input(42);
output(6, 225) <= input(43);
output(6, 226) <= input(38);
output(6, 227) <= input(36);
output(6, 228) <= input(0);
output(6, 229) <= input(1);
output(6, 230) <= input(2);
output(6, 231) <= input(3);
output(6, 232) <= input(4);
output(6, 233) <= input(5);
output(6, 234) <= input(6);
output(6, 235) <= input(7);
output(6, 236) <= input(8);
output(6, 237) <= input(9);
output(6, 238) <= input(10);
output(6, 239) <= input(11);
output(6, 240) <= input(42);
output(6, 241) <= input(43);
output(6, 242) <= input(38);
output(6, 243) <= input(36);
output(6, 244) <= input(0);
output(6, 245) <= input(1);
output(6, 246) <= input(2);
output(6, 247) <= input(3);
output(6, 248) <= input(4);
output(6, 249) <= input(5);
output(6, 250) <= input(6);
output(6, 251) <= input(7);
output(6, 252) <= input(8);
output(6, 253) <= input(9);
output(6, 254) <= input(10);
output(6, 255) <= input(11);
output(7, 0) <= input(44);
output(7, 1) <= input(45);
output(7, 2) <= input(38);
output(7, 3) <= input(36);
output(7, 4) <= input(0);
output(7, 5) <= input(1);
output(7, 6) <= input(2);
output(7, 7) <= input(3);
output(7, 8) <= input(4);
output(7, 9) <= input(5);
output(7, 10) <= input(6);
output(7, 11) <= input(7);
output(7, 12) <= input(8);
output(7, 13) <= input(9);
output(7, 14) <= input(10);
output(7, 15) <= input(11);
output(7, 16) <= input(44);
output(7, 17) <= input(45);
output(7, 18) <= input(38);
output(7, 19) <= input(36);
output(7, 20) <= input(0);
output(7, 21) <= input(1);
output(7, 22) <= input(2);
output(7, 23) <= input(3);
output(7, 24) <= input(4);
output(7, 25) <= input(5);
output(7, 26) <= input(6);
output(7, 27) <= input(7);
output(7, 28) <= input(8);
output(7, 29) <= input(9);
output(7, 30) <= input(10);
output(7, 31) <= input(11);
output(7, 32) <= input(44);
output(7, 33) <= input(45);
output(7, 34) <= input(38);
output(7, 35) <= input(36);
output(7, 36) <= input(0);
output(7, 37) <= input(1);
output(7, 38) <= input(2);
output(7, 39) <= input(3);
output(7, 40) <= input(4);
output(7, 41) <= input(5);
output(7, 42) <= input(6);
output(7, 43) <= input(7);
output(7, 44) <= input(8);
output(7, 45) <= input(9);
output(7, 46) <= input(10);
output(7, 47) <= input(11);
output(7, 48) <= input(44);
output(7, 49) <= input(45);
output(7, 50) <= input(38);
output(7, 51) <= input(36);
output(7, 52) <= input(0);
output(7, 53) <= input(1);
output(7, 54) <= input(2);
output(7, 55) <= input(3);
output(7, 56) <= input(4);
output(7, 57) <= input(5);
output(7, 58) <= input(6);
output(7, 59) <= input(7);
output(7, 60) <= input(8);
output(7, 61) <= input(9);
output(7, 62) <= input(10);
output(7, 63) <= input(11);
output(7, 64) <= input(44);
output(7, 65) <= input(45);
output(7, 66) <= input(38);
output(7, 67) <= input(36);
output(7, 68) <= input(0);
output(7, 69) <= input(1);
output(7, 70) <= input(2);
output(7, 71) <= input(3);
output(7, 72) <= input(4);
output(7, 73) <= input(5);
output(7, 74) <= input(6);
output(7, 75) <= input(7);
output(7, 76) <= input(8);
output(7, 77) <= input(9);
output(7, 78) <= input(10);
output(7, 79) <= input(11);
output(7, 80) <= input(46);
output(7, 81) <= input(47);
output(7, 82) <= input(48);
output(7, 83) <= input(37);
output(7, 84) <= input(35);
output(7, 85) <= input(16);
output(7, 86) <= input(17);
output(7, 87) <= input(18);
output(7, 88) <= input(19);
output(7, 89) <= input(20);
output(7, 90) <= input(21);
output(7, 91) <= input(22);
output(7, 92) <= input(23);
output(7, 93) <= input(24);
output(7, 94) <= input(25);
output(7, 95) <= input(26);
output(7, 96) <= input(46);
output(7, 97) <= input(47);
output(7, 98) <= input(48);
output(7, 99) <= input(37);
output(7, 100) <= input(35);
output(7, 101) <= input(16);
output(7, 102) <= input(17);
output(7, 103) <= input(18);
output(7, 104) <= input(19);
output(7, 105) <= input(20);
output(7, 106) <= input(21);
output(7, 107) <= input(22);
output(7, 108) <= input(23);
output(7, 109) <= input(24);
output(7, 110) <= input(25);
output(7, 111) <= input(26);
output(7, 112) <= input(46);
output(7, 113) <= input(47);
output(7, 114) <= input(48);
output(7, 115) <= input(37);
output(7, 116) <= input(35);
output(7, 117) <= input(16);
output(7, 118) <= input(17);
output(7, 119) <= input(18);
output(7, 120) <= input(19);
output(7, 121) <= input(20);
output(7, 122) <= input(21);
output(7, 123) <= input(22);
output(7, 124) <= input(23);
output(7, 125) <= input(24);
output(7, 126) <= input(25);
output(7, 127) <= input(26);
output(7, 128) <= input(46);
output(7, 129) <= input(47);
output(7, 130) <= input(48);
output(7, 131) <= input(37);
output(7, 132) <= input(35);
output(7, 133) <= input(16);
output(7, 134) <= input(17);
output(7, 135) <= input(18);
output(7, 136) <= input(19);
output(7, 137) <= input(20);
output(7, 138) <= input(21);
output(7, 139) <= input(22);
output(7, 140) <= input(23);
output(7, 141) <= input(24);
output(7, 142) <= input(25);
output(7, 143) <= input(26);
output(7, 144) <= input(46);
output(7, 145) <= input(47);
output(7, 146) <= input(48);
output(7, 147) <= input(37);
output(7, 148) <= input(35);
output(7, 149) <= input(16);
output(7, 150) <= input(17);
output(7, 151) <= input(18);
output(7, 152) <= input(19);
output(7, 153) <= input(20);
output(7, 154) <= input(21);
output(7, 155) <= input(22);
output(7, 156) <= input(23);
output(7, 157) <= input(24);
output(7, 158) <= input(25);
output(7, 159) <= input(26);
output(7, 160) <= input(49);
output(7, 161) <= input(44);
output(7, 162) <= input(45);
output(7, 163) <= input(38);
output(7, 164) <= input(36);
output(7, 165) <= input(0);
output(7, 166) <= input(1);
output(7, 167) <= input(2);
output(7, 168) <= input(3);
output(7, 169) <= input(4);
output(7, 170) <= input(5);
output(7, 171) <= input(6);
output(7, 172) <= input(7);
output(7, 173) <= input(8);
output(7, 174) <= input(9);
output(7, 175) <= input(10);
output(7, 176) <= input(49);
output(7, 177) <= input(44);
output(7, 178) <= input(45);
output(7, 179) <= input(38);
output(7, 180) <= input(36);
output(7, 181) <= input(0);
output(7, 182) <= input(1);
output(7, 183) <= input(2);
output(7, 184) <= input(3);
output(7, 185) <= input(4);
output(7, 186) <= input(5);
output(7, 187) <= input(6);
output(7, 188) <= input(7);
output(7, 189) <= input(8);
output(7, 190) <= input(9);
output(7, 191) <= input(10);
output(7, 192) <= input(49);
output(7, 193) <= input(44);
output(7, 194) <= input(45);
output(7, 195) <= input(38);
output(7, 196) <= input(36);
output(7, 197) <= input(0);
output(7, 198) <= input(1);
output(7, 199) <= input(2);
output(7, 200) <= input(3);
output(7, 201) <= input(4);
output(7, 202) <= input(5);
output(7, 203) <= input(6);
output(7, 204) <= input(7);
output(7, 205) <= input(8);
output(7, 206) <= input(9);
output(7, 207) <= input(10);
output(7, 208) <= input(49);
output(7, 209) <= input(44);
output(7, 210) <= input(45);
output(7, 211) <= input(38);
output(7, 212) <= input(36);
output(7, 213) <= input(0);
output(7, 214) <= input(1);
output(7, 215) <= input(2);
output(7, 216) <= input(3);
output(7, 217) <= input(4);
output(7, 218) <= input(5);
output(7, 219) <= input(6);
output(7, 220) <= input(7);
output(7, 221) <= input(8);
output(7, 222) <= input(9);
output(7, 223) <= input(10);
output(7, 224) <= input(49);
output(7, 225) <= input(44);
output(7, 226) <= input(45);
output(7, 227) <= input(38);
output(7, 228) <= input(36);
output(7, 229) <= input(0);
output(7, 230) <= input(1);
output(7, 231) <= input(2);
output(7, 232) <= input(3);
output(7, 233) <= input(4);
output(7, 234) <= input(5);
output(7, 235) <= input(6);
output(7, 236) <= input(7);
output(7, 237) <= input(8);
output(7, 238) <= input(9);
output(7, 239) <= input(10);
output(7, 240) <= input(49);
output(7, 241) <= input(44);
output(7, 242) <= input(45);
output(7, 243) <= input(38);
output(7, 244) <= input(36);
output(7, 245) <= input(0);
output(7, 246) <= input(1);
output(7, 247) <= input(2);
output(7, 248) <= input(3);
output(7, 249) <= input(4);
output(7, 250) <= input(5);
output(7, 251) <= input(6);
output(7, 252) <= input(7);
output(7, 253) <= input(8);
output(7, 254) <= input(9);
output(7, 255) <= input(10);
when "0011" =>
output(0, 0) <= input(0);
output(0, 1) <= input(1);
output(0, 2) <= input(2);
output(0, 3) <= input(3);
output(0, 4) <= input(4);
output(0, 5) <= input(5);
output(0, 6) <= input(6);
output(0, 7) <= input(7);
output(0, 8) <= input(8);
output(0, 9) <= input(9);
output(0, 10) <= input(10);
output(0, 11) <= input(11);
output(0, 12) <= input(12);
output(0, 13) <= input(13);
output(0, 14) <= input(14);
output(0, 15) <= input(15);
output(0, 16) <= input(0);
output(0, 17) <= input(1);
output(0, 18) <= input(2);
output(0, 19) <= input(3);
output(0, 20) <= input(4);
output(0, 21) <= input(5);
output(0, 22) <= input(6);
output(0, 23) <= input(7);
output(0, 24) <= input(8);
output(0, 25) <= input(9);
output(0, 26) <= input(10);
output(0, 27) <= input(11);
output(0, 28) <= input(12);
output(0, 29) <= input(13);
output(0, 30) <= input(14);
output(0, 31) <= input(15);
output(0, 32) <= input(0);
output(0, 33) <= input(1);
output(0, 34) <= input(2);
output(0, 35) <= input(3);
output(0, 36) <= input(4);
output(0, 37) <= input(5);
output(0, 38) <= input(6);
output(0, 39) <= input(7);
output(0, 40) <= input(8);
output(0, 41) <= input(9);
output(0, 42) <= input(10);
output(0, 43) <= input(11);
output(0, 44) <= input(12);
output(0, 45) <= input(13);
output(0, 46) <= input(14);
output(0, 47) <= input(15);
output(0, 48) <= input(0);
output(0, 49) <= input(1);
output(0, 50) <= input(2);
output(0, 51) <= input(3);
output(0, 52) <= input(4);
output(0, 53) <= input(5);
output(0, 54) <= input(6);
output(0, 55) <= input(7);
output(0, 56) <= input(8);
output(0, 57) <= input(9);
output(0, 58) <= input(10);
output(0, 59) <= input(11);
output(0, 60) <= input(12);
output(0, 61) <= input(13);
output(0, 62) <= input(14);
output(0, 63) <= input(15);
output(0, 64) <= input(16);
output(0, 65) <= input(17);
output(0, 66) <= input(18);
output(0, 67) <= input(19);
output(0, 68) <= input(20);
output(0, 69) <= input(21);
output(0, 70) <= input(22);
output(0, 71) <= input(23);
output(0, 72) <= input(24);
output(0, 73) <= input(25);
output(0, 74) <= input(26);
output(0, 75) <= input(27);
output(0, 76) <= input(28);
output(0, 77) <= input(29);
output(0, 78) <= input(30);
output(0, 79) <= input(31);
output(0, 80) <= input(16);
output(0, 81) <= input(17);
output(0, 82) <= input(18);
output(0, 83) <= input(19);
output(0, 84) <= input(20);
output(0, 85) <= input(21);
output(0, 86) <= input(22);
output(0, 87) <= input(23);
output(0, 88) <= input(24);
output(0, 89) <= input(25);
output(0, 90) <= input(26);
output(0, 91) <= input(27);
output(0, 92) <= input(28);
output(0, 93) <= input(29);
output(0, 94) <= input(30);
output(0, 95) <= input(31);
output(0, 96) <= input(16);
output(0, 97) <= input(17);
output(0, 98) <= input(18);
output(0, 99) <= input(19);
output(0, 100) <= input(20);
output(0, 101) <= input(21);
output(0, 102) <= input(22);
output(0, 103) <= input(23);
output(0, 104) <= input(24);
output(0, 105) <= input(25);
output(0, 106) <= input(26);
output(0, 107) <= input(27);
output(0, 108) <= input(28);
output(0, 109) <= input(29);
output(0, 110) <= input(30);
output(0, 111) <= input(31);
output(0, 112) <= input(16);
output(0, 113) <= input(17);
output(0, 114) <= input(18);
output(0, 115) <= input(19);
output(0, 116) <= input(20);
output(0, 117) <= input(21);
output(0, 118) <= input(22);
output(0, 119) <= input(23);
output(0, 120) <= input(24);
output(0, 121) <= input(25);
output(0, 122) <= input(26);
output(0, 123) <= input(27);
output(0, 124) <= input(28);
output(0, 125) <= input(29);
output(0, 126) <= input(30);
output(0, 127) <= input(31);
output(0, 128) <= input(32);
output(0, 129) <= input(0);
output(0, 130) <= input(1);
output(0, 131) <= input(2);
output(0, 132) <= input(3);
output(0, 133) <= input(4);
output(0, 134) <= input(5);
output(0, 135) <= input(6);
output(0, 136) <= input(7);
output(0, 137) <= input(8);
output(0, 138) <= input(9);
output(0, 139) <= input(10);
output(0, 140) <= input(11);
output(0, 141) <= input(12);
output(0, 142) <= input(13);
output(0, 143) <= input(14);
output(0, 144) <= input(32);
output(0, 145) <= input(0);
output(0, 146) <= input(1);
output(0, 147) <= input(2);
output(0, 148) <= input(3);
output(0, 149) <= input(4);
output(0, 150) <= input(5);
output(0, 151) <= input(6);
output(0, 152) <= input(7);
output(0, 153) <= input(8);
output(0, 154) <= input(9);
output(0, 155) <= input(10);
output(0, 156) <= input(11);
output(0, 157) <= input(12);
output(0, 158) <= input(13);
output(0, 159) <= input(14);
output(0, 160) <= input(32);
output(0, 161) <= input(0);
output(0, 162) <= input(1);
output(0, 163) <= input(2);
output(0, 164) <= input(3);
output(0, 165) <= input(4);
output(0, 166) <= input(5);
output(0, 167) <= input(6);
output(0, 168) <= input(7);
output(0, 169) <= input(8);
output(0, 170) <= input(9);
output(0, 171) <= input(10);
output(0, 172) <= input(11);
output(0, 173) <= input(12);
output(0, 174) <= input(13);
output(0, 175) <= input(14);
output(0, 176) <= input(32);
output(0, 177) <= input(0);
output(0, 178) <= input(1);
output(0, 179) <= input(2);
output(0, 180) <= input(3);
output(0, 181) <= input(4);
output(0, 182) <= input(5);
output(0, 183) <= input(6);
output(0, 184) <= input(7);
output(0, 185) <= input(8);
output(0, 186) <= input(9);
output(0, 187) <= input(10);
output(0, 188) <= input(11);
output(0, 189) <= input(12);
output(0, 190) <= input(13);
output(0, 191) <= input(14);
output(0, 192) <= input(33);
output(0, 193) <= input(16);
output(0, 194) <= input(17);
output(0, 195) <= input(18);
output(0, 196) <= input(19);
output(0, 197) <= input(20);
output(0, 198) <= input(21);
output(0, 199) <= input(22);
output(0, 200) <= input(23);
output(0, 201) <= input(24);
output(0, 202) <= input(25);
output(0, 203) <= input(26);
output(0, 204) <= input(27);
output(0, 205) <= input(28);
output(0, 206) <= input(29);
output(0, 207) <= input(30);
output(0, 208) <= input(33);
output(0, 209) <= input(16);
output(0, 210) <= input(17);
output(0, 211) <= input(18);
output(0, 212) <= input(19);
output(0, 213) <= input(20);
output(0, 214) <= input(21);
output(0, 215) <= input(22);
output(0, 216) <= input(23);
output(0, 217) <= input(24);
output(0, 218) <= input(25);
output(0, 219) <= input(26);
output(0, 220) <= input(27);
output(0, 221) <= input(28);
output(0, 222) <= input(29);
output(0, 223) <= input(30);
output(0, 224) <= input(33);
output(0, 225) <= input(16);
output(0, 226) <= input(17);
output(0, 227) <= input(18);
output(0, 228) <= input(19);
output(0, 229) <= input(20);
output(0, 230) <= input(21);
output(0, 231) <= input(22);
output(0, 232) <= input(23);
output(0, 233) <= input(24);
output(0, 234) <= input(25);
output(0, 235) <= input(26);
output(0, 236) <= input(27);
output(0, 237) <= input(28);
output(0, 238) <= input(29);
output(0, 239) <= input(30);
output(0, 240) <= input(33);
output(0, 241) <= input(16);
output(0, 242) <= input(17);
output(0, 243) <= input(18);
output(0, 244) <= input(19);
output(0, 245) <= input(20);
output(0, 246) <= input(21);
output(0, 247) <= input(22);
output(0, 248) <= input(23);
output(0, 249) <= input(24);
output(0, 250) <= input(25);
output(0, 251) <= input(26);
output(0, 252) <= input(27);
output(0, 253) <= input(28);
output(0, 254) <= input(29);
output(0, 255) <= input(30);
output(1, 0) <= input(34);
output(1, 1) <= input(35);
output(1, 2) <= input(36);
output(1, 3) <= input(37);
output(1, 4) <= input(3);
output(1, 5) <= input(4);
output(1, 6) <= input(5);
output(1, 7) <= input(6);
output(1, 8) <= input(7);
output(1, 9) <= input(8);
output(1, 10) <= input(9);
output(1, 11) <= input(10);
output(1, 12) <= input(11);
output(1, 13) <= input(12);
output(1, 14) <= input(13);
output(1, 15) <= input(14);
output(1, 16) <= input(34);
output(1, 17) <= input(35);
output(1, 18) <= input(36);
output(1, 19) <= input(37);
output(1, 20) <= input(3);
output(1, 21) <= input(4);
output(1, 22) <= input(5);
output(1, 23) <= input(6);
output(1, 24) <= input(7);
output(1, 25) <= input(8);
output(1, 26) <= input(9);
output(1, 27) <= input(10);
output(1, 28) <= input(11);
output(1, 29) <= input(12);
output(1, 30) <= input(13);
output(1, 31) <= input(14);
output(1, 32) <= input(38);
output(1, 33) <= input(39);
output(1, 34) <= input(40);
output(1, 35) <= input(41);
output(1, 36) <= input(19);
output(1, 37) <= input(20);
output(1, 38) <= input(21);
output(1, 39) <= input(22);
output(1, 40) <= input(23);
output(1, 41) <= input(24);
output(1, 42) <= input(25);
output(1, 43) <= input(26);
output(1, 44) <= input(27);
output(1, 45) <= input(28);
output(1, 46) <= input(29);
output(1, 47) <= input(30);
output(1, 48) <= input(38);
output(1, 49) <= input(39);
output(1, 50) <= input(40);
output(1, 51) <= input(41);
output(1, 52) <= input(19);
output(1, 53) <= input(20);
output(1, 54) <= input(21);
output(1, 55) <= input(22);
output(1, 56) <= input(23);
output(1, 57) <= input(24);
output(1, 58) <= input(25);
output(1, 59) <= input(26);
output(1, 60) <= input(27);
output(1, 61) <= input(28);
output(1, 62) <= input(29);
output(1, 63) <= input(30);
output(1, 64) <= input(38);
output(1, 65) <= input(39);
output(1, 66) <= input(40);
output(1, 67) <= input(41);
output(1, 68) <= input(19);
output(1, 69) <= input(20);
output(1, 70) <= input(21);
output(1, 71) <= input(22);
output(1, 72) <= input(23);
output(1, 73) <= input(24);
output(1, 74) <= input(25);
output(1, 75) <= input(26);
output(1, 76) <= input(27);
output(1, 77) <= input(28);
output(1, 78) <= input(29);
output(1, 79) <= input(30);
output(1, 80) <= input(42);
output(1, 81) <= input(34);
output(1, 82) <= input(35);
output(1, 83) <= input(36);
output(1, 84) <= input(37);
output(1, 85) <= input(3);
output(1, 86) <= input(4);
output(1, 87) <= input(5);
output(1, 88) <= input(6);
output(1, 89) <= input(7);
output(1, 90) <= input(8);
output(1, 91) <= input(9);
output(1, 92) <= input(10);
output(1, 93) <= input(11);
output(1, 94) <= input(12);
output(1, 95) <= input(13);
output(1, 96) <= input(42);
output(1, 97) <= input(34);
output(1, 98) <= input(35);
output(1, 99) <= input(36);
output(1, 100) <= input(37);
output(1, 101) <= input(3);
output(1, 102) <= input(4);
output(1, 103) <= input(5);
output(1, 104) <= input(6);
output(1, 105) <= input(7);
output(1, 106) <= input(8);
output(1, 107) <= input(9);
output(1, 108) <= input(10);
output(1, 109) <= input(11);
output(1, 110) <= input(12);
output(1, 111) <= input(13);
output(1, 112) <= input(42);
output(1, 113) <= input(34);
output(1, 114) <= input(35);
output(1, 115) <= input(36);
output(1, 116) <= input(37);
output(1, 117) <= input(3);
output(1, 118) <= input(4);
output(1, 119) <= input(5);
output(1, 120) <= input(6);
output(1, 121) <= input(7);
output(1, 122) <= input(8);
output(1, 123) <= input(9);
output(1, 124) <= input(10);
output(1, 125) <= input(11);
output(1, 126) <= input(12);
output(1, 127) <= input(13);
output(1, 128) <= input(43);
output(1, 129) <= input(38);
output(1, 130) <= input(39);
output(1, 131) <= input(40);
output(1, 132) <= input(41);
output(1, 133) <= input(19);
output(1, 134) <= input(20);
output(1, 135) <= input(21);
output(1, 136) <= input(22);
output(1, 137) <= input(23);
output(1, 138) <= input(24);
output(1, 139) <= input(25);
output(1, 140) <= input(26);
output(1, 141) <= input(27);
output(1, 142) <= input(28);
output(1, 143) <= input(29);
output(1, 144) <= input(43);
output(1, 145) <= input(38);
output(1, 146) <= input(39);
output(1, 147) <= input(40);
output(1, 148) <= input(41);
output(1, 149) <= input(19);
output(1, 150) <= input(20);
output(1, 151) <= input(21);
output(1, 152) <= input(22);
output(1, 153) <= input(23);
output(1, 154) <= input(24);
output(1, 155) <= input(25);
output(1, 156) <= input(26);
output(1, 157) <= input(27);
output(1, 158) <= input(28);
output(1, 159) <= input(29);
output(1, 160) <= input(44);
output(1, 161) <= input(42);
output(1, 162) <= input(34);
output(1, 163) <= input(35);
output(1, 164) <= input(36);
output(1, 165) <= input(37);
output(1, 166) <= input(3);
output(1, 167) <= input(4);
output(1, 168) <= input(5);
output(1, 169) <= input(6);
output(1, 170) <= input(7);
output(1, 171) <= input(8);
output(1, 172) <= input(9);
output(1, 173) <= input(10);
output(1, 174) <= input(11);
output(1, 175) <= input(12);
output(1, 176) <= input(44);
output(1, 177) <= input(42);
output(1, 178) <= input(34);
output(1, 179) <= input(35);
output(1, 180) <= input(36);
output(1, 181) <= input(37);
output(1, 182) <= input(3);
output(1, 183) <= input(4);
output(1, 184) <= input(5);
output(1, 185) <= input(6);
output(1, 186) <= input(7);
output(1, 187) <= input(8);
output(1, 188) <= input(9);
output(1, 189) <= input(10);
output(1, 190) <= input(11);
output(1, 191) <= input(12);
output(1, 192) <= input(44);
output(1, 193) <= input(42);
output(1, 194) <= input(34);
output(1, 195) <= input(35);
output(1, 196) <= input(36);
output(1, 197) <= input(37);
output(1, 198) <= input(3);
output(1, 199) <= input(4);
output(1, 200) <= input(5);
output(1, 201) <= input(6);
output(1, 202) <= input(7);
output(1, 203) <= input(8);
output(1, 204) <= input(9);
output(1, 205) <= input(10);
output(1, 206) <= input(11);
output(1, 207) <= input(12);
output(1, 208) <= input(45);
output(1, 209) <= input(43);
output(1, 210) <= input(38);
output(1, 211) <= input(39);
output(1, 212) <= input(40);
output(1, 213) <= input(41);
output(1, 214) <= input(19);
output(1, 215) <= input(20);
output(1, 216) <= input(21);
output(1, 217) <= input(22);
output(1, 218) <= input(23);
output(1, 219) <= input(24);
output(1, 220) <= input(25);
output(1, 221) <= input(26);
output(1, 222) <= input(27);
output(1, 223) <= input(28);
output(1, 224) <= input(45);
output(1, 225) <= input(43);
output(1, 226) <= input(38);
output(1, 227) <= input(39);
output(1, 228) <= input(40);
output(1, 229) <= input(41);
output(1, 230) <= input(19);
output(1, 231) <= input(20);
output(1, 232) <= input(21);
output(1, 233) <= input(22);
output(1, 234) <= input(23);
output(1, 235) <= input(24);
output(1, 236) <= input(25);
output(1, 237) <= input(26);
output(1, 238) <= input(27);
output(1, 239) <= input(28);
output(1, 240) <= input(45);
output(1, 241) <= input(43);
output(1, 242) <= input(38);
output(1, 243) <= input(39);
output(1, 244) <= input(40);
output(1, 245) <= input(41);
output(1, 246) <= input(19);
output(1, 247) <= input(20);
output(1, 248) <= input(21);
output(1, 249) <= input(22);
output(1, 250) <= input(23);
output(1, 251) <= input(24);
output(1, 252) <= input(25);
output(1, 253) <= input(26);
output(1, 254) <= input(27);
output(1, 255) <= input(28);
output(2, 0) <= input(46);
output(2, 1) <= input(47);
output(2, 2) <= input(48);
output(2, 3) <= input(49);
output(2, 4) <= input(50);
output(2, 5) <= input(3);
output(2, 6) <= input(4);
output(2, 7) <= input(5);
output(2, 8) <= input(6);
output(2, 9) <= input(7);
output(2, 10) <= input(8);
output(2, 11) <= input(9);
output(2, 12) <= input(10);
output(2, 13) <= input(11);
output(2, 14) <= input(12);
output(2, 15) <= input(13);
output(2, 16) <= input(46);
output(2, 17) <= input(47);
output(2, 18) <= input(48);
output(2, 19) <= input(49);
output(2, 20) <= input(50);
output(2, 21) <= input(3);
output(2, 22) <= input(4);
output(2, 23) <= input(5);
output(2, 24) <= input(6);
output(2, 25) <= input(7);
output(2, 26) <= input(8);
output(2, 27) <= input(9);
output(2, 28) <= input(10);
output(2, 29) <= input(11);
output(2, 30) <= input(12);
output(2, 31) <= input(13);
output(2, 32) <= input(51);
output(2, 33) <= input(52);
output(2, 34) <= input(53);
output(2, 35) <= input(54);
output(2, 36) <= input(55);
output(2, 37) <= input(19);
output(2, 38) <= input(20);
output(2, 39) <= input(21);
output(2, 40) <= input(22);
output(2, 41) <= input(23);
output(2, 42) <= input(24);
output(2, 43) <= input(25);
output(2, 44) <= input(26);
output(2, 45) <= input(27);
output(2, 46) <= input(28);
output(2, 47) <= input(29);
output(2, 48) <= input(51);
output(2, 49) <= input(52);
output(2, 50) <= input(53);
output(2, 51) <= input(54);
output(2, 52) <= input(55);
output(2, 53) <= input(19);
output(2, 54) <= input(20);
output(2, 55) <= input(21);
output(2, 56) <= input(22);
output(2, 57) <= input(23);
output(2, 58) <= input(24);
output(2, 59) <= input(25);
output(2, 60) <= input(26);
output(2, 61) <= input(27);
output(2, 62) <= input(28);
output(2, 63) <= input(29);
output(2, 64) <= input(56);
output(2, 65) <= input(46);
output(2, 66) <= input(47);
output(2, 67) <= input(48);
output(2, 68) <= input(49);
output(2, 69) <= input(50);
output(2, 70) <= input(3);
output(2, 71) <= input(4);
output(2, 72) <= input(5);
output(2, 73) <= input(6);
output(2, 74) <= input(7);
output(2, 75) <= input(8);
output(2, 76) <= input(9);
output(2, 77) <= input(10);
output(2, 78) <= input(11);
output(2, 79) <= input(12);
output(2, 80) <= input(56);
output(2, 81) <= input(46);
output(2, 82) <= input(47);
output(2, 83) <= input(48);
output(2, 84) <= input(49);
output(2, 85) <= input(50);
output(2, 86) <= input(3);
output(2, 87) <= input(4);
output(2, 88) <= input(5);
output(2, 89) <= input(6);
output(2, 90) <= input(7);
output(2, 91) <= input(8);
output(2, 92) <= input(9);
output(2, 93) <= input(10);
output(2, 94) <= input(11);
output(2, 95) <= input(12);
output(2, 96) <= input(57);
output(2, 97) <= input(51);
output(2, 98) <= input(52);
output(2, 99) <= input(53);
output(2, 100) <= input(54);
output(2, 101) <= input(55);
output(2, 102) <= input(19);
output(2, 103) <= input(20);
output(2, 104) <= input(21);
output(2, 105) <= input(22);
output(2, 106) <= input(23);
output(2, 107) <= input(24);
output(2, 108) <= input(25);
output(2, 109) <= input(26);
output(2, 110) <= input(27);
output(2, 111) <= input(28);
output(2, 112) <= input(57);
output(2, 113) <= input(51);
output(2, 114) <= input(52);
output(2, 115) <= input(53);
output(2, 116) <= input(54);
output(2, 117) <= input(55);
output(2, 118) <= input(19);
output(2, 119) <= input(20);
output(2, 120) <= input(21);
output(2, 121) <= input(22);
output(2, 122) <= input(23);
output(2, 123) <= input(24);
output(2, 124) <= input(25);
output(2, 125) <= input(26);
output(2, 126) <= input(27);
output(2, 127) <= input(28);
output(2, 128) <= input(58);
output(2, 129) <= input(56);
output(2, 130) <= input(46);
output(2, 131) <= input(47);
output(2, 132) <= input(48);
output(2, 133) <= input(49);
output(2, 134) <= input(50);
output(2, 135) <= input(3);
output(2, 136) <= input(4);
output(2, 137) <= input(5);
output(2, 138) <= input(6);
output(2, 139) <= input(7);
output(2, 140) <= input(8);
output(2, 141) <= input(9);
output(2, 142) <= input(10);
output(2, 143) <= input(11);
output(2, 144) <= input(58);
output(2, 145) <= input(56);
output(2, 146) <= input(46);
output(2, 147) <= input(47);
output(2, 148) <= input(48);
output(2, 149) <= input(49);
output(2, 150) <= input(50);
output(2, 151) <= input(3);
output(2, 152) <= input(4);
output(2, 153) <= input(5);
output(2, 154) <= input(6);
output(2, 155) <= input(7);
output(2, 156) <= input(8);
output(2, 157) <= input(9);
output(2, 158) <= input(10);
output(2, 159) <= input(11);
output(2, 160) <= input(59);
output(2, 161) <= input(57);
output(2, 162) <= input(51);
output(2, 163) <= input(52);
output(2, 164) <= input(53);
output(2, 165) <= input(54);
output(2, 166) <= input(55);
output(2, 167) <= input(19);
output(2, 168) <= input(20);
output(2, 169) <= input(21);
output(2, 170) <= input(22);
output(2, 171) <= input(23);
output(2, 172) <= input(24);
output(2, 173) <= input(25);
output(2, 174) <= input(26);
output(2, 175) <= input(27);
output(2, 176) <= input(59);
output(2, 177) <= input(57);
output(2, 178) <= input(51);
output(2, 179) <= input(52);
output(2, 180) <= input(53);
output(2, 181) <= input(54);
output(2, 182) <= input(55);
output(2, 183) <= input(19);
output(2, 184) <= input(20);
output(2, 185) <= input(21);
output(2, 186) <= input(22);
output(2, 187) <= input(23);
output(2, 188) <= input(24);
output(2, 189) <= input(25);
output(2, 190) <= input(26);
output(2, 191) <= input(27);
output(2, 192) <= input(60);
output(2, 193) <= input(58);
output(2, 194) <= input(56);
output(2, 195) <= input(46);
output(2, 196) <= input(47);
output(2, 197) <= input(48);
output(2, 198) <= input(49);
output(2, 199) <= input(50);
output(2, 200) <= input(3);
output(2, 201) <= input(4);
output(2, 202) <= input(5);
output(2, 203) <= input(6);
output(2, 204) <= input(7);
output(2, 205) <= input(8);
output(2, 206) <= input(9);
output(2, 207) <= input(10);
output(2, 208) <= input(60);
output(2, 209) <= input(58);
output(2, 210) <= input(56);
output(2, 211) <= input(46);
output(2, 212) <= input(47);
output(2, 213) <= input(48);
output(2, 214) <= input(49);
output(2, 215) <= input(50);
output(2, 216) <= input(3);
output(2, 217) <= input(4);
output(2, 218) <= input(5);
output(2, 219) <= input(6);
output(2, 220) <= input(7);
output(2, 221) <= input(8);
output(2, 222) <= input(9);
output(2, 223) <= input(10);
output(2, 224) <= input(61);
output(2, 225) <= input(59);
output(2, 226) <= input(57);
output(2, 227) <= input(51);
output(2, 228) <= input(52);
output(2, 229) <= input(53);
output(2, 230) <= input(54);
output(2, 231) <= input(55);
output(2, 232) <= input(19);
output(2, 233) <= input(20);
output(2, 234) <= input(21);
output(2, 235) <= input(22);
output(2, 236) <= input(23);
output(2, 237) <= input(24);
output(2, 238) <= input(25);
output(2, 239) <= input(26);
output(2, 240) <= input(61);
output(2, 241) <= input(59);
output(2, 242) <= input(57);
output(2, 243) <= input(51);
output(2, 244) <= input(52);
output(2, 245) <= input(53);
output(2, 246) <= input(54);
output(2, 247) <= input(55);
output(2, 248) <= input(19);
output(2, 249) <= input(20);
output(2, 250) <= input(21);
output(2, 251) <= input(22);
output(2, 252) <= input(23);
output(2, 253) <= input(24);
output(2, 254) <= input(25);
output(2, 255) <= input(26);
when "0100" =>
output(0, 0) <= input(0);
output(0, 1) <= input(1);
output(0, 2) <= input(2);
output(0, 3) <= input(3);
output(0, 4) <= input(4);
output(0, 5) <= input(5);
output(0, 6) <= input(6);
output(0, 7) <= input(7);
output(0, 8) <= input(8);
output(0, 9) <= input(9);
output(0, 10) <= input(10);
output(0, 11) <= input(11);
output(0, 12) <= input(12);
output(0, 13) <= input(13);
output(0, 14) <= input(14);
output(0, 15) <= input(15);
output(0, 16) <= input(16);
output(0, 17) <= input(17);
output(0, 18) <= input(18);
output(0, 19) <= input(19);
output(0, 20) <= input(20);
output(0, 21) <= input(21);
output(0, 22) <= input(22);
output(0, 23) <= input(23);
output(0, 24) <= input(24);
output(0, 25) <= input(25);
output(0, 26) <= input(26);
output(0, 27) <= input(27);
output(0, 28) <= input(28);
output(0, 29) <= input(29);
output(0, 30) <= input(30);
output(0, 31) <= input(31);
output(0, 32) <= input(16);
output(0, 33) <= input(17);
output(0, 34) <= input(18);
output(0, 35) <= input(19);
output(0, 36) <= input(20);
output(0, 37) <= input(21);
output(0, 38) <= input(22);
output(0, 39) <= input(23);
output(0, 40) <= input(24);
output(0, 41) <= input(25);
output(0, 42) <= input(26);
output(0, 43) <= input(27);
output(0, 44) <= input(28);
output(0, 45) <= input(29);
output(0, 46) <= input(30);
output(0, 47) <= input(31);
output(0, 48) <= input(32);
output(0, 49) <= input(0);
output(0, 50) <= input(1);
output(0, 51) <= input(2);
output(0, 52) <= input(3);
output(0, 53) <= input(4);
output(0, 54) <= input(5);
output(0, 55) <= input(6);
output(0, 56) <= input(7);
output(0, 57) <= input(8);
output(0, 58) <= input(9);
output(0, 59) <= input(10);
output(0, 60) <= input(11);
output(0, 61) <= input(12);
output(0, 62) <= input(13);
output(0, 63) <= input(14);
output(0, 64) <= input(33);
output(0, 65) <= input(16);
output(0, 66) <= input(17);
output(0, 67) <= input(18);
output(0, 68) <= input(19);
output(0, 69) <= input(20);
output(0, 70) <= input(21);
output(0, 71) <= input(22);
output(0, 72) <= input(23);
output(0, 73) <= input(24);
output(0, 74) <= input(25);
output(0, 75) <= input(26);
output(0, 76) <= input(27);
output(0, 77) <= input(28);
output(0, 78) <= input(29);
output(0, 79) <= input(30);
output(0, 80) <= input(33);
output(0, 81) <= input(16);
output(0, 82) <= input(17);
output(0, 83) <= input(18);
output(0, 84) <= input(19);
output(0, 85) <= input(20);
output(0, 86) <= input(21);
output(0, 87) <= input(22);
output(0, 88) <= input(23);
output(0, 89) <= input(24);
output(0, 90) <= input(25);
output(0, 91) <= input(26);
output(0, 92) <= input(27);
output(0, 93) <= input(28);
output(0, 94) <= input(29);
output(0, 95) <= input(30);
output(0, 96) <= input(34);
output(0, 97) <= input(32);
output(0, 98) <= input(0);
output(0, 99) <= input(1);
output(0, 100) <= input(2);
output(0, 101) <= input(3);
output(0, 102) <= input(4);
output(0, 103) <= input(5);
output(0, 104) <= input(6);
output(0, 105) <= input(7);
output(0, 106) <= input(8);
output(0, 107) <= input(9);
output(0, 108) <= input(10);
output(0, 109) <= input(11);
output(0, 110) <= input(12);
output(0, 111) <= input(13);
output(0, 112) <= input(34);
output(0, 113) <= input(32);
output(0, 114) <= input(0);
output(0, 115) <= input(1);
output(0, 116) <= input(2);
output(0, 117) <= input(3);
output(0, 118) <= input(4);
output(0, 119) <= input(5);
output(0, 120) <= input(6);
output(0, 121) <= input(7);
output(0, 122) <= input(8);
output(0, 123) <= input(9);
output(0, 124) <= input(10);
output(0, 125) <= input(11);
output(0, 126) <= input(12);
output(0, 127) <= input(13);
output(0, 128) <= input(35);
output(0, 129) <= input(33);
output(0, 130) <= input(16);
output(0, 131) <= input(17);
output(0, 132) <= input(18);
output(0, 133) <= input(19);
output(0, 134) <= input(20);
output(0, 135) <= input(21);
output(0, 136) <= input(22);
output(0, 137) <= input(23);
output(0, 138) <= input(24);
output(0, 139) <= input(25);
output(0, 140) <= input(26);
output(0, 141) <= input(27);
output(0, 142) <= input(28);
output(0, 143) <= input(29);
output(0, 144) <= input(36);
output(0, 145) <= input(34);
output(0, 146) <= input(32);
output(0, 147) <= input(0);
output(0, 148) <= input(1);
output(0, 149) <= input(2);
output(0, 150) <= input(3);
output(0, 151) <= input(4);
output(0, 152) <= input(5);
output(0, 153) <= input(6);
output(0, 154) <= input(7);
output(0, 155) <= input(8);
output(0, 156) <= input(9);
output(0, 157) <= input(10);
output(0, 158) <= input(11);
output(0, 159) <= input(12);
output(0, 160) <= input(36);
output(0, 161) <= input(34);
output(0, 162) <= input(32);
output(0, 163) <= input(0);
output(0, 164) <= input(1);
output(0, 165) <= input(2);
output(0, 166) <= input(3);
output(0, 167) <= input(4);
output(0, 168) <= input(5);
output(0, 169) <= input(6);
output(0, 170) <= input(7);
output(0, 171) <= input(8);
output(0, 172) <= input(9);
output(0, 173) <= input(10);
output(0, 174) <= input(11);
output(0, 175) <= input(12);
output(0, 176) <= input(37);
output(0, 177) <= input(35);
output(0, 178) <= input(33);
output(0, 179) <= input(16);
output(0, 180) <= input(17);
output(0, 181) <= input(18);
output(0, 182) <= input(19);
output(0, 183) <= input(20);
output(0, 184) <= input(21);
output(0, 185) <= input(22);
output(0, 186) <= input(23);
output(0, 187) <= input(24);
output(0, 188) <= input(25);
output(0, 189) <= input(26);
output(0, 190) <= input(27);
output(0, 191) <= input(28);
output(0, 192) <= input(38);
output(0, 193) <= input(36);
output(0, 194) <= input(34);
output(0, 195) <= input(32);
output(0, 196) <= input(0);
output(0, 197) <= input(1);
output(0, 198) <= input(2);
output(0, 199) <= input(3);
output(0, 200) <= input(4);
output(0, 201) <= input(5);
output(0, 202) <= input(6);
output(0, 203) <= input(7);
output(0, 204) <= input(8);
output(0, 205) <= input(9);
output(0, 206) <= input(10);
output(0, 207) <= input(11);
output(0, 208) <= input(38);
output(0, 209) <= input(36);
output(0, 210) <= input(34);
output(0, 211) <= input(32);
output(0, 212) <= input(0);
output(0, 213) <= input(1);
output(0, 214) <= input(2);
output(0, 215) <= input(3);
output(0, 216) <= input(4);
output(0, 217) <= input(5);
output(0, 218) <= input(6);
output(0, 219) <= input(7);
output(0, 220) <= input(8);
output(0, 221) <= input(9);
output(0, 222) <= input(10);
output(0, 223) <= input(11);
output(0, 224) <= input(39);
output(0, 225) <= input(37);
output(0, 226) <= input(35);
output(0, 227) <= input(33);
output(0, 228) <= input(16);
output(0, 229) <= input(17);
output(0, 230) <= input(18);
output(0, 231) <= input(19);
output(0, 232) <= input(20);
output(0, 233) <= input(21);
output(0, 234) <= input(22);
output(0, 235) <= input(23);
output(0, 236) <= input(24);
output(0, 237) <= input(25);
output(0, 238) <= input(26);
output(0, 239) <= input(27);
output(0, 240) <= input(39);
output(0, 241) <= input(37);
output(0, 242) <= input(35);
output(0, 243) <= input(33);
output(0, 244) <= input(16);
output(0, 245) <= input(17);
output(0, 246) <= input(18);
output(0, 247) <= input(19);
output(0, 248) <= input(20);
output(0, 249) <= input(21);
output(0, 250) <= input(22);
output(0, 251) <= input(23);
output(0, 252) <= input(24);
output(0, 253) <= input(25);
output(0, 254) <= input(26);
output(0, 255) <= input(27);
output(1, 0) <= input(40);
output(1, 1) <= input(41);
output(1, 2) <= input(42);
output(1, 3) <= input(43);
output(1, 4) <= input(44);
output(1, 5) <= input(45);
output(1, 6) <= input(5);
output(1, 7) <= input(6);
output(1, 8) <= input(7);
output(1, 9) <= input(8);
output(1, 10) <= input(9);
output(1, 11) <= input(10);
output(1, 12) <= input(11);
output(1, 13) <= input(12);
output(1, 14) <= input(13);
output(1, 15) <= input(14);
output(1, 16) <= input(46);
output(1, 17) <= input(47);
output(1, 18) <= input(48);
output(1, 19) <= input(49);
output(1, 20) <= input(50);
output(1, 21) <= input(51);
output(1, 22) <= input(21);
output(1, 23) <= input(22);
output(1, 24) <= input(23);
output(1, 25) <= input(24);
output(1, 26) <= input(25);
output(1, 27) <= input(26);
output(1, 28) <= input(27);
output(1, 29) <= input(28);
output(1, 30) <= input(29);
output(1, 31) <= input(30);
output(1, 32) <= input(52);
output(1, 33) <= input(40);
output(1, 34) <= input(41);
output(1, 35) <= input(42);
output(1, 36) <= input(43);
output(1, 37) <= input(44);
output(1, 38) <= input(45);
output(1, 39) <= input(5);
output(1, 40) <= input(6);
output(1, 41) <= input(7);
output(1, 42) <= input(8);
output(1, 43) <= input(9);
output(1, 44) <= input(10);
output(1, 45) <= input(11);
output(1, 46) <= input(12);
output(1, 47) <= input(13);
output(1, 48) <= input(52);
output(1, 49) <= input(40);
output(1, 50) <= input(41);
output(1, 51) <= input(42);
output(1, 52) <= input(43);
output(1, 53) <= input(44);
output(1, 54) <= input(45);
output(1, 55) <= input(5);
output(1, 56) <= input(6);
output(1, 57) <= input(7);
output(1, 58) <= input(8);
output(1, 59) <= input(9);
output(1, 60) <= input(10);
output(1, 61) <= input(11);
output(1, 62) <= input(12);
output(1, 63) <= input(13);
output(1, 64) <= input(53);
output(1, 65) <= input(46);
output(1, 66) <= input(47);
output(1, 67) <= input(48);
output(1, 68) <= input(49);
output(1, 69) <= input(50);
output(1, 70) <= input(51);
output(1, 71) <= input(21);
output(1, 72) <= input(22);
output(1, 73) <= input(23);
output(1, 74) <= input(24);
output(1, 75) <= input(25);
output(1, 76) <= input(26);
output(1, 77) <= input(27);
output(1, 78) <= input(28);
output(1, 79) <= input(29);
output(1, 80) <= input(54);
output(1, 81) <= input(52);
output(1, 82) <= input(40);
output(1, 83) <= input(41);
output(1, 84) <= input(42);
output(1, 85) <= input(43);
output(1, 86) <= input(44);
output(1, 87) <= input(45);
output(1, 88) <= input(5);
output(1, 89) <= input(6);
output(1, 90) <= input(7);
output(1, 91) <= input(8);
output(1, 92) <= input(9);
output(1, 93) <= input(10);
output(1, 94) <= input(11);
output(1, 95) <= input(12);
output(1, 96) <= input(55);
output(1, 97) <= input(53);
output(1, 98) <= input(46);
output(1, 99) <= input(47);
output(1, 100) <= input(48);
output(1, 101) <= input(49);
output(1, 102) <= input(50);
output(1, 103) <= input(51);
output(1, 104) <= input(21);
output(1, 105) <= input(22);
output(1, 106) <= input(23);
output(1, 107) <= input(24);
output(1, 108) <= input(25);
output(1, 109) <= input(26);
output(1, 110) <= input(27);
output(1, 111) <= input(28);
output(1, 112) <= input(55);
output(1, 113) <= input(53);
output(1, 114) <= input(46);
output(1, 115) <= input(47);
output(1, 116) <= input(48);
output(1, 117) <= input(49);
output(1, 118) <= input(50);
output(1, 119) <= input(51);
output(1, 120) <= input(21);
output(1, 121) <= input(22);
output(1, 122) <= input(23);
output(1, 123) <= input(24);
output(1, 124) <= input(25);
output(1, 125) <= input(26);
output(1, 126) <= input(27);
output(1, 127) <= input(28);
output(1, 128) <= input(56);
output(1, 129) <= input(54);
output(1, 130) <= input(52);
output(1, 131) <= input(40);
output(1, 132) <= input(41);
output(1, 133) <= input(42);
output(1, 134) <= input(43);
output(1, 135) <= input(44);
output(1, 136) <= input(45);
output(1, 137) <= input(5);
output(1, 138) <= input(6);
output(1, 139) <= input(7);
output(1, 140) <= input(8);
output(1, 141) <= input(9);
output(1, 142) <= input(10);
output(1, 143) <= input(11);
output(1, 144) <= input(57);
output(1, 145) <= input(55);
output(1, 146) <= input(53);
output(1, 147) <= input(46);
output(1, 148) <= input(47);
output(1, 149) <= input(48);
output(1, 150) <= input(49);
output(1, 151) <= input(50);
output(1, 152) <= input(51);
output(1, 153) <= input(21);
output(1, 154) <= input(22);
output(1, 155) <= input(23);
output(1, 156) <= input(24);
output(1, 157) <= input(25);
output(1, 158) <= input(26);
output(1, 159) <= input(27);
output(1, 160) <= input(58);
output(1, 161) <= input(56);
output(1, 162) <= input(54);
output(1, 163) <= input(52);
output(1, 164) <= input(40);
output(1, 165) <= input(41);
output(1, 166) <= input(42);
output(1, 167) <= input(43);
output(1, 168) <= input(44);
output(1, 169) <= input(45);
output(1, 170) <= input(5);
output(1, 171) <= input(6);
output(1, 172) <= input(7);
output(1, 173) <= input(8);
output(1, 174) <= input(9);
output(1, 175) <= input(10);
output(1, 176) <= input(58);
output(1, 177) <= input(56);
output(1, 178) <= input(54);
output(1, 179) <= input(52);
output(1, 180) <= input(40);
output(1, 181) <= input(41);
output(1, 182) <= input(42);
output(1, 183) <= input(43);
output(1, 184) <= input(44);
output(1, 185) <= input(45);
output(1, 186) <= input(5);
output(1, 187) <= input(6);
output(1, 188) <= input(7);
output(1, 189) <= input(8);
output(1, 190) <= input(9);
output(1, 191) <= input(10);
output(1, 192) <= input(59);
output(1, 193) <= input(57);
output(1, 194) <= input(55);
output(1, 195) <= input(53);
output(1, 196) <= input(46);
output(1, 197) <= input(47);
output(1, 198) <= input(48);
output(1, 199) <= input(49);
output(1, 200) <= input(50);
output(1, 201) <= input(51);
output(1, 202) <= input(21);
output(1, 203) <= input(22);
output(1, 204) <= input(23);
output(1, 205) <= input(24);
output(1, 206) <= input(25);
output(1, 207) <= input(26);
output(1, 208) <= input(60);
output(1, 209) <= input(58);
output(1, 210) <= input(56);
output(1, 211) <= input(54);
output(1, 212) <= input(52);
output(1, 213) <= input(40);
output(1, 214) <= input(41);
output(1, 215) <= input(42);
output(1, 216) <= input(43);
output(1, 217) <= input(44);
output(1, 218) <= input(45);
output(1, 219) <= input(5);
output(1, 220) <= input(6);
output(1, 221) <= input(7);
output(1, 222) <= input(8);
output(1, 223) <= input(9);
output(1, 224) <= input(61);
output(1, 225) <= input(59);
output(1, 226) <= input(57);
output(1, 227) <= input(55);
output(1, 228) <= input(53);
output(1, 229) <= input(46);
output(1, 230) <= input(47);
output(1, 231) <= input(48);
output(1, 232) <= input(49);
output(1, 233) <= input(50);
output(1, 234) <= input(51);
output(1, 235) <= input(21);
output(1, 236) <= input(22);
output(1, 237) <= input(23);
output(1, 238) <= input(24);
output(1, 239) <= input(25);
output(1, 240) <= input(61);
output(1, 241) <= input(59);
output(1, 242) <= input(57);
output(1, 243) <= input(55);
output(1, 244) <= input(53);
output(1, 245) <= input(46);
output(1, 246) <= input(47);
output(1, 247) <= input(48);
output(1, 248) <= input(49);
output(1, 249) <= input(50);
output(1, 250) <= input(51);
output(1, 251) <= input(21);
output(1, 252) <= input(22);
output(1, 253) <= input(23);
output(1, 254) <= input(24);
output(1, 255) <= input(25);
output(2, 0) <= input(62);
output(2, 1) <= input(63);
output(2, 2) <= input(64);
output(2, 3) <= input(65);
output(2, 4) <= input(66);
output(2, 5) <= input(67);
output(2, 6) <= input(68);
output(2, 7) <= input(69);
output(2, 8) <= input(6);
output(2, 9) <= input(7);
output(2, 10) <= input(8);
output(2, 11) <= input(9);
output(2, 12) <= input(10);
output(2, 13) <= input(11);
output(2, 14) <= input(12);
output(2, 15) <= input(13);
output(2, 16) <= input(70);
output(2, 17) <= input(71);
output(2, 18) <= input(72);
output(2, 19) <= input(73);
output(2, 20) <= input(74);
output(2, 21) <= input(75);
output(2, 22) <= input(76);
output(2, 23) <= input(77);
output(2, 24) <= input(22);
output(2, 25) <= input(23);
output(2, 26) <= input(24);
output(2, 27) <= input(25);
output(2, 28) <= input(26);
output(2, 29) <= input(27);
output(2, 30) <= input(28);
output(2, 31) <= input(29);
output(2, 32) <= input(78);
output(2, 33) <= input(62);
output(2, 34) <= input(63);
output(2, 35) <= input(64);
output(2, 36) <= input(65);
output(2, 37) <= input(66);
output(2, 38) <= input(67);
output(2, 39) <= input(68);
output(2, 40) <= input(69);
output(2, 41) <= input(6);
output(2, 42) <= input(7);
output(2, 43) <= input(8);
output(2, 44) <= input(9);
output(2, 45) <= input(10);
output(2, 46) <= input(11);
output(2, 47) <= input(12);
output(2, 48) <= input(79);
output(2, 49) <= input(70);
output(2, 50) <= input(71);
output(2, 51) <= input(72);
output(2, 52) <= input(73);
output(2, 53) <= input(74);
output(2, 54) <= input(75);
output(2, 55) <= input(76);
output(2, 56) <= input(77);
output(2, 57) <= input(22);
output(2, 58) <= input(23);
output(2, 59) <= input(24);
output(2, 60) <= input(25);
output(2, 61) <= input(26);
output(2, 62) <= input(27);
output(2, 63) <= input(28);
output(2, 64) <= input(80);
output(2, 65) <= input(78);
output(2, 66) <= input(62);
output(2, 67) <= input(63);
output(2, 68) <= input(64);
output(2, 69) <= input(65);
output(2, 70) <= input(66);
output(2, 71) <= input(67);
output(2, 72) <= input(68);
output(2, 73) <= input(69);
output(2, 74) <= input(6);
output(2, 75) <= input(7);
output(2, 76) <= input(8);
output(2, 77) <= input(9);
output(2, 78) <= input(10);
output(2, 79) <= input(11);
output(2, 80) <= input(81);
output(2, 81) <= input(79);
output(2, 82) <= input(70);
output(2, 83) <= input(71);
output(2, 84) <= input(72);
output(2, 85) <= input(73);
output(2, 86) <= input(74);
output(2, 87) <= input(75);
output(2, 88) <= input(76);
output(2, 89) <= input(77);
output(2, 90) <= input(22);
output(2, 91) <= input(23);
output(2, 92) <= input(24);
output(2, 93) <= input(25);
output(2, 94) <= input(26);
output(2, 95) <= input(27);
output(2, 96) <= input(82);
output(2, 97) <= input(80);
output(2, 98) <= input(78);
output(2, 99) <= input(62);
output(2, 100) <= input(63);
output(2, 101) <= input(64);
output(2, 102) <= input(65);
output(2, 103) <= input(66);
output(2, 104) <= input(67);
output(2, 105) <= input(68);
output(2, 106) <= input(69);
output(2, 107) <= input(6);
output(2, 108) <= input(7);
output(2, 109) <= input(8);
output(2, 110) <= input(9);
output(2, 111) <= input(10);
output(2, 112) <= input(82);
output(2, 113) <= input(80);
output(2, 114) <= input(78);
output(2, 115) <= input(62);
output(2, 116) <= input(63);
output(2, 117) <= input(64);
output(2, 118) <= input(65);
output(2, 119) <= input(66);
output(2, 120) <= input(67);
output(2, 121) <= input(68);
output(2, 122) <= input(69);
output(2, 123) <= input(6);
output(2, 124) <= input(7);
output(2, 125) <= input(8);
output(2, 126) <= input(9);
output(2, 127) <= input(10);
output(2, 128) <= input(83);
output(2, 129) <= input(81);
output(2, 130) <= input(79);
output(2, 131) <= input(70);
output(2, 132) <= input(71);
output(2, 133) <= input(72);
output(2, 134) <= input(73);
output(2, 135) <= input(74);
output(2, 136) <= input(75);
output(2, 137) <= input(76);
output(2, 138) <= input(77);
output(2, 139) <= input(22);
output(2, 140) <= input(23);
output(2, 141) <= input(24);
output(2, 142) <= input(25);
output(2, 143) <= input(26);
output(2, 144) <= input(84);
output(2, 145) <= input(82);
output(2, 146) <= input(80);
output(2, 147) <= input(78);
output(2, 148) <= input(62);
output(2, 149) <= input(63);
output(2, 150) <= input(64);
output(2, 151) <= input(65);
output(2, 152) <= input(66);
output(2, 153) <= input(67);
output(2, 154) <= input(68);
output(2, 155) <= input(69);
output(2, 156) <= input(6);
output(2, 157) <= input(7);
output(2, 158) <= input(8);
output(2, 159) <= input(9);
output(2, 160) <= input(85);
output(2, 161) <= input(83);
output(2, 162) <= input(81);
output(2, 163) <= input(79);
output(2, 164) <= input(70);
output(2, 165) <= input(71);
output(2, 166) <= input(72);
output(2, 167) <= input(73);
output(2, 168) <= input(74);
output(2, 169) <= input(75);
output(2, 170) <= input(76);
output(2, 171) <= input(77);
output(2, 172) <= input(22);
output(2, 173) <= input(23);
output(2, 174) <= input(24);
output(2, 175) <= input(25);
output(2, 176) <= input(86);
output(2, 177) <= input(84);
output(2, 178) <= input(82);
output(2, 179) <= input(80);
output(2, 180) <= input(78);
output(2, 181) <= input(62);
output(2, 182) <= input(63);
output(2, 183) <= input(64);
output(2, 184) <= input(65);
output(2, 185) <= input(66);
output(2, 186) <= input(67);
output(2, 187) <= input(68);
output(2, 188) <= input(69);
output(2, 189) <= input(6);
output(2, 190) <= input(7);
output(2, 191) <= input(8);
output(2, 192) <= input(87);
output(2, 193) <= input(85);
output(2, 194) <= input(83);
output(2, 195) <= input(81);
output(2, 196) <= input(79);
output(2, 197) <= input(70);
output(2, 198) <= input(71);
output(2, 199) <= input(72);
output(2, 200) <= input(73);
output(2, 201) <= input(74);
output(2, 202) <= input(75);
output(2, 203) <= input(76);
output(2, 204) <= input(77);
output(2, 205) <= input(22);
output(2, 206) <= input(23);
output(2, 207) <= input(24);
output(2, 208) <= input(88);
output(2, 209) <= input(86);
output(2, 210) <= input(84);
output(2, 211) <= input(82);
output(2, 212) <= input(80);
output(2, 213) <= input(78);
output(2, 214) <= input(62);
output(2, 215) <= input(63);
output(2, 216) <= input(64);
output(2, 217) <= input(65);
output(2, 218) <= input(66);
output(2, 219) <= input(67);
output(2, 220) <= input(68);
output(2, 221) <= input(69);
output(2, 222) <= input(6);
output(2, 223) <= input(7);
output(2, 224) <= input(89);
output(2, 225) <= input(87);
output(2, 226) <= input(85);
output(2, 227) <= input(83);
output(2, 228) <= input(81);
output(2, 229) <= input(79);
output(2, 230) <= input(70);
output(2, 231) <= input(71);
output(2, 232) <= input(72);
output(2, 233) <= input(73);
output(2, 234) <= input(74);
output(2, 235) <= input(75);
output(2, 236) <= input(76);
output(2, 237) <= input(77);
output(2, 238) <= input(22);
output(2, 239) <= input(23);
output(2, 240) <= input(89);
output(2, 241) <= input(87);
output(2, 242) <= input(85);
output(2, 243) <= input(83);
output(2, 244) <= input(81);
output(2, 245) <= input(79);
output(2, 246) <= input(70);
output(2, 247) <= input(71);
output(2, 248) <= input(72);
output(2, 249) <= input(73);
output(2, 250) <= input(74);
output(2, 251) <= input(75);
output(2, 252) <= input(76);
output(2, 253) <= input(77);
output(2, 254) <= input(22);
output(2, 255) <= input(23);
when "0101" =>
output(0, 0) <= input(0);
output(0, 1) <= input(1);
output(0, 2) <= input(2);
output(0, 3) <= input(3);
output(0, 4) <= input(4);
output(0, 5) <= input(5);
output(0, 6) <= input(6);
output(0, 7) <= input(7);
output(0, 8) <= input(8);
output(0, 9) <= input(9);
output(0, 10) <= input(10);
output(0, 11) <= input(11);
output(0, 12) <= input(12);
output(0, 13) <= input(13);
output(0, 14) <= input(14);
output(0, 15) <= input(15);
output(0, 16) <= input(16);
output(0, 17) <= input(17);
output(0, 18) <= input(18);
output(0, 19) <= input(19);
output(0, 20) <= input(20);
output(0, 21) <= input(21);
output(0, 22) <= input(22);
output(0, 23) <= input(23);
output(0, 24) <= input(24);
output(0, 25) <= input(25);
output(0, 26) <= input(26);
output(0, 27) <= input(27);
output(0, 28) <= input(28);
output(0, 29) <= input(29);
output(0, 30) <= input(30);
output(0, 31) <= input(31);
output(0, 32) <= input(32);
output(0, 33) <= input(0);
output(0, 34) <= input(1);
output(0, 35) <= input(2);
output(0, 36) <= input(3);
output(0, 37) <= input(4);
output(0, 38) <= input(5);
output(0, 39) <= input(6);
output(0, 40) <= input(7);
output(0, 41) <= input(8);
output(0, 42) <= input(9);
output(0, 43) <= input(10);
output(0, 44) <= input(11);
output(0, 45) <= input(12);
output(0, 46) <= input(13);
output(0, 47) <= input(14);
output(0, 48) <= input(33);
output(0, 49) <= input(16);
output(0, 50) <= input(17);
output(0, 51) <= input(18);
output(0, 52) <= input(19);
output(0, 53) <= input(20);
output(0, 54) <= input(21);
output(0, 55) <= input(22);
output(0, 56) <= input(23);
output(0, 57) <= input(24);
output(0, 58) <= input(25);
output(0, 59) <= input(26);
output(0, 60) <= input(27);
output(0, 61) <= input(28);
output(0, 62) <= input(29);
output(0, 63) <= input(30);
output(0, 64) <= input(34);
output(0, 65) <= input(32);
output(0, 66) <= input(0);
output(0, 67) <= input(1);
output(0, 68) <= input(2);
output(0, 69) <= input(3);
output(0, 70) <= input(4);
output(0, 71) <= input(5);
output(0, 72) <= input(6);
output(0, 73) <= input(7);
output(0, 74) <= input(8);
output(0, 75) <= input(9);
output(0, 76) <= input(10);
output(0, 77) <= input(11);
output(0, 78) <= input(12);
output(0, 79) <= input(13);
output(0, 80) <= input(35);
output(0, 81) <= input(33);
output(0, 82) <= input(16);
output(0, 83) <= input(17);
output(0, 84) <= input(18);
output(0, 85) <= input(19);
output(0, 86) <= input(20);
output(0, 87) <= input(21);
output(0, 88) <= input(22);
output(0, 89) <= input(23);
output(0, 90) <= input(24);
output(0, 91) <= input(25);
output(0, 92) <= input(26);
output(0, 93) <= input(27);
output(0, 94) <= input(28);
output(0, 95) <= input(29);
output(0, 96) <= input(36);
output(0, 97) <= input(34);
output(0, 98) <= input(32);
output(0, 99) <= input(0);
output(0, 100) <= input(1);
output(0, 101) <= input(2);
output(0, 102) <= input(3);
output(0, 103) <= input(4);
output(0, 104) <= input(5);
output(0, 105) <= input(6);
output(0, 106) <= input(7);
output(0, 107) <= input(8);
output(0, 108) <= input(9);
output(0, 109) <= input(10);
output(0, 110) <= input(11);
output(0, 111) <= input(12);
output(0, 112) <= input(37);
output(0, 113) <= input(35);
output(0, 114) <= input(33);
output(0, 115) <= input(16);
output(0, 116) <= input(17);
output(0, 117) <= input(18);
output(0, 118) <= input(19);
output(0, 119) <= input(20);
output(0, 120) <= input(21);
output(0, 121) <= input(22);
output(0, 122) <= input(23);
output(0, 123) <= input(24);
output(0, 124) <= input(25);
output(0, 125) <= input(26);
output(0, 126) <= input(27);
output(0, 127) <= input(28);
output(0, 128) <= input(38);
output(0, 129) <= input(36);
output(0, 130) <= input(34);
output(0, 131) <= input(32);
output(0, 132) <= input(0);
output(0, 133) <= input(1);
output(0, 134) <= input(2);
output(0, 135) <= input(3);
output(0, 136) <= input(4);
output(0, 137) <= input(5);
output(0, 138) <= input(6);
output(0, 139) <= input(7);
output(0, 140) <= input(8);
output(0, 141) <= input(9);
output(0, 142) <= input(10);
output(0, 143) <= input(11);
output(0, 144) <= input(39);
output(0, 145) <= input(37);
output(0, 146) <= input(35);
output(0, 147) <= input(33);
output(0, 148) <= input(16);
output(0, 149) <= input(17);
output(0, 150) <= input(18);
output(0, 151) <= input(19);
output(0, 152) <= input(20);
output(0, 153) <= input(21);
output(0, 154) <= input(22);
output(0, 155) <= input(23);
output(0, 156) <= input(24);
output(0, 157) <= input(25);
output(0, 158) <= input(26);
output(0, 159) <= input(27);
output(0, 160) <= input(40);
output(0, 161) <= input(38);
output(0, 162) <= input(36);
output(0, 163) <= input(34);
output(0, 164) <= input(32);
output(0, 165) <= input(0);
output(0, 166) <= input(1);
output(0, 167) <= input(2);
output(0, 168) <= input(3);
output(0, 169) <= input(4);
output(0, 170) <= input(5);
output(0, 171) <= input(6);
output(0, 172) <= input(7);
output(0, 173) <= input(8);
output(0, 174) <= input(9);
output(0, 175) <= input(10);
output(0, 176) <= input(41);
output(0, 177) <= input(39);
output(0, 178) <= input(37);
output(0, 179) <= input(35);
output(0, 180) <= input(33);
output(0, 181) <= input(16);
output(0, 182) <= input(17);
output(0, 183) <= input(18);
output(0, 184) <= input(19);
output(0, 185) <= input(20);
output(0, 186) <= input(21);
output(0, 187) <= input(22);
output(0, 188) <= input(23);
output(0, 189) <= input(24);
output(0, 190) <= input(25);
output(0, 191) <= input(26);
output(0, 192) <= input(42);
output(0, 193) <= input(40);
output(0, 194) <= input(38);
output(0, 195) <= input(36);
output(0, 196) <= input(34);
output(0, 197) <= input(32);
output(0, 198) <= input(0);
output(0, 199) <= input(1);
output(0, 200) <= input(2);
output(0, 201) <= input(3);
output(0, 202) <= input(4);
output(0, 203) <= input(5);
output(0, 204) <= input(6);
output(0, 205) <= input(7);
output(0, 206) <= input(8);
output(0, 207) <= input(9);
output(0, 208) <= input(43);
output(0, 209) <= input(41);
output(0, 210) <= input(39);
output(0, 211) <= input(37);
output(0, 212) <= input(35);
output(0, 213) <= input(33);
output(0, 214) <= input(16);
output(0, 215) <= input(17);
output(0, 216) <= input(18);
output(0, 217) <= input(19);
output(0, 218) <= input(20);
output(0, 219) <= input(21);
output(0, 220) <= input(22);
output(0, 221) <= input(23);
output(0, 222) <= input(24);
output(0, 223) <= input(25);
output(0, 224) <= input(44);
output(0, 225) <= input(42);
output(0, 226) <= input(40);
output(0, 227) <= input(38);
output(0, 228) <= input(36);
output(0, 229) <= input(34);
output(0, 230) <= input(32);
output(0, 231) <= input(0);
output(0, 232) <= input(1);
output(0, 233) <= input(2);
output(0, 234) <= input(3);
output(0, 235) <= input(4);
output(0, 236) <= input(5);
output(0, 237) <= input(6);
output(0, 238) <= input(7);
output(0, 239) <= input(8);
output(0, 240) <= input(45);
output(0, 241) <= input(43);
output(0, 242) <= input(41);
output(0, 243) <= input(39);
output(0, 244) <= input(37);
output(0, 245) <= input(35);
output(0, 246) <= input(33);
output(0, 247) <= input(16);
output(0, 248) <= input(17);
output(0, 249) <= input(18);
output(0, 250) <= input(19);
output(0, 251) <= input(20);
output(0, 252) <= input(21);
output(0, 253) <= input(22);
output(0, 254) <= input(23);
output(0, 255) <= input(24);
output(1, 0) <= input(16);
output(1, 1) <= input(46);
output(1, 2) <= input(47);
output(1, 3) <= input(48);
output(1, 4) <= input(49);
output(1, 5) <= input(50);
output(1, 6) <= input(51);
output(1, 7) <= input(52);
output(1, 8) <= input(23);
output(1, 9) <= input(24);
output(1, 10) <= input(25);
output(1, 11) <= input(26);
output(1, 12) <= input(27);
output(1, 13) <= input(28);
output(1, 14) <= input(29);
output(1, 15) <= input(30);
output(1, 16) <= input(32);
output(1, 17) <= input(0);
output(1, 18) <= input(53);
output(1, 19) <= input(54);
output(1, 20) <= input(55);
output(1, 21) <= input(56);
output(1, 22) <= input(57);
output(1, 23) <= input(58);
output(1, 24) <= input(59);
output(1, 25) <= input(7);
output(1, 26) <= input(8);
output(1, 27) <= input(9);
output(1, 28) <= input(10);
output(1, 29) <= input(11);
output(1, 30) <= input(12);
output(1, 31) <= input(13);
output(1, 32) <= input(33);
output(1, 33) <= input(16);
output(1, 34) <= input(46);
output(1, 35) <= input(47);
output(1, 36) <= input(48);
output(1, 37) <= input(49);
output(1, 38) <= input(50);
output(1, 39) <= input(51);
output(1, 40) <= input(52);
output(1, 41) <= input(23);
output(1, 42) <= input(24);
output(1, 43) <= input(25);
output(1, 44) <= input(26);
output(1, 45) <= input(27);
output(1, 46) <= input(28);
output(1, 47) <= input(29);
output(1, 48) <= input(60);
output(1, 49) <= input(32);
output(1, 50) <= input(0);
output(1, 51) <= input(53);
output(1, 52) <= input(54);
output(1, 53) <= input(55);
output(1, 54) <= input(56);
output(1, 55) <= input(57);
output(1, 56) <= input(58);
output(1, 57) <= input(59);
output(1, 58) <= input(7);
output(1, 59) <= input(8);
output(1, 60) <= input(9);
output(1, 61) <= input(10);
output(1, 62) <= input(11);
output(1, 63) <= input(12);
output(1, 64) <= input(61);
output(1, 65) <= input(33);
output(1, 66) <= input(16);
output(1, 67) <= input(46);
output(1, 68) <= input(47);
output(1, 69) <= input(48);
output(1, 70) <= input(49);
output(1, 71) <= input(50);
output(1, 72) <= input(51);
output(1, 73) <= input(52);
output(1, 74) <= input(23);
output(1, 75) <= input(24);
output(1, 76) <= input(25);
output(1, 77) <= input(26);
output(1, 78) <= input(27);
output(1, 79) <= input(28);
output(1, 80) <= input(62);
output(1, 81) <= input(60);
output(1, 82) <= input(32);
output(1, 83) <= input(0);
output(1, 84) <= input(53);
output(1, 85) <= input(54);
output(1, 86) <= input(55);
output(1, 87) <= input(56);
output(1, 88) <= input(57);
output(1, 89) <= input(58);
output(1, 90) <= input(59);
output(1, 91) <= input(7);
output(1, 92) <= input(8);
output(1, 93) <= input(9);
output(1, 94) <= input(10);
output(1, 95) <= input(11);
output(1, 96) <= input(63);
output(1, 97) <= input(61);
output(1, 98) <= input(33);
output(1, 99) <= input(16);
output(1, 100) <= input(46);
output(1, 101) <= input(47);
output(1, 102) <= input(48);
output(1, 103) <= input(49);
output(1, 104) <= input(50);
output(1, 105) <= input(51);
output(1, 106) <= input(52);
output(1, 107) <= input(23);
output(1, 108) <= input(24);
output(1, 109) <= input(25);
output(1, 110) <= input(26);
output(1, 111) <= input(27);
output(1, 112) <= input(64);
output(1, 113) <= input(62);
output(1, 114) <= input(60);
output(1, 115) <= input(32);
output(1, 116) <= input(0);
output(1, 117) <= input(53);
output(1, 118) <= input(54);
output(1, 119) <= input(55);
output(1, 120) <= input(56);
output(1, 121) <= input(57);
output(1, 122) <= input(58);
output(1, 123) <= input(59);
output(1, 124) <= input(7);
output(1, 125) <= input(8);
output(1, 126) <= input(9);
output(1, 127) <= input(10);
output(1, 128) <= input(65);
output(1, 129) <= input(64);
output(1, 130) <= input(62);
output(1, 131) <= input(60);
output(1, 132) <= input(32);
output(1, 133) <= input(0);
output(1, 134) <= input(53);
output(1, 135) <= input(54);
output(1, 136) <= input(55);
output(1, 137) <= input(56);
output(1, 138) <= input(57);
output(1, 139) <= input(58);
output(1, 140) <= input(59);
output(1, 141) <= input(7);
output(1, 142) <= input(8);
output(1, 143) <= input(9);
output(1, 144) <= input(66);
output(1, 145) <= input(67);
output(1, 146) <= input(63);
output(1, 147) <= input(61);
output(1, 148) <= input(33);
output(1, 149) <= input(16);
output(1, 150) <= input(46);
output(1, 151) <= input(47);
output(1, 152) <= input(48);
output(1, 153) <= input(49);
output(1, 154) <= input(50);
output(1, 155) <= input(51);
output(1, 156) <= input(52);
output(1, 157) <= input(23);
output(1, 158) <= input(24);
output(1, 159) <= input(25);
output(1, 160) <= input(68);
output(1, 161) <= input(65);
output(1, 162) <= input(64);
output(1, 163) <= input(62);
output(1, 164) <= input(60);
output(1, 165) <= input(32);
output(1, 166) <= input(0);
output(1, 167) <= input(53);
output(1, 168) <= input(54);
output(1, 169) <= input(55);
output(1, 170) <= input(56);
output(1, 171) <= input(57);
output(1, 172) <= input(58);
output(1, 173) <= input(59);
output(1, 174) <= input(7);
output(1, 175) <= input(8);
output(1, 176) <= input(69);
output(1, 177) <= input(66);
output(1, 178) <= input(67);
output(1, 179) <= input(63);
output(1, 180) <= input(61);
output(1, 181) <= input(33);
output(1, 182) <= input(16);
output(1, 183) <= input(46);
output(1, 184) <= input(47);
output(1, 185) <= input(48);
output(1, 186) <= input(49);
output(1, 187) <= input(50);
output(1, 188) <= input(51);
output(1, 189) <= input(52);
output(1, 190) <= input(23);
output(1, 191) <= input(24);
output(1, 192) <= input(70);
output(1, 193) <= input(68);
output(1, 194) <= input(65);
output(1, 195) <= input(64);
output(1, 196) <= input(62);
output(1, 197) <= input(60);
output(1, 198) <= input(32);
output(1, 199) <= input(0);
output(1, 200) <= input(53);
output(1, 201) <= input(54);
output(1, 202) <= input(55);
output(1, 203) <= input(56);
output(1, 204) <= input(57);
output(1, 205) <= input(58);
output(1, 206) <= input(59);
output(1, 207) <= input(7);
output(1, 208) <= input(71);
output(1, 209) <= input(69);
output(1, 210) <= input(66);
output(1, 211) <= input(67);
output(1, 212) <= input(63);
output(1, 213) <= input(61);
output(1, 214) <= input(33);
output(1, 215) <= input(16);
output(1, 216) <= input(46);
output(1, 217) <= input(47);
output(1, 218) <= input(48);
output(1, 219) <= input(49);
output(1, 220) <= input(50);
output(1, 221) <= input(51);
output(1, 222) <= input(52);
output(1, 223) <= input(23);
output(1, 224) <= input(72);
output(1, 225) <= input(70);
output(1, 226) <= input(68);
output(1, 227) <= input(65);
output(1, 228) <= input(64);
output(1, 229) <= input(62);
output(1, 230) <= input(60);
output(1, 231) <= input(32);
output(1, 232) <= input(0);
output(1, 233) <= input(53);
output(1, 234) <= input(54);
output(1, 235) <= input(55);
output(1, 236) <= input(56);
output(1, 237) <= input(57);
output(1, 238) <= input(58);
output(1, 239) <= input(59);
output(1, 240) <= input(73);
output(1, 241) <= input(71);
output(1, 242) <= input(69);
output(1, 243) <= input(66);
output(1, 244) <= input(67);
output(1, 245) <= input(63);
output(1, 246) <= input(61);
output(1, 247) <= input(33);
output(1, 248) <= input(16);
output(1, 249) <= input(46);
output(1, 250) <= input(47);
output(1, 251) <= input(48);
output(1, 252) <= input(49);
output(1, 253) <= input(50);
output(1, 254) <= input(51);
output(1, 255) <= input(52);
when "0110" =>
output(0, 0) <= input(0);
output(0, 1) <= input(1);
output(0, 2) <= input(2);
output(0, 3) <= input(3);
output(0, 4) <= input(4);
output(0, 5) <= input(5);
output(0, 6) <= input(6);
output(0, 7) <= input(7);
output(0, 8) <= input(8);
output(0, 9) <= input(9);
output(0, 10) <= input(10);
output(0, 11) <= input(11);
output(0, 12) <= input(12);
output(0, 13) <= input(13);
output(0, 14) <= input(14);
output(0, 15) <= input(15);
output(0, 16) <= input(16);
output(0, 17) <= input(17);
output(0, 18) <= input(18);
output(0, 19) <= input(19);
output(0, 20) <= input(20);
output(0, 21) <= input(21);
output(0, 22) <= input(22);
output(0, 23) <= input(23);
output(0, 24) <= input(24);
output(0, 25) <= input(25);
output(0, 26) <= input(26);
output(0, 27) <= input(27);
output(0, 28) <= input(28);
output(0, 29) <= input(29);
output(0, 30) <= input(30);
output(0, 31) <= input(31);
output(0, 32) <= input(32);
output(0, 33) <= input(0);
output(0, 34) <= input(1);
output(0, 35) <= input(2);
output(0, 36) <= input(3);
output(0, 37) <= input(4);
output(0, 38) <= input(5);
output(0, 39) <= input(6);
output(0, 40) <= input(7);
output(0, 41) <= input(8);
output(0, 42) <= input(9);
output(0, 43) <= input(10);
output(0, 44) <= input(11);
output(0, 45) <= input(12);
output(0, 46) <= input(13);
output(0, 47) <= input(14);
output(0, 48) <= input(33);
output(0, 49) <= input(16);
output(0, 50) <= input(17);
output(0, 51) <= input(18);
output(0, 52) <= input(19);
output(0, 53) <= input(20);
output(0, 54) <= input(21);
output(0, 55) <= input(22);
output(0, 56) <= input(23);
output(0, 57) <= input(24);
output(0, 58) <= input(25);
output(0, 59) <= input(26);
output(0, 60) <= input(27);
output(0, 61) <= input(28);
output(0, 62) <= input(29);
output(0, 63) <= input(30);
output(0, 64) <= input(34);
output(0, 65) <= input(33);
output(0, 66) <= input(16);
output(0, 67) <= input(17);
output(0, 68) <= input(18);
output(0, 69) <= input(19);
output(0, 70) <= input(20);
output(0, 71) <= input(21);
output(0, 72) <= input(22);
output(0, 73) <= input(23);
output(0, 74) <= input(24);
output(0, 75) <= input(25);
output(0, 76) <= input(26);
output(0, 77) <= input(27);
output(0, 78) <= input(28);
output(0, 79) <= input(29);
output(0, 80) <= input(35);
output(0, 81) <= input(36);
output(0, 82) <= input(32);
output(0, 83) <= input(0);
output(0, 84) <= input(1);
output(0, 85) <= input(2);
output(0, 86) <= input(3);
output(0, 87) <= input(4);
output(0, 88) <= input(5);
output(0, 89) <= input(6);
output(0, 90) <= input(7);
output(0, 91) <= input(8);
output(0, 92) <= input(9);
output(0, 93) <= input(10);
output(0, 94) <= input(11);
output(0, 95) <= input(12);
output(0, 96) <= input(37);
output(0, 97) <= input(34);
output(0, 98) <= input(33);
output(0, 99) <= input(16);
output(0, 100) <= input(17);
output(0, 101) <= input(18);
output(0, 102) <= input(19);
output(0, 103) <= input(20);
output(0, 104) <= input(21);
output(0, 105) <= input(22);
output(0, 106) <= input(23);
output(0, 107) <= input(24);
output(0, 108) <= input(25);
output(0, 109) <= input(26);
output(0, 110) <= input(27);
output(0, 111) <= input(28);
output(0, 112) <= input(38);
output(0, 113) <= input(35);
output(0, 114) <= input(36);
output(0, 115) <= input(32);
output(0, 116) <= input(0);
output(0, 117) <= input(1);
output(0, 118) <= input(2);
output(0, 119) <= input(3);
output(0, 120) <= input(4);
output(0, 121) <= input(5);
output(0, 122) <= input(6);
output(0, 123) <= input(7);
output(0, 124) <= input(8);
output(0, 125) <= input(9);
output(0, 126) <= input(10);
output(0, 127) <= input(11);
output(0, 128) <= input(39);
output(0, 129) <= input(38);
output(0, 130) <= input(35);
output(0, 131) <= input(36);
output(0, 132) <= input(32);
output(0, 133) <= input(0);
output(0, 134) <= input(1);
output(0, 135) <= input(2);
output(0, 136) <= input(3);
output(0, 137) <= input(4);
output(0, 138) <= input(5);
output(0, 139) <= input(6);
output(0, 140) <= input(7);
output(0, 141) <= input(8);
output(0, 142) <= input(9);
output(0, 143) <= input(10);
output(0, 144) <= input(40);
output(0, 145) <= input(41);
output(0, 146) <= input(37);
output(0, 147) <= input(34);
output(0, 148) <= input(33);
output(0, 149) <= input(16);
output(0, 150) <= input(17);
output(0, 151) <= input(18);
output(0, 152) <= input(19);
output(0, 153) <= input(20);
output(0, 154) <= input(21);
output(0, 155) <= input(22);
output(0, 156) <= input(23);
output(0, 157) <= input(24);
output(0, 158) <= input(25);
output(0, 159) <= input(26);
output(0, 160) <= input(42);
output(0, 161) <= input(39);
output(0, 162) <= input(38);
output(0, 163) <= input(35);
output(0, 164) <= input(36);
output(0, 165) <= input(32);
output(0, 166) <= input(0);
output(0, 167) <= input(1);
output(0, 168) <= input(2);
output(0, 169) <= input(3);
output(0, 170) <= input(4);
output(0, 171) <= input(5);
output(0, 172) <= input(6);
output(0, 173) <= input(7);
output(0, 174) <= input(8);
output(0, 175) <= input(9);
output(0, 176) <= input(43);
output(0, 177) <= input(40);
output(0, 178) <= input(41);
output(0, 179) <= input(37);
output(0, 180) <= input(34);
output(0, 181) <= input(33);
output(0, 182) <= input(16);
output(0, 183) <= input(17);
output(0, 184) <= input(18);
output(0, 185) <= input(19);
output(0, 186) <= input(20);
output(0, 187) <= input(21);
output(0, 188) <= input(22);
output(0, 189) <= input(23);
output(0, 190) <= input(24);
output(0, 191) <= input(25);
output(0, 192) <= input(44);
output(0, 193) <= input(43);
output(0, 194) <= input(40);
output(0, 195) <= input(41);
output(0, 196) <= input(37);
output(0, 197) <= input(34);
output(0, 198) <= input(33);
output(0, 199) <= input(16);
output(0, 200) <= input(17);
output(0, 201) <= input(18);
output(0, 202) <= input(19);
output(0, 203) <= input(20);
output(0, 204) <= input(21);
output(0, 205) <= input(22);
output(0, 206) <= input(23);
output(0, 207) <= input(24);
output(0, 208) <= input(45);
output(0, 209) <= input(46);
output(0, 210) <= input(42);
output(0, 211) <= input(39);
output(0, 212) <= input(38);
output(0, 213) <= input(35);
output(0, 214) <= input(36);
output(0, 215) <= input(32);
output(0, 216) <= input(0);
output(0, 217) <= input(1);
output(0, 218) <= input(2);
output(0, 219) <= input(3);
output(0, 220) <= input(4);
output(0, 221) <= input(5);
output(0, 222) <= input(6);
output(0, 223) <= input(7);
output(0, 224) <= input(47);
output(0, 225) <= input(44);
output(0, 226) <= input(43);
output(0, 227) <= input(40);
output(0, 228) <= input(41);
output(0, 229) <= input(37);
output(0, 230) <= input(34);
output(0, 231) <= input(33);
output(0, 232) <= input(16);
output(0, 233) <= input(17);
output(0, 234) <= input(18);
output(0, 235) <= input(19);
output(0, 236) <= input(20);
output(0, 237) <= input(21);
output(0, 238) <= input(22);
output(0, 239) <= input(23);
output(0, 240) <= input(48);
output(0, 241) <= input(45);
output(0, 242) <= input(46);
output(0, 243) <= input(42);
output(0, 244) <= input(39);
output(0, 245) <= input(38);
output(0, 246) <= input(35);
output(0, 247) <= input(36);
output(0, 248) <= input(32);
output(0, 249) <= input(0);
output(0, 250) <= input(1);
output(0, 251) <= input(2);
output(0, 252) <= input(3);
output(0, 253) <= input(4);
output(0, 254) <= input(5);
output(0, 255) <= input(6);
output(1, 0) <= input(49);
output(1, 1) <= input(50);
output(1, 2) <= input(51);
output(1, 3) <= input(19);
output(1, 4) <= input(20);
output(1, 5) <= input(52);
output(1, 6) <= input(53);
output(1, 7) <= input(54);
output(1, 8) <= input(55);
output(1, 9) <= input(56);
output(1, 10) <= input(57);
output(1, 11) <= input(58);
output(1, 12) <= input(59);
output(1, 13) <= input(28);
output(1, 14) <= input(29);
output(1, 15) <= input(30);
output(1, 16) <= input(60);
output(1, 17) <= input(61);
output(1, 18) <= input(62);
output(1, 19) <= input(2);
output(1, 20) <= input(3);
output(1, 21) <= input(63);
output(1, 22) <= input(64);
output(1, 23) <= input(65);
output(1, 24) <= input(66);
output(1, 25) <= input(67);
output(1, 26) <= input(68);
output(1, 27) <= input(69);
output(1, 28) <= input(70);
output(1, 29) <= input(11);
output(1, 30) <= input(12);
output(1, 31) <= input(13);
output(1, 32) <= input(71);
output(1, 33) <= input(60);
output(1, 34) <= input(61);
output(1, 35) <= input(62);
output(1, 36) <= input(2);
output(1, 37) <= input(3);
output(1, 38) <= input(63);
output(1, 39) <= input(64);
output(1, 40) <= input(65);
output(1, 41) <= input(66);
output(1, 42) <= input(67);
output(1, 43) <= input(68);
output(1, 44) <= input(69);
output(1, 45) <= input(70);
output(1, 46) <= input(11);
output(1, 47) <= input(12);
output(1, 48) <= input(72);
output(1, 49) <= input(73);
output(1, 50) <= input(49);
output(1, 51) <= input(50);
output(1, 52) <= input(51);
output(1, 53) <= input(19);
output(1, 54) <= input(20);
output(1, 55) <= input(52);
output(1, 56) <= input(53);
output(1, 57) <= input(54);
output(1, 58) <= input(55);
output(1, 59) <= input(56);
output(1, 60) <= input(57);
output(1, 61) <= input(58);
output(1, 62) <= input(59);
output(1, 63) <= input(28);
output(1, 64) <= input(34);
output(1, 65) <= input(72);
output(1, 66) <= input(73);
output(1, 67) <= input(49);
output(1, 68) <= input(50);
output(1, 69) <= input(51);
output(1, 70) <= input(19);
output(1, 71) <= input(20);
output(1, 72) <= input(52);
output(1, 73) <= input(53);
output(1, 74) <= input(54);
output(1, 75) <= input(55);
output(1, 76) <= input(56);
output(1, 77) <= input(57);
output(1, 78) <= input(58);
output(1, 79) <= input(59);
output(1, 80) <= input(35);
output(1, 81) <= input(74);
output(1, 82) <= input(71);
output(1, 83) <= input(60);
output(1, 84) <= input(61);
output(1, 85) <= input(62);
output(1, 86) <= input(2);
output(1, 87) <= input(3);
output(1, 88) <= input(63);
output(1, 89) <= input(64);
output(1, 90) <= input(65);
output(1, 91) <= input(66);
output(1, 92) <= input(67);
output(1, 93) <= input(68);
output(1, 94) <= input(69);
output(1, 95) <= input(70);
output(1, 96) <= input(38);
output(1, 97) <= input(35);
output(1, 98) <= input(74);
output(1, 99) <= input(71);
output(1, 100) <= input(60);
output(1, 101) <= input(61);
output(1, 102) <= input(62);
output(1, 103) <= input(2);
output(1, 104) <= input(3);
output(1, 105) <= input(63);
output(1, 106) <= input(64);
output(1, 107) <= input(65);
output(1, 108) <= input(66);
output(1, 109) <= input(67);
output(1, 110) <= input(68);
output(1, 111) <= input(69);
output(1, 112) <= input(75);
output(1, 113) <= input(37);
output(1, 114) <= input(34);
output(1, 115) <= input(72);
output(1, 116) <= input(73);
output(1, 117) <= input(49);
output(1, 118) <= input(50);
output(1, 119) <= input(51);
output(1, 120) <= input(19);
output(1, 121) <= input(20);
output(1, 122) <= input(52);
output(1, 123) <= input(53);
output(1, 124) <= input(54);
output(1, 125) <= input(55);
output(1, 126) <= input(56);
output(1, 127) <= input(57);
output(1, 128) <= input(76);
output(1, 129) <= input(38);
output(1, 130) <= input(35);
output(1, 131) <= input(74);
output(1, 132) <= input(71);
output(1, 133) <= input(60);
output(1, 134) <= input(61);
output(1, 135) <= input(62);
output(1, 136) <= input(2);
output(1, 137) <= input(3);
output(1, 138) <= input(63);
output(1, 139) <= input(64);
output(1, 140) <= input(65);
output(1, 141) <= input(66);
output(1, 142) <= input(67);
output(1, 143) <= input(68);
output(1, 144) <= input(77);
output(1, 145) <= input(76);
output(1, 146) <= input(38);
output(1, 147) <= input(35);
output(1, 148) <= input(74);
output(1, 149) <= input(71);
output(1, 150) <= input(60);
output(1, 151) <= input(61);
output(1, 152) <= input(62);
output(1, 153) <= input(2);
output(1, 154) <= input(3);
output(1, 155) <= input(63);
output(1, 156) <= input(64);
output(1, 157) <= input(65);
output(1, 158) <= input(66);
output(1, 159) <= input(67);
output(1, 160) <= input(78);
output(1, 161) <= input(79);
output(1, 162) <= input(75);
output(1, 163) <= input(37);
output(1, 164) <= input(34);
output(1, 165) <= input(72);
output(1, 166) <= input(73);
output(1, 167) <= input(49);
output(1, 168) <= input(50);
output(1, 169) <= input(51);
output(1, 170) <= input(19);
output(1, 171) <= input(20);
output(1, 172) <= input(52);
output(1, 173) <= input(53);
output(1, 174) <= input(54);
output(1, 175) <= input(55);
output(1, 176) <= input(80);
output(1, 177) <= input(78);
output(1, 178) <= input(79);
output(1, 179) <= input(75);
output(1, 180) <= input(37);
output(1, 181) <= input(34);
output(1, 182) <= input(72);
output(1, 183) <= input(73);
output(1, 184) <= input(49);
output(1, 185) <= input(50);
output(1, 186) <= input(51);
output(1, 187) <= input(19);
output(1, 188) <= input(20);
output(1, 189) <= input(52);
output(1, 190) <= input(53);
output(1, 191) <= input(54);
output(1, 192) <= input(81);
output(1, 193) <= input(82);
output(1, 194) <= input(77);
output(1, 195) <= input(76);
output(1, 196) <= input(38);
output(1, 197) <= input(35);
output(1, 198) <= input(74);
output(1, 199) <= input(71);
output(1, 200) <= input(60);
output(1, 201) <= input(61);
output(1, 202) <= input(62);
output(1, 203) <= input(2);
output(1, 204) <= input(3);
output(1, 205) <= input(63);
output(1, 206) <= input(64);
output(1, 207) <= input(65);
output(1, 208) <= input(83);
output(1, 209) <= input(81);
output(1, 210) <= input(82);
output(1, 211) <= input(77);
output(1, 212) <= input(76);
output(1, 213) <= input(38);
output(1, 214) <= input(35);
output(1, 215) <= input(74);
output(1, 216) <= input(71);
output(1, 217) <= input(60);
output(1, 218) <= input(61);
output(1, 219) <= input(62);
output(1, 220) <= input(2);
output(1, 221) <= input(3);
output(1, 222) <= input(63);
output(1, 223) <= input(64);
output(1, 224) <= input(84);
output(1, 225) <= input(85);
output(1, 226) <= input(80);
output(1, 227) <= input(78);
output(1, 228) <= input(79);
output(1, 229) <= input(75);
output(1, 230) <= input(37);
output(1, 231) <= input(34);
output(1, 232) <= input(72);
output(1, 233) <= input(73);
output(1, 234) <= input(49);
output(1, 235) <= input(50);
output(1, 236) <= input(51);
output(1, 237) <= input(19);
output(1, 238) <= input(20);
output(1, 239) <= input(52);
output(1, 240) <= input(86);
output(1, 241) <= input(83);
output(1, 242) <= input(81);
output(1, 243) <= input(82);
output(1, 244) <= input(77);
output(1, 245) <= input(76);
output(1, 246) <= input(38);
output(1, 247) <= input(35);
output(1, 248) <= input(74);
output(1, 249) <= input(71);
output(1, 250) <= input(60);
output(1, 251) <= input(61);
output(1, 252) <= input(62);
output(1, 253) <= input(2);
output(1, 254) <= input(3);
output(1, 255) <= input(63);
output(2, 0) <= input(87);
output(2, 1) <= input(88);
output(2, 2) <= input(89);
output(2, 3) <= input(90);
output(2, 4) <= input(91);
output(2, 5) <= input(92);
output(2, 6) <= input(93);
output(2, 7) <= input(94);
output(2, 8) <= input(95);
output(2, 9) <= input(96);
output(2, 10) <= input(97);
output(2, 11) <= input(98);
output(2, 12) <= input(99);
output(2, 13) <= input(70);
output(2, 14) <= input(11);
output(2, 15) <= input(12);
output(2, 16) <= input(100);
output(2, 17) <= input(87);
output(2, 18) <= input(88);
output(2, 19) <= input(89);
output(2, 20) <= input(90);
output(2, 21) <= input(91);
output(2, 22) <= input(92);
output(2, 23) <= input(93);
output(2, 24) <= input(94);
output(2, 25) <= input(95);
output(2, 26) <= input(96);
output(2, 27) <= input(97);
output(2, 28) <= input(98);
output(2, 29) <= input(99);
output(2, 30) <= input(70);
output(2, 31) <= input(11);
output(2, 32) <= input(101);
output(2, 33) <= input(102);
output(2, 34) <= input(103);
output(2, 35) <= input(104);
output(2, 36) <= input(105);
output(2, 37) <= input(106);
output(2, 38) <= input(107);
output(2, 39) <= input(108);
output(2, 40) <= input(109);
output(2, 41) <= input(110);
output(2, 42) <= input(111);
output(2, 43) <= input(112);
output(2, 44) <= input(113);
output(2, 45) <= input(114);
output(2, 46) <= input(115);
output(2, 47) <= input(59);
output(2, 48) <= input(116);
output(2, 49) <= input(101);
output(2, 50) <= input(102);
output(2, 51) <= input(103);
output(2, 52) <= input(104);
output(2, 53) <= input(105);
output(2, 54) <= input(106);
output(2, 55) <= input(107);
output(2, 56) <= input(108);
output(2, 57) <= input(109);
output(2, 58) <= input(110);
output(2, 59) <= input(111);
output(2, 60) <= input(112);
output(2, 61) <= input(113);
output(2, 62) <= input(114);
output(2, 63) <= input(115);
output(2, 64) <= input(117);
output(2, 65) <= input(116);
output(2, 66) <= input(101);
output(2, 67) <= input(102);
output(2, 68) <= input(103);
output(2, 69) <= input(104);
output(2, 70) <= input(105);
output(2, 71) <= input(106);
output(2, 72) <= input(107);
output(2, 73) <= input(108);
output(2, 74) <= input(109);
output(2, 75) <= input(110);
output(2, 76) <= input(111);
output(2, 77) <= input(112);
output(2, 78) <= input(113);
output(2, 79) <= input(114);
output(2, 80) <= input(118);
output(2, 81) <= input(119);
output(2, 82) <= input(120);
output(2, 83) <= input(100);
output(2, 84) <= input(87);
output(2, 85) <= input(88);
output(2, 86) <= input(89);
output(2, 87) <= input(90);
output(2, 88) <= input(91);
output(2, 89) <= input(92);
output(2, 90) <= input(93);
output(2, 91) <= input(94);
output(2, 92) <= input(95);
output(2, 93) <= input(96);
output(2, 94) <= input(97);
output(2, 95) <= input(98);
output(2, 96) <= input(121);
output(2, 97) <= input(118);
output(2, 98) <= input(119);
output(2, 99) <= input(120);
output(2, 100) <= input(100);
output(2, 101) <= input(87);
output(2, 102) <= input(88);
output(2, 103) <= input(89);
output(2, 104) <= input(90);
output(2, 105) <= input(91);
output(2, 106) <= input(92);
output(2, 107) <= input(93);
output(2, 108) <= input(94);
output(2, 109) <= input(95);
output(2, 110) <= input(96);
output(2, 111) <= input(97);
output(2, 112) <= input(122);
output(2, 113) <= input(123);
output(2, 114) <= input(117);
output(2, 115) <= input(116);
output(2, 116) <= input(101);
output(2, 117) <= input(102);
output(2, 118) <= input(103);
output(2, 119) <= input(104);
output(2, 120) <= input(105);
output(2, 121) <= input(106);
output(2, 122) <= input(107);
output(2, 123) <= input(108);
output(2, 124) <= input(109);
output(2, 125) <= input(110);
output(2, 126) <= input(111);
output(2, 127) <= input(112);
output(2, 128) <= input(124);
output(2, 129) <= input(122);
output(2, 130) <= input(123);
output(2, 131) <= input(117);
output(2, 132) <= input(116);
output(2, 133) <= input(101);
output(2, 134) <= input(102);
output(2, 135) <= input(103);
output(2, 136) <= input(104);
output(2, 137) <= input(105);
output(2, 138) <= input(106);
output(2, 139) <= input(107);
output(2, 140) <= input(108);
output(2, 141) <= input(109);
output(2, 142) <= input(110);
output(2, 143) <= input(111);
output(2, 144) <= input(125);
output(2, 145) <= input(124);
output(2, 146) <= input(122);
output(2, 147) <= input(123);
output(2, 148) <= input(117);
output(2, 149) <= input(116);
output(2, 150) <= input(101);
output(2, 151) <= input(102);
output(2, 152) <= input(103);
output(2, 153) <= input(104);
output(2, 154) <= input(105);
output(2, 155) <= input(106);
output(2, 156) <= input(107);
output(2, 157) <= input(108);
output(2, 158) <= input(109);
output(2, 159) <= input(110);
output(2, 160) <= input(126);
output(2, 161) <= input(127);
output(2, 162) <= input(128);
output(2, 163) <= input(121);
output(2, 164) <= input(118);
output(2, 165) <= input(119);
output(2, 166) <= input(120);
output(2, 167) <= input(100);
output(2, 168) <= input(87);
output(2, 169) <= input(88);
output(2, 170) <= input(89);
output(2, 171) <= input(90);
output(2, 172) <= input(91);
output(2, 173) <= input(92);
output(2, 174) <= input(93);
output(2, 175) <= input(94);
output(2, 176) <= input(129);
output(2, 177) <= input(126);
output(2, 178) <= input(127);
output(2, 179) <= input(128);
output(2, 180) <= input(121);
output(2, 181) <= input(118);
output(2, 182) <= input(119);
output(2, 183) <= input(120);
output(2, 184) <= input(100);
output(2, 185) <= input(87);
output(2, 186) <= input(88);
output(2, 187) <= input(89);
output(2, 188) <= input(90);
output(2, 189) <= input(91);
output(2, 190) <= input(92);
output(2, 191) <= input(93);
output(2, 192) <= input(130);
output(2, 193) <= input(129);
output(2, 194) <= input(126);
output(2, 195) <= input(127);
output(2, 196) <= input(128);
output(2, 197) <= input(121);
output(2, 198) <= input(118);
output(2, 199) <= input(119);
output(2, 200) <= input(120);
output(2, 201) <= input(100);
output(2, 202) <= input(87);
output(2, 203) <= input(88);
output(2, 204) <= input(89);
output(2, 205) <= input(90);
output(2, 206) <= input(91);
output(2, 207) <= input(92);
output(2, 208) <= input(131);
output(2, 209) <= input(132);
output(2, 210) <= input(133);
output(2, 211) <= input(125);
output(2, 212) <= input(124);
output(2, 213) <= input(122);
output(2, 214) <= input(123);
output(2, 215) <= input(117);
output(2, 216) <= input(116);
output(2, 217) <= input(101);
output(2, 218) <= input(102);
output(2, 219) <= input(103);
output(2, 220) <= input(104);
output(2, 221) <= input(105);
output(2, 222) <= input(106);
output(2, 223) <= input(107);
output(2, 224) <= input(134);
output(2, 225) <= input(131);
output(2, 226) <= input(132);
output(2, 227) <= input(133);
output(2, 228) <= input(125);
output(2, 229) <= input(124);
output(2, 230) <= input(122);
output(2, 231) <= input(123);
output(2, 232) <= input(117);
output(2, 233) <= input(116);
output(2, 234) <= input(101);
output(2, 235) <= input(102);
output(2, 236) <= input(103);
output(2, 237) <= input(104);
output(2, 238) <= input(105);
output(2, 239) <= input(106);
output(2, 240) <= input(135);
output(2, 241) <= input(136);
output(2, 242) <= input(130);
output(2, 243) <= input(129);
output(2, 244) <= input(126);
output(2, 245) <= input(127);
output(2, 246) <= input(128);
output(2, 247) <= input(121);
output(2, 248) <= input(118);
output(2, 249) <= input(119);
output(2, 250) <= input(120);
output(2, 251) <= input(100);
output(2, 252) <= input(87);
output(2, 253) <= input(88);
output(2, 254) <= input(89);
output(2, 255) <= input(90);
when "0111" =>
output(0, 0) <= input(0);
output(0, 1) <= input(1);
output(0, 2) <= input(2);
output(0, 3) <= input(3);
output(0, 4) <= input(4);
output(0, 5) <= input(5);
output(0, 6) <= input(6);
output(0, 7) <= input(7);
output(0, 8) <= input(8);
output(0, 9) <= input(9);
output(0, 10) <= input(10);
output(0, 11) <= input(11);
output(0, 12) <= input(12);
output(0, 13) <= input(13);
output(0, 14) <= input(14);
output(0, 15) <= input(15);
output(0, 16) <= input(16);
output(0, 17) <= input(0);
output(0, 18) <= input(1);
output(0, 19) <= input(2);
output(0, 20) <= input(3);
output(0, 21) <= input(4);
output(0, 22) <= input(5);
output(0, 23) <= input(6);
output(0, 24) <= input(7);
output(0, 25) <= input(8);
output(0, 26) <= input(9);
output(0, 27) <= input(10);
output(0, 28) <= input(11);
output(0, 29) <= input(12);
output(0, 30) <= input(13);
output(0, 31) <= input(14);
output(0, 32) <= input(17);
output(0, 33) <= input(16);
output(0, 34) <= input(0);
output(0, 35) <= input(1);
output(0, 36) <= input(2);
output(0, 37) <= input(3);
output(0, 38) <= input(4);
output(0, 39) <= input(5);
output(0, 40) <= input(6);
output(0, 41) <= input(7);
output(0, 42) <= input(8);
output(0, 43) <= input(9);
output(0, 44) <= input(10);
output(0, 45) <= input(11);
output(0, 46) <= input(12);
output(0, 47) <= input(13);
output(0, 48) <= input(18);
output(0, 49) <= input(17);
output(0, 50) <= input(16);
output(0, 51) <= input(0);
output(0, 52) <= input(1);
output(0, 53) <= input(2);
output(0, 54) <= input(3);
output(0, 55) <= input(4);
output(0, 56) <= input(5);
output(0, 57) <= input(6);
output(0, 58) <= input(7);
output(0, 59) <= input(8);
output(0, 60) <= input(9);
output(0, 61) <= input(10);
output(0, 62) <= input(11);
output(0, 63) <= input(12);
output(0, 64) <= input(19);
output(0, 65) <= input(18);
output(0, 66) <= input(17);
output(0, 67) <= input(16);
output(0, 68) <= input(0);
output(0, 69) <= input(1);
output(0, 70) <= input(2);
output(0, 71) <= input(3);
output(0, 72) <= input(4);
output(0, 73) <= input(5);
output(0, 74) <= input(6);
output(0, 75) <= input(7);
output(0, 76) <= input(8);
output(0, 77) <= input(9);
output(0, 78) <= input(10);
output(0, 79) <= input(11);
output(0, 80) <= input(20);
output(0, 81) <= input(21);
output(0, 82) <= input(22);
output(0, 83) <= input(23);
output(0, 84) <= input(24);
output(0, 85) <= input(25);
output(0, 86) <= input(26);
output(0, 87) <= input(27);
output(0, 88) <= input(28);
output(0, 89) <= input(29);
output(0, 90) <= input(30);
output(0, 91) <= input(31);
output(0, 92) <= input(32);
output(0, 93) <= input(33);
output(0, 94) <= input(34);
output(0, 95) <= input(35);
output(0, 96) <= input(36);
output(0, 97) <= input(20);
output(0, 98) <= input(21);
output(0, 99) <= input(22);
output(0, 100) <= input(23);
output(0, 101) <= input(24);
output(0, 102) <= input(25);
output(0, 103) <= input(26);
output(0, 104) <= input(27);
output(0, 105) <= input(28);
output(0, 106) <= input(29);
output(0, 107) <= input(30);
output(0, 108) <= input(31);
output(0, 109) <= input(32);
output(0, 110) <= input(33);
output(0, 111) <= input(34);
output(0, 112) <= input(37);
output(0, 113) <= input(36);
output(0, 114) <= input(20);
output(0, 115) <= input(21);
output(0, 116) <= input(22);
output(0, 117) <= input(23);
output(0, 118) <= input(24);
output(0, 119) <= input(25);
output(0, 120) <= input(26);
output(0, 121) <= input(27);
output(0, 122) <= input(28);
output(0, 123) <= input(29);
output(0, 124) <= input(30);
output(0, 125) <= input(31);
output(0, 126) <= input(32);
output(0, 127) <= input(33);
output(0, 128) <= input(38);
output(0, 129) <= input(37);
output(0, 130) <= input(36);
output(0, 131) <= input(20);
output(0, 132) <= input(21);
output(0, 133) <= input(22);
output(0, 134) <= input(23);
output(0, 135) <= input(24);
output(0, 136) <= input(25);
output(0, 137) <= input(26);
output(0, 138) <= input(27);
output(0, 139) <= input(28);
output(0, 140) <= input(29);
output(0, 141) <= input(30);
output(0, 142) <= input(31);
output(0, 143) <= input(32);
output(0, 144) <= input(39);
output(0, 145) <= input(38);
output(0, 146) <= input(37);
output(0, 147) <= input(36);
output(0, 148) <= input(20);
output(0, 149) <= input(21);
output(0, 150) <= input(22);
output(0, 151) <= input(23);
output(0, 152) <= input(24);
output(0, 153) <= input(25);
output(0, 154) <= input(26);
output(0, 155) <= input(27);
output(0, 156) <= input(28);
output(0, 157) <= input(29);
output(0, 158) <= input(30);
output(0, 159) <= input(31);
output(0, 160) <= input(40);
output(0, 161) <= input(41);
output(0, 162) <= input(42);
output(0, 163) <= input(43);
output(0, 164) <= input(44);
output(0, 165) <= input(19);
output(0, 166) <= input(18);
output(0, 167) <= input(17);
output(0, 168) <= input(16);
output(0, 169) <= input(0);
output(0, 170) <= input(1);
output(0, 171) <= input(2);
output(0, 172) <= input(3);
output(0, 173) <= input(4);
output(0, 174) <= input(5);
output(0, 175) <= input(6);
output(0, 176) <= input(45);
output(0, 177) <= input(40);
output(0, 178) <= input(41);
output(0, 179) <= input(42);
output(0, 180) <= input(43);
output(0, 181) <= input(44);
output(0, 182) <= input(19);
output(0, 183) <= input(18);
output(0, 184) <= input(17);
output(0, 185) <= input(16);
output(0, 186) <= input(0);
output(0, 187) <= input(1);
output(0, 188) <= input(2);
output(0, 189) <= input(3);
output(0, 190) <= input(4);
output(0, 191) <= input(5);
output(0, 192) <= input(46);
output(0, 193) <= input(45);
output(0, 194) <= input(40);
output(0, 195) <= input(41);
output(0, 196) <= input(42);
output(0, 197) <= input(43);
output(0, 198) <= input(44);
output(0, 199) <= input(19);
output(0, 200) <= input(18);
output(0, 201) <= input(17);
output(0, 202) <= input(16);
output(0, 203) <= input(0);
output(0, 204) <= input(1);
output(0, 205) <= input(2);
output(0, 206) <= input(3);
output(0, 207) <= input(4);
output(0, 208) <= input(47);
output(0, 209) <= input(46);
output(0, 210) <= input(45);
output(0, 211) <= input(40);
output(0, 212) <= input(41);
output(0, 213) <= input(42);
output(0, 214) <= input(43);
output(0, 215) <= input(44);
output(0, 216) <= input(19);
output(0, 217) <= input(18);
output(0, 218) <= input(17);
output(0, 219) <= input(16);
output(0, 220) <= input(0);
output(0, 221) <= input(1);
output(0, 222) <= input(2);
output(0, 223) <= input(3);
output(0, 224) <= input(48);
output(0, 225) <= input(47);
output(0, 226) <= input(46);
output(0, 227) <= input(45);
output(0, 228) <= input(40);
output(0, 229) <= input(41);
output(0, 230) <= input(42);
output(0, 231) <= input(43);
output(0, 232) <= input(44);
output(0, 233) <= input(19);
output(0, 234) <= input(18);
output(0, 235) <= input(17);
output(0, 236) <= input(16);
output(0, 237) <= input(0);
output(0, 238) <= input(1);
output(0, 239) <= input(2);
output(0, 240) <= input(49);
output(0, 241) <= input(50);
output(0, 242) <= input(51);
output(0, 243) <= input(52);
output(0, 244) <= input(53);
output(0, 245) <= input(39);
output(0, 246) <= input(38);
output(0, 247) <= input(37);
output(0, 248) <= input(36);
output(0, 249) <= input(20);
output(0, 250) <= input(21);
output(0, 251) <= input(22);
output(0, 252) <= input(23);
output(0, 253) <= input(24);
output(0, 254) <= input(25);
output(0, 255) <= input(26);
output(1, 0) <= input(54);
output(1, 1) <= input(55);
output(1, 2) <= input(56);
output(1, 3) <= input(57);
output(1, 4) <= input(58);
output(1, 5) <= input(59);
output(1, 6) <= input(60);
output(1, 7) <= input(61);
output(1, 8) <= input(62);
output(1, 9) <= input(63);
output(1, 10) <= input(64);
output(1, 11) <= input(65);
output(1, 12) <= input(66);
output(1, 13) <= input(67);
output(1, 14) <= input(68);
output(1, 15) <= input(69);
output(1, 16) <= input(70);
output(1, 17) <= input(54);
output(1, 18) <= input(55);
output(1, 19) <= input(56);
output(1, 20) <= input(57);
output(1, 21) <= input(58);
output(1, 22) <= input(59);
output(1, 23) <= input(60);
output(1, 24) <= input(61);
output(1, 25) <= input(62);
output(1, 26) <= input(63);
output(1, 27) <= input(64);
output(1, 28) <= input(65);
output(1, 29) <= input(66);
output(1, 30) <= input(67);
output(1, 31) <= input(68);
output(1, 32) <= input(71);
output(1, 33) <= input(70);
output(1, 34) <= input(54);
output(1, 35) <= input(55);
output(1, 36) <= input(56);
output(1, 37) <= input(57);
output(1, 38) <= input(58);
output(1, 39) <= input(59);
output(1, 40) <= input(60);
output(1, 41) <= input(61);
output(1, 42) <= input(62);
output(1, 43) <= input(63);
output(1, 44) <= input(64);
output(1, 45) <= input(65);
output(1, 46) <= input(66);
output(1, 47) <= input(67);
output(1, 48) <= input(72);
output(1, 49) <= input(71);
output(1, 50) <= input(70);
output(1, 51) <= input(54);
output(1, 52) <= input(55);
output(1, 53) <= input(56);
output(1, 54) <= input(57);
output(1, 55) <= input(58);
output(1, 56) <= input(59);
output(1, 57) <= input(60);
output(1, 58) <= input(61);
output(1, 59) <= input(62);
output(1, 60) <= input(63);
output(1, 61) <= input(64);
output(1, 62) <= input(65);
output(1, 63) <= input(66);
output(1, 64) <= input(73);
output(1, 65) <= input(72);
output(1, 66) <= input(71);
output(1, 67) <= input(70);
output(1, 68) <= input(54);
output(1, 69) <= input(55);
output(1, 70) <= input(56);
output(1, 71) <= input(57);
output(1, 72) <= input(58);
output(1, 73) <= input(59);
output(1, 74) <= input(60);
output(1, 75) <= input(61);
output(1, 76) <= input(62);
output(1, 77) <= input(63);
output(1, 78) <= input(64);
output(1, 79) <= input(65);
output(1, 80) <= input(74);
output(1, 81) <= input(73);
output(1, 82) <= input(72);
output(1, 83) <= input(71);
output(1, 84) <= input(70);
output(1, 85) <= input(54);
output(1, 86) <= input(55);
output(1, 87) <= input(56);
output(1, 88) <= input(57);
output(1, 89) <= input(58);
output(1, 90) <= input(59);
output(1, 91) <= input(60);
output(1, 92) <= input(61);
output(1, 93) <= input(62);
output(1, 94) <= input(63);
output(1, 95) <= input(64);
output(1, 96) <= input(75);
output(1, 97) <= input(74);
output(1, 98) <= input(73);
output(1, 99) <= input(72);
output(1, 100) <= input(71);
output(1, 101) <= input(70);
output(1, 102) <= input(54);
output(1, 103) <= input(55);
output(1, 104) <= input(56);
output(1, 105) <= input(57);
output(1, 106) <= input(58);
output(1, 107) <= input(59);
output(1, 108) <= input(60);
output(1, 109) <= input(61);
output(1, 110) <= input(62);
output(1, 111) <= input(63);
output(1, 112) <= input(76);
output(1, 113) <= input(75);
output(1, 114) <= input(74);
output(1, 115) <= input(73);
output(1, 116) <= input(72);
output(1, 117) <= input(71);
output(1, 118) <= input(70);
output(1, 119) <= input(54);
output(1, 120) <= input(55);
output(1, 121) <= input(56);
output(1, 122) <= input(57);
output(1, 123) <= input(58);
output(1, 124) <= input(59);
output(1, 125) <= input(60);
output(1, 126) <= input(61);
output(1, 127) <= input(62);
output(1, 128) <= input(77);
output(1, 129) <= input(76);
output(1, 130) <= input(75);
output(1, 131) <= input(74);
output(1, 132) <= input(73);
output(1, 133) <= input(72);
output(1, 134) <= input(71);
output(1, 135) <= input(70);
output(1, 136) <= input(54);
output(1, 137) <= input(55);
output(1, 138) <= input(56);
output(1, 139) <= input(57);
output(1, 140) <= input(58);
output(1, 141) <= input(59);
output(1, 142) <= input(60);
output(1, 143) <= input(61);
output(1, 144) <= input(78);
output(1, 145) <= input(77);
output(1, 146) <= input(76);
output(1, 147) <= input(75);
output(1, 148) <= input(74);
output(1, 149) <= input(73);
output(1, 150) <= input(72);
output(1, 151) <= input(71);
output(1, 152) <= input(70);
output(1, 153) <= input(54);
output(1, 154) <= input(55);
output(1, 155) <= input(56);
output(1, 156) <= input(57);
output(1, 157) <= input(58);
output(1, 158) <= input(59);
output(1, 159) <= input(60);
output(1, 160) <= input(79);
output(1, 161) <= input(78);
output(1, 162) <= input(77);
output(1, 163) <= input(76);
output(1, 164) <= input(75);
output(1, 165) <= input(74);
output(1, 166) <= input(73);
output(1, 167) <= input(72);
output(1, 168) <= input(71);
output(1, 169) <= input(70);
output(1, 170) <= input(54);
output(1, 171) <= input(55);
output(1, 172) <= input(56);
output(1, 173) <= input(57);
output(1, 174) <= input(58);
output(1, 175) <= input(59);
output(1, 176) <= input(80);
output(1, 177) <= input(79);
output(1, 178) <= input(78);
output(1, 179) <= input(77);
output(1, 180) <= input(76);
output(1, 181) <= input(75);
output(1, 182) <= input(74);
output(1, 183) <= input(73);
output(1, 184) <= input(72);
output(1, 185) <= input(71);
output(1, 186) <= input(70);
output(1, 187) <= input(54);
output(1, 188) <= input(55);
output(1, 189) <= input(56);
output(1, 190) <= input(57);
output(1, 191) <= input(58);
output(1, 192) <= input(81);
output(1, 193) <= input(80);
output(1, 194) <= input(79);
output(1, 195) <= input(78);
output(1, 196) <= input(77);
output(1, 197) <= input(76);
output(1, 198) <= input(75);
output(1, 199) <= input(74);
output(1, 200) <= input(73);
output(1, 201) <= input(72);
output(1, 202) <= input(71);
output(1, 203) <= input(70);
output(1, 204) <= input(54);
output(1, 205) <= input(55);
output(1, 206) <= input(56);
output(1, 207) <= input(57);
output(1, 208) <= input(82);
output(1, 209) <= input(81);
output(1, 210) <= input(80);
output(1, 211) <= input(79);
output(1, 212) <= input(78);
output(1, 213) <= input(77);
output(1, 214) <= input(76);
output(1, 215) <= input(75);
output(1, 216) <= input(74);
output(1, 217) <= input(73);
output(1, 218) <= input(72);
output(1, 219) <= input(71);
output(1, 220) <= input(70);
output(1, 221) <= input(54);
output(1, 222) <= input(55);
output(1, 223) <= input(56);
output(1, 224) <= input(83);
output(1, 225) <= input(82);
output(1, 226) <= input(81);
output(1, 227) <= input(80);
output(1, 228) <= input(79);
output(1, 229) <= input(78);
output(1, 230) <= input(77);
output(1, 231) <= input(76);
output(1, 232) <= input(75);
output(1, 233) <= input(74);
output(1, 234) <= input(73);
output(1, 235) <= input(72);
output(1, 236) <= input(71);
output(1, 237) <= input(70);
output(1, 238) <= input(54);
output(1, 239) <= input(55);
output(1, 240) <= input(84);
output(1, 241) <= input(83);
output(1, 242) <= input(82);
output(1, 243) <= input(81);
output(1, 244) <= input(80);
output(1, 245) <= input(79);
output(1, 246) <= input(78);
output(1, 247) <= input(77);
output(1, 248) <= input(76);
output(1, 249) <= input(75);
output(1, 250) <= input(74);
output(1, 251) <= input(73);
output(1, 252) <= input(72);
output(1, 253) <= input(71);
output(1, 254) <= input(70);
output(1, 255) <= input(54);
when "1000" =>
output(0, 0) <= input(0);
output(0, 1) <= input(1);
output(0, 2) <= input(2);
output(0, 3) <= input(3);
output(0, 4) <= input(4);
output(0, 5) <= input(5);
output(0, 6) <= input(6);
output(0, 7) <= input(7);
output(0, 8) <= input(8);
output(0, 9) <= input(9);
output(0, 10) <= input(10);
output(0, 11) <= input(11);
output(0, 12) <= input(12);
output(0, 13) <= input(13);
output(0, 14) <= input(14);
output(0, 15) <= input(15);
output(0, 16) <= input(16);
output(0, 17) <= input(0);
output(0, 18) <= input(1);
output(0, 19) <= input(2);
output(0, 20) <= input(3);
output(0, 21) <= input(4);
output(0, 22) <= input(5);
output(0, 23) <= input(6);
output(0, 24) <= input(7);
output(0, 25) <= input(8);
output(0, 26) <= input(9);
output(0, 27) <= input(10);
output(0, 28) <= input(11);
output(0, 29) <= input(12);
output(0, 30) <= input(13);
output(0, 31) <= input(14);
output(0, 32) <= input(17);
output(0, 33) <= input(16);
output(0, 34) <= input(0);
output(0, 35) <= input(1);
output(0, 36) <= input(2);
output(0, 37) <= input(3);
output(0, 38) <= input(4);
output(0, 39) <= input(5);
output(0, 40) <= input(6);
output(0, 41) <= input(7);
output(0, 42) <= input(8);
output(0, 43) <= input(9);
output(0, 44) <= input(10);
output(0, 45) <= input(11);
output(0, 46) <= input(12);
output(0, 47) <= input(13);
output(0, 48) <= input(18);
output(0, 49) <= input(17);
output(0, 50) <= input(16);
output(0, 51) <= input(0);
output(0, 52) <= input(1);
output(0, 53) <= input(2);
output(0, 54) <= input(3);
output(0, 55) <= input(4);
output(0, 56) <= input(5);
output(0, 57) <= input(6);
output(0, 58) <= input(7);
output(0, 59) <= input(8);
output(0, 60) <= input(9);
output(0, 61) <= input(10);
output(0, 62) <= input(11);
output(0, 63) <= input(12);
output(0, 64) <= input(19);
output(0, 65) <= input(18);
output(0, 66) <= input(17);
output(0, 67) <= input(16);
output(0, 68) <= input(0);
output(0, 69) <= input(1);
output(0, 70) <= input(2);
output(0, 71) <= input(3);
output(0, 72) <= input(4);
output(0, 73) <= input(5);
output(0, 74) <= input(6);
output(0, 75) <= input(7);
output(0, 76) <= input(8);
output(0, 77) <= input(9);
output(0, 78) <= input(10);
output(0, 79) <= input(11);
output(0, 80) <= input(20);
output(0, 81) <= input(21);
output(0, 82) <= input(22);
output(0, 83) <= input(23);
output(0, 84) <= input(24);
output(0, 85) <= input(25);
output(0, 86) <= input(26);
output(0, 87) <= input(27);
output(0, 88) <= input(28);
output(0, 89) <= input(29);
output(0, 90) <= input(30);
output(0, 91) <= input(31);
output(0, 92) <= input(32);
output(0, 93) <= input(33);
output(0, 94) <= input(34);
output(0, 95) <= input(35);
output(0, 96) <= input(36);
output(0, 97) <= input(20);
output(0, 98) <= input(21);
output(0, 99) <= input(22);
output(0, 100) <= input(23);
output(0, 101) <= input(24);
output(0, 102) <= input(25);
output(0, 103) <= input(26);
output(0, 104) <= input(27);
output(0, 105) <= input(28);
output(0, 106) <= input(29);
output(0, 107) <= input(30);
output(0, 108) <= input(31);
output(0, 109) <= input(32);
output(0, 110) <= input(33);
output(0, 111) <= input(34);
output(0, 112) <= input(37);
output(0, 113) <= input(36);
output(0, 114) <= input(20);
output(0, 115) <= input(21);
output(0, 116) <= input(22);
output(0, 117) <= input(23);
output(0, 118) <= input(24);
output(0, 119) <= input(25);
output(0, 120) <= input(26);
output(0, 121) <= input(27);
output(0, 122) <= input(28);
output(0, 123) <= input(29);
output(0, 124) <= input(30);
output(0, 125) <= input(31);
output(0, 126) <= input(32);
output(0, 127) <= input(33);
output(0, 128) <= input(38);
output(0, 129) <= input(37);
output(0, 130) <= input(36);
output(0, 131) <= input(20);
output(0, 132) <= input(21);
output(0, 133) <= input(22);
output(0, 134) <= input(23);
output(0, 135) <= input(24);
output(0, 136) <= input(25);
output(0, 137) <= input(26);
output(0, 138) <= input(27);
output(0, 139) <= input(28);
output(0, 140) <= input(29);
output(0, 141) <= input(30);
output(0, 142) <= input(31);
output(0, 143) <= input(32);
output(0, 144) <= input(39);
output(0, 145) <= input(38);
output(0, 146) <= input(37);
output(0, 147) <= input(36);
output(0, 148) <= input(20);
output(0, 149) <= input(21);
output(0, 150) <= input(22);
output(0, 151) <= input(23);
output(0, 152) <= input(24);
output(0, 153) <= input(25);
output(0, 154) <= input(26);
output(0, 155) <= input(27);
output(0, 156) <= input(28);
output(0, 157) <= input(29);
output(0, 158) <= input(30);
output(0, 159) <= input(31);
output(0, 160) <= input(40);
output(0, 161) <= input(41);
output(0, 162) <= input(42);
output(0, 163) <= input(43);
output(0, 164) <= input(44);
output(0, 165) <= input(19);
output(0, 166) <= input(18);
output(0, 167) <= input(17);
output(0, 168) <= input(16);
output(0, 169) <= input(0);
output(0, 170) <= input(1);
output(0, 171) <= input(2);
output(0, 172) <= input(3);
output(0, 173) <= input(4);
output(0, 174) <= input(5);
output(0, 175) <= input(6);
output(0, 176) <= input(45);
output(0, 177) <= input(40);
output(0, 178) <= input(41);
output(0, 179) <= input(42);
output(0, 180) <= input(43);
output(0, 181) <= input(44);
output(0, 182) <= input(19);
output(0, 183) <= input(18);
output(0, 184) <= input(17);
output(0, 185) <= input(16);
output(0, 186) <= input(0);
output(0, 187) <= input(1);
output(0, 188) <= input(2);
output(0, 189) <= input(3);
output(0, 190) <= input(4);
output(0, 191) <= input(5);
output(0, 192) <= input(46);
output(0, 193) <= input(45);
output(0, 194) <= input(40);
output(0, 195) <= input(41);
output(0, 196) <= input(42);
output(0, 197) <= input(43);
output(0, 198) <= input(44);
output(0, 199) <= input(19);
output(0, 200) <= input(18);
output(0, 201) <= input(17);
output(0, 202) <= input(16);
output(0, 203) <= input(0);
output(0, 204) <= input(1);
output(0, 205) <= input(2);
output(0, 206) <= input(3);
output(0, 207) <= input(4);
output(0, 208) <= input(47);
output(0, 209) <= input(46);
output(0, 210) <= input(45);
output(0, 211) <= input(40);
output(0, 212) <= input(41);
output(0, 213) <= input(42);
output(0, 214) <= input(43);
output(0, 215) <= input(44);
output(0, 216) <= input(19);
output(0, 217) <= input(18);
output(0, 218) <= input(17);
output(0, 219) <= input(16);
output(0, 220) <= input(0);
output(0, 221) <= input(1);
output(0, 222) <= input(2);
output(0, 223) <= input(3);
output(0, 224) <= input(48);
output(0, 225) <= input(47);
output(0, 226) <= input(46);
output(0, 227) <= input(45);
output(0, 228) <= input(40);
output(0, 229) <= input(41);
output(0, 230) <= input(42);
output(0, 231) <= input(43);
output(0, 232) <= input(44);
output(0, 233) <= input(19);
output(0, 234) <= input(18);
output(0, 235) <= input(17);
output(0, 236) <= input(16);
output(0, 237) <= input(0);
output(0, 238) <= input(1);
output(0, 239) <= input(2);
output(0, 240) <= input(49);
output(0, 241) <= input(50);
output(0, 242) <= input(51);
output(0, 243) <= input(52);
output(0, 244) <= input(53);
output(0, 245) <= input(39);
output(0, 246) <= input(38);
output(0, 247) <= input(37);
output(0, 248) <= input(36);
output(0, 249) <= input(20);
output(0, 250) <= input(21);
output(0, 251) <= input(22);
output(0, 252) <= input(23);
output(0, 253) <= input(24);
output(0, 254) <= input(25);
output(0, 255) <= input(26);
when "1001" =>
output(0, 0) <= input(0);
output(0, 1) <= input(1);
output(0, 2) <= input(2);
output(0, 3) <= input(3);
output(0, 4) <= input(4);
output(0, 5) <= input(5);
output(0, 6) <= input(6);
output(0, 7) <= input(7);
output(0, 8) <= input(8);
output(0, 9) <= input(9);
output(0, 10) <= input(10);
output(0, 11) <= input(11);
output(0, 12) <= input(12);
output(0, 13) <= input(13);
output(0, 14) <= input(14);
output(0, 15) <= input(15);
output(0, 16) <= input(16);
output(0, 17) <= input(0);
output(0, 18) <= input(1);
output(0, 19) <= input(2);
output(0, 20) <= input(3);
output(0, 21) <= input(4);
output(0, 22) <= input(5);
output(0, 23) <= input(6);
output(0, 24) <= input(7);
output(0, 25) <= input(8);
output(0, 26) <= input(9);
output(0, 27) <= input(10);
output(0, 28) <= input(11);
output(0, 29) <= input(12);
output(0, 30) <= input(13);
output(0, 31) <= input(14);
output(0, 32) <= input(17);
output(0, 33) <= input(18);
output(0, 34) <= input(19);
output(0, 35) <= input(20);
output(0, 36) <= input(21);
output(0, 37) <= input(22);
output(0, 38) <= input(23);
output(0, 39) <= input(24);
output(0, 40) <= input(25);
output(0, 41) <= input(26);
output(0, 42) <= input(27);
output(0, 43) <= input(28);
output(0, 44) <= input(29);
output(0, 45) <= input(30);
output(0, 46) <= input(31);
output(0, 47) <= input(32);
output(0, 48) <= input(33);
output(0, 49) <= input(17);
output(0, 50) <= input(18);
output(0, 51) <= input(19);
output(0, 52) <= input(20);
output(0, 53) <= input(21);
output(0, 54) <= input(22);
output(0, 55) <= input(23);
output(0, 56) <= input(24);
output(0, 57) <= input(25);
output(0, 58) <= input(26);
output(0, 59) <= input(27);
output(0, 60) <= input(28);
output(0, 61) <= input(29);
output(0, 62) <= input(30);
output(0, 63) <= input(31);
output(0, 64) <= input(34);
output(0, 65) <= input(33);
output(0, 66) <= input(17);
output(0, 67) <= input(18);
output(0, 68) <= input(19);
output(0, 69) <= input(20);
output(0, 70) <= input(21);
output(0, 71) <= input(22);
output(0, 72) <= input(23);
output(0, 73) <= input(24);
output(0, 74) <= input(25);
output(0, 75) <= input(26);
output(0, 76) <= input(27);
output(0, 77) <= input(28);
output(0, 78) <= input(29);
output(0, 79) <= input(30);
output(0, 80) <= input(35);
output(0, 81) <= input(36);
output(0, 82) <= input(37);
output(0, 83) <= input(16);
output(0, 84) <= input(0);
output(0, 85) <= input(1);
output(0, 86) <= input(2);
output(0, 87) <= input(3);
output(0, 88) <= input(4);
output(0, 89) <= input(5);
output(0, 90) <= input(6);
output(0, 91) <= input(7);
output(0, 92) <= input(8);
output(0, 93) <= input(9);
output(0, 94) <= input(10);
output(0, 95) <= input(11);
output(0, 96) <= input(38);
output(0, 97) <= input(35);
output(0, 98) <= input(36);
output(0, 99) <= input(37);
output(0, 100) <= input(16);
output(0, 101) <= input(0);
output(0, 102) <= input(1);
output(0, 103) <= input(2);
output(0, 104) <= input(3);
output(0, 105) <= input(4);
output(0, 106) <= input(5);
output(0, 107) <= input(6);
output(0, 108) <= input(7);
output(0, 109) <= input(8);
output(0, 110) <= input(9);
output(0, 111) <= input(10);
output(0, 112) <= input(39);
output(0, 113) <= input(40);
output(0, 114) <= input(34);
output(0, 115) <= input(33);
output(0, 116) <= input(17);
output(0, 117) <= input(18);
output(0, 118) <= input(19);
output(0, 119) <= input(20);
output(0, 120) <= input(21);
output(0, 121) <= input(22);
output(0, 122) <= input(23);
output(0, 123) <= input(24);
output(0, 124) <= input(25);
output(0, 125) <= input(26);
output(0, 126) <= input(27);
output(0, 127) <= input(28);
output(0, 128) <= input(41);
output(0, 129) <= input(39);
output(0, 130) <= input(40);
output(0, 131) <= input(34);
output(0, 132) <= input(33);
output(0, 133) <= input(17);
output(0, 134) <= input(18);
output(0, 135) <= input(19);
output(0, 136) <= input(20);
output(0, 137) <= input(21);
output(0, 138) <= input(22);
output(0, 139) <= input(23);
output(0, 140) <= input(24);
output(0, 141) <= input(25);
output(0, 142) <= input(26);
output(0, 143) <= input(27);
output(0, 144) <= input(42);
output(0, 145) <= input(41);
output(0, 146) <= input(39);
output(0, 147) <= input(40);
output(0, 148) <= input(34);
output(0, 149) <= input(33);
output(0, 150) <= input(17);
output(0, 151) <= input(18);
output(0, 152) <= input(19);
output(0, 153) <= input(20);
output(0, 154) <= input(21);
output(0, 155) <= input(22);
output(0, 156) <= input(23);
output(0, 157) <= input(24);
output(0, 158) <= input(25);
output(0, 159) <= input(26);
output(0, 160) <= input(43);
output(0, 161) <= input(44);
output(0, 162) <= input(45);
output(0, 163) <= input(38);
output(0, 164) <= input(35);
output(0, 165) <= input(36);
output(0, 166) <= input(37);
output(0, 167) <= input(16);
output(0, 168) <= input(0);
output(0, 169) <= input(1);
output(0, 170) <= input(2);
output(0, 171) <= input(3);
output(0, 172) <= input(4);
output(0, 173) <= input(5);
output(0, 174) <= input(6);
output(0, 175) <= input(7);
output(0, 176) <= input(46);
output(0, 177) <= input(43);
output(0, 178) <= input(44);
output(0, 179) <= input(45);
output(0, 180) <= input(38);
output(0, 181) <= input(35);
output(0, 182) <= input(36);
output(0, 183) <= input(37);
output(0, 184) <= input(16);
output(0, 185) <= input(0);
output(0, 186) <= input(1);
output(0, 187) <= input(2);
output(0, 188) <= input(3);
output(0, 189) <= input(4);
output(0, 190) <= input(5);
output(0, 191) <= input(6);
output(0, 192) <= input(47);
output(0, 193) <= input(46);
output(0, 194) <= input(43);
output(0, 195) <= input(44);
output(0, 196) <= input(45);
output(0, 197) <= input(38);
output(0, 198) <= input(35);
output(0, 199) <= input(36);
output(0, 200) <= input(37);
output(0, 201) <= input(16);
output(0, 202) <= input(0);
output(0, 203) <= input(1);
output(0, 204) <= input(2);
output(0, 205) <= input(3);
output(0, 206) <= input(4);
output(0, 207) <= input(5);
output(0, 208) <= input(48);
output(0, 209) <= input(49);
output(0, 210) <= input(50);
output(0, 211) <= input(42);
output(0, 212) <= input(41);
output(0, 213) <= input(39);
output(0, 214) <= input(40);
output(0, 215) <= input(34);
output(0, 216) <= input(33);
output(0, 217) <= input(17);
output(0, 218) <= input(18);
output(0, 219) <= input(19);
output(0, 220) <= input(20);
output(0, 221) <= input(21);
output(0, 222) <= input(22);
output(0, 223) <= input(23);
output(0, 224) <= input(51);
output(0, 225) <= input(48);
output(0, 226) <= input(49);
output(0, 227) <= input(50);
output(0, 228) <= input(42);
output(0, 229) <= input(41);
output(0, 230) <= input(39);
output(0, 231) <= input(40);
output(0, 232) <= input(34);
output(0, 233) <= input(33);
output(0, 234) <= input(17);
output(0, 235) <= input(18);
output(0, 236) <= input(19);
output(0, 237) <= input(20);
output(0, 238) <= input(21);
output(0, 239) <= input(22);
output(0, 240) <= input(52);
output(0, 241) <= input(53);
output(0, 242) <= input(47);
output(0, 243) <= input(46);
output(0, 244) <= input(43);
output(0, 245) <= input(44);
output(0, 246) <= input(45);
output(0, 247) <= input(38);
output(0, 248) <= input(35);
output(0, 249) <= input(36);
output(0, 250) <= input(37);
output(0, 251) <= input(16);
output(0, 252) <= input(0);
output(0, 253) <= input(1);
output(0, 254) <= input(2);
output(0, 255) <= input(3);
output(1, 0) <= input(54);
output(1, 1) <= input(55);
output(1, 2) <= input(56);
output(1, 3) <= input(57);
output(1, 4) <= input(58);
output(1, 5) <= input(59);
output(1, 6) <= input(60);
output(1, 7) <= input(61);
output(1, 8) <= input(62);
output(1, 9) <= input(63);
output(1, 10) <= input(64);
output(1, 11) <= input(65);
output(1, 12) <= input(32);
output(1, 13) <= input(66);
output(1, 14) <= input(67);
output(1, 15) <= input(68);
output(1, 16) <= input(69);
output(1, 17) <= input(70);
output(1, 18) <= input(71);
output(1, 19) <= input(72);
output(1, 20) <= input(73);
output(1, 21) <= input(74);
output(1, 22) <= input(75);
output(1, 23) <= input(76);
output(1, 24) <= input(77);
output(1, 25) <= input(78);
output(1, 26) <= input(79);
output(1, 27) <= input(80);
output(1, 28) <= input(13);
output(1, 29) <= input(14);
output(1, 30) <= input(15);
output(1, 31) <= input(81);
output(1, 32) <= input(82);
output(1, 33) <= input(69);
output(1, 34) <= input(70);
output(1, 35) <= input(71);
output(1, 36) <= input(72);
output(1, 37) <= input(73);
output(1, 38) <= input(74);
output(1, 39) <= input(75);
output(1, 40) <= input(76);
output(1, 41) <= input(77);
output(1, 42) <= input(78);
output(1, 43) <= input(79);
output(1, 44) <= input(80);
output(1, 45) <= input(13);
output(1, 46) <= input(14);
output(1, 47) <= input(15);
output(1, 48) <= input(83);
output(1, 49) <= input(84);
output(1, 50) <= input(54);
output(1, 51) <= input(55);
output(1, 52) <= input(56);
output(1, 53) <= input(57);
output(1, 54) <= input(58);
output(1, 55) <= input(59);
output(1, 56) <= input(60);
output(1, 57) <= input(61);
output(1, 58) <= input(62);
output(1, 59) <= input(63);
output(1, 60) <= input(64);
output(1, 61) <= input(65);
output(1, 62) <= input(32);
output(1, 63) <= input(66);
output(1, 64) <= input(85);
output(1, 65) <= input(83);
output(1, 66) <= input(84);
output(1, 67) <= input(54);
output(1, 68) <= input(55);
output(1, 69) <= input(56);
output(1, 70) <= input(57);
output(1, 71) <= input(58);
output(1, 72) <= input(59);
output(1, 73) <= input(60);
output(1, 74) <= input(61);
output(1, 75) <= input(62);
output(1, 76) <= input(63);
output(1, 77) <= input(64);
output(1, 78) <= input(65);
output(1, 79) <= input(32);
output(1, 80) <= input(86);
output(1, 81) <= input(87);
output(1, 82) <= input(82);
output(1, 83) <= input(69);
output(1, 84) <= input(70);
output(1, 85) <= input(71);
output(1, 86) <= input(72);
output(1, 87) <= input(73);
output(1, 88) <= input(74);
output(1, 89) <= input(75);
output(1, 90) <= input(76);
output(1, 91) <= input(77);
output(1, 92) <= input(78);
output(1, 93) <= input(79);
output(1, 94) <= input(80);
output(1, 95) <= input(13);
output(1, 96) <= input(88);
output(1, 97) <= input(86);
output(1, 98) <= input(87);
output(1, 99) <= input(82);
output(1, 100) <= input(69);
output(1, 101) <= input(70);
output(1, 102) <= input(71);
output(1, 103) <= input(72);
output(1, 104) <= input(73);
output(1, 105) <= input(74);
output(1, 106) <= input(75);
output(1, 107) <= input(76);
output(1, 108) <= input(77);
output(1, 109) <= input(78);
output(1, 110) <= input(79);
output(1, 111) <= input(80);
output(1, 112) <= input(89);
output(1, 113) <= input(90);
output(1, 114) <= input(85);
output(1, 115) <= input(83);
output(1, 116) <= input(84);
output(1, 117) <= input(54);
output(1, 118) <= input(55);
output(1, 119) <= input(56);
output(1, 120) <= input(57);
output(1, 121) <= input(58);
output(1, 122) <= input(59);
output(1, 123) <= input(60);
output(1, 124) <= input(61);
output(1, 125) <= input(62);
output(1, 126) <= input(63);
output(1, 127) <= input(64);
output(1, 128) <= input(91);
output(1, 129) <= input(88);
output(1, 130) <= input(86);
output(1, 131) <= input(87);
output(1, 132) <= input(82);
output(1, 133) <= input(69);
output(1, 134) <= input(70);
output(1, 135) <= input(71);
output(1, 136) <= input(72);
output(1, 137) <= input(73);
output(1, 138) <= input(74);
output(1, 139) <= input(75);
output(1, 140) <= input(76);
output(1, 141) <= input(77);
output(1, 142) <= input(78);
output(1, 143) <= input(79);
output(1, 144) <= input(92);
output(1, 145) <= input(91);
output(1, 146) <= input(88);
output(1, 147) <= input(86);
output(1, 148) <= input(87);
output(1, 149) <= input(82);
output(1, 150) <= input(69);
output(1, 151) <= input(70);
output(1, 152) <= input(71);
output(1, 153) <= input(72);
output(1, 154) <= input(73);
output(1, 155) <= input(74);
output(1, 156) <= input(75);
output(1, 157) <= input(76);
output(1, 158) <= input(77);
output(1, 159) <= input(78);
output(1, 160) <= input(93);
output(1, 161) <= input(94);
output(1, 162) <= input(89);
output(1, 163) <= input(90);
output(1, 164) <= input(85);
output(1, 165) <= input(83);
output(1, 166) <= input(84);
output(1, 167) <= input(54);
output(1, 168) <= input(55);
output(1, 169) <= input(56);
output(1, 170) <= input(57);
output(1, 171) <= input(58);
output(1, 172) <= input(59);
output(1, 173) <= input(60);
output(1, 174) <= input(61);
output(1, 175) <= input(62);
output(1, 176) <= input(95);
output(1, 177) <= input(93);
output(1, 178) <= input(94);
output(1, 179) <= input(89);
output(1, 180) <= input(90);
output(1, 181) <= input(85);
output(1, 182) <= input(83);
output(1, 183) <= input(84);
output(1, 184) <= input(54);
output(1, 185) <= input(55);
output(1, 186) <= input(56);
output(1, 187) <= input(57);
output(1, 188) <= input(58);
output(1, 189) <= input(59);
output(1, 190) <= input(60);
output(1, 191) <= input(61);
output(1, 192) <= input(96);
output(1, 193) <= input(97);
output(1, 194) <= input(92);
output(1, 195) <= input(91);
output(1, 196) <= input(88);
output(1, 197) <= input(86);
output(1, 198) <= input(87);
output(1, 199) <= input(82);
output(1, 200) <= input(69);
output(1, 201) <= input(70);
output(1, 202) <= input(71);
output(1, 203) <= input(72);
output(1, 204) <= input(73);
output(1, 205) <= input(74);
output(1, 206) <= input(75);
output(1, 207) <= input(76);
output(1, 208) <= input(98);
output(1, 209) <= input(96);
output(1, 210) <= input(97);
output(1, 211) <= input(92);
output(1, 212) <= input(91);
output(1, 213) <= input(88);
output(1, 214) <= input(86);
output(1, 215) <= input(87);
output(1, 216) <= input(82);
output(1, 217) <= input(69);
output(1, 218) <= input(70);
output(1, 219) <= input(71);
output(1, 220) <= input(72);
output(1, 221) <= input(73);
output(1, 222) <= input(74);
output(1, 223) <= input(75);
output(1, 224) <= input(99);
output(1, 225) <= input(100);
output(1, 226) <= input(95);
output(1, 227) <= input(93);
output(1, 228) <= input(94);
output(1, 229) <= input(89);
output(1, 230) <= input(90);
output(1, 231) <= input(85);
output(1, 232) <= input(83);
output(1, 233) <= input(84);
output(1, 234) <= input(54);
output(1, 235) <= input(55);
output(1, 236) <= input(56);
output(1, 237) <= input(57);
output(1, 238) <= input(58);
output(1, 239) <= input(59);
output(1, 240) <= input(101);
output(1, 241) <= input(98);
output(1, 242) <= input(96);
output(1, 243) <= input(97);
output(1, 244) <= input(92);
output(1, 245) <= input(91);
output(1, 246) <= input(88);
output(1, 247) <= input(86);
output(1, 248) <= input(87);
output(1, 249) <= input(82);
output(1, 250) <= input(69);
output(1, 251) <= input(70);
output(1, 252) <= input(71);
output(1, 253) <= input(72);
output(1, 254) <= input(73);
output(1, 255) <= input(74);
output(2, 0) <= input(102);
output(2, 1) <= input(103);
output(2, 2) <= input(72);
output(2, 3) <= input(73);
output(2, 4) <= input(104);
output(2, 5) <= input(105);
output(2, 6) <= input(106);
output(2, 7) <= input(107);
output(2, 8) <= input(108);
output(2, 9) <= input(109);
output(2, 10) <= input(110);
output(2, 11) <= input(14);
output(2, 12) <= input(15);
output(2, 13) <= input(81);
output(2, 14) <= input(111);
output(2, 15) <= input(112);
output(2, 16) <= input(113);
output(2, 17) <= input(114);
output(2, 18) <= input(115);
output(2, 19) <= input(57);
output(2, 20) <= input(58);
output(2, 21) <= input(116);
output(2, 22) <= input(117);
output(2, 23) <= input(118);
output(2, 24) <= input(119);
output(2, 25) <= input(120);
output(2, 26) <= input(121);
output(2, 27) <= input(122);
output(2, 28) <= input(66);
output(2, 29) <= input(67);
output(2, 30) <= input(68);
output(2, 31) <= input(123);
output(2, 32) <= input(124);
output(2, 33) <= input(102);
output(2, 34) <= input(103);
output(2, 35) <= input(72);
output(2, 36) <= input(73);
output(2, 37) <= input(104);
output(2, 38) <= input(105);
output(2, 39) <= input(106);
output(2, 40) <= input(107);
output(2, 41) <= input(108);
output(2, 42) <= input(109);
output(2, 43) <= input(110);
output(2, 44) <= input(14);
output(2, 45) <= input(15);
output(2, 46) <= input(81);
output(2, 47) <= input(111);
output(2, 48) <= input(125);
output(2, 49) <= input(113);
output(2, 50) <= input(114);
output(2, 51) <= input(115);
output(2, 52) <= input(57);
output(2, 53) <= input(58);
output(2, 54) <= input(116);
output(2, 55) <= input(117);
output(2, 56) <= input(118);
output(2, 57) <= input(119);
output(2, 58) <= input(120);
output(2, 59) <= input(121);
output(2, 60) <= input(122);
output(2, 61) <= input(66);
output(2, 62) <= input(67);
output(2, 63) <= input(68);
output(2, 64) <= input(85);
output(2, 65) <= input(125);
output(2, 66) <= input(113);
output(2, 67) <= input(114);
output(2, 68) <= input(115);
output(2, 69) <= input(57);
output(2, 70) <= input(58);
output(2, 71) <= input(116);
output(2, 72) <= input(117);
output(2, 73) <= input(118);
output(2, 74) <= input(119);
output(2, 75) <= input(120);
output(2, 76) <= input(121);
output(2, 77) <= input(122);
output(2, 78) <= input(66);
output(2, 79) <= input(67);
output(2, 80) <= input(86);
output(2, 81) <= input(126);
output(2, 82) <= input(124);
output(2, 83) <= input(102);
output(2, 84) <= input(103);
output(2, 85) <= input(72);
output(2, 86) <= input(73);
output(2, 87) <= input(104);
output(2, 88) <= input(105);
output(2, 89) <= input(106);
output(2, 90) <= input(107);
output(2, 91) <= input(108);
output(2, 92) <= input(109);
output(2, 93) <= input(110);
output(2, 94) <= input(14);
output(2, 95) <= input(15);
output(2, 96) <= input(90);
output(2, 97) <= input(85);
output(2, 98) <= input(125);
output(2, 99) <= input(113);
output(2, 100) <= input(114);
output(2, 101) <= input(115);
output(2, 102) <= input(57);
output(2, 103) <= input(58);
output(2, 104) <= input(116);
output(2, 105) <= input(117);
output(2, 106) <= input(118);
output(2, 107) <= input(119);
output(2, 108) <= input(120);
output(2, 109) <= input(121);
output(2, 110) <= input(122);
output(2, 111) <= input(66);
output(2, 112) <= input(88);
output(2, 113) <= input(86);
output(2, 114) <= input(126);
output(2, 115) <= input(124);
output(2, 116) <= input(102);
output(2, 117) <= input(103);
output(2, 118) <= input(72);
output(2, 119) <= input(73);
output(2, 120) <= input(104);
output(2, 121) <= input(105);
output(2, 122) <= input(106);
output(2, 123) <= input(107);
output(2, 124) <= input(108);
output(2, 125) <= input(109);
output(2, 126) <= input(110);
output(2, 127) <= input(14);
output(2, 128) <= input(127);
output(2, 129) <= input(88);
output(2, 130) <= input(86);
output(2, 131) <= input(126);
output(2, 132) <= input(124);
output(2, 133) <= input(102);
output(2, 134) <= input(103);
output(2, 135) <= input(72);
output(2, 136) <= input(73);
output(2, 137) <= input(104);
output(2, 138) <= input(105);
output(2, 139) <= input(106);
output(2, 140) <= input(107);
output(2, 141) <= input(108);
output(2, 142) <= input(109);
output(2, 143) <= input(110);
output(2, 144) <= input(128);
output(2, 145) <= input(129);
output(2, 146) <= input(90);
output(2, 147) <= input(85);
output(2, 148) <= input(125);
output(2, 149) <= input(113);
output(2, 150) <= input(114);
output(2, 151) <= input(115);
output(2, 152) <= input(57);
output(2, 153) <= input(58);
output(2, 154) <= input(116);
output(2, 155) <= input(117);
output(2, 156) <= input(118);
output(2, 157) <= input(119);
output(2, 158) <= input(120);
output(2, 159) <= input(121);
output(2, 160) <= input(130);
output(2, 161) <= input(127);
output(2, 162) <= input(88);
output(2, 163) <= input(86);
output(2, 164) <= input(126);
output(2, 165) <= input(124);
output(2, 166) <= input(102);
output(2, 167) <= input(103);
output(2, 168) <= input(72);
output(2, 169) <= input(73);
output(2, 170) <= input(104);
output(2, 171) <= input(105);
output(2, 172) <= input(106);
output(2, 173) <= input(107);
output(2, 174) <= input(108);
output(2, 175) <= input(109);
output(2, 176) <= input(131);
output(2, 177) <= input(128);
output(2, 178) <= input(129);
output(2, 179) <= input(90);
output(2, 180) <= input(85);
output(2, 181) <= input(125);
output(2, 182) <= input(113);
output(2, 183) <= input(114);
output(2, 184) <= input(115);
output(2, 185) <= input(57);
output(2, 186) <= input(58);
output(2, 187) <= input(116);
output(2, 188) <= input(117);
output(2, 189) <= input(118);
output(2, 190) <= input(119);
output(2, 191) <= input(120);
output(2, 192) <= input(132);
output(2, 193) <= input(131);
output(2, 194) <= input(128);
output(2, 195) <= input(129);
output(2, 196) <= input(90);
output(2, 197) <= input(85);
output(2, 198) <= input(125);
output(2, 199) <= input(113);
output(2, 200) <= input(114);
output(2, 201) <= input(115);
output(2, 202) <= input(57);
output(2, 203) <= input(58);
output(2, 204) <= input(116);
output(2, 205) <= input(117);
output(2, 206) <= input(118);
output(2, 207) <= input(119);
output(2, 208) <= input(133);
output(2, 209) <= input(134);
output(2, 210) <= input(130);
output(2, 211) <= input(127);
output(2, 212) <= input(88);
output(2, 213) <= input(86);
output(2, 214) <= input(126);
output(2, 215) <= input(124);
output(2, 216) <= input(102);
output(2, 217) <= input(103);
output(2, 218) <= input(72);
output(2, 219) <= input(73);
output(2, 220) <= input(104);
output(2, 221) <= input(105);
output(2, 222) <= input(106);
output(2, 223) <= input(107);
output(2, 224) <= input(135);
output(2, 225) <= input(132);
output(2, 226) <= input(131);
output(2, 227) <= input(128);
output(2, 228) <= input(129);
output(2, 229) <= input(90);
output(2, 230) <= input(85);
output(2, 231) <= input(125);
output(2, 232) <= input(113);
output(2, 233) <= input(114);
output(2, 234) <= input(115);
output(2, 235) <= input(57);
output(2, 236) <= input(58);
output(2, 237) <= input(116);
output(2, 238) <= input(117);
output(2, 239) <= input(118);
output(2, 240) <= input(136);
output(2, 241) <= input(133);
output(2, 242) <= input(134);
output(2, 243) <= input(130);
output(2, 244) <= input(127);
output(2, 245) <= input(88);
output(2, 246) <= input(86);
output(2, 247) <= input(126);
output(2, 248) <= input(124);
output(2, 249) <= input(102);
output(2, 250) <= input(103);
output(2, 251) <= input(72);
output(2, 252) <= input(73);
output(2, 253) <= input(104);
output(2, 254) <= input(105);
output(2, 255) <= input(106);
when "1010" =>
output(0, 0) <= input(0);
output(0, 1) <= input(1);
output(0, 2) <= input(2);
output(0, 3) <= input(3);
output(0, 4) <= input(4);
output(0, 5) <= input(5);
output(0, 6) <= input(6);
output(0, 7) <= input(7);
output(0, 8) <= input(8);
output(0, 9) <= input(9);
output(0, 10) <= input(10);
output(0, 11) <= input(11);
output(0, 12) <= input(12);
output(0, 13) <= input(13);
output(0, 14) <= input(14);
output(0, 15) <= input(15);
output(0, 16) <= input(16);
output(0, 17) <= input(17);
output(0, 18) <= input(18);
output(0, 19) <= input(19);
output(0, 20) <= input(20);
output(0, 21) <= input(21);
output(0, 22) <= input(22);
output(0, 23) <= input(23);
output(0, 24) <= input(24);
output(0, 25) <= input(25);
output(0, 26) <= input(26);
output(0, 27) <= input(27);
output(0, 28) <= input(28);
output(0, 29) <= input(29);
output(0, 30) <= input(30);
output(0, 31) <= input(31);
output(0, 32) <= input(32);
output(0, 33) <= input(0);
output(0, 34) <= input(1);
output(0, 35) <= input(2);
output(0, 36) <= input(3);
output(0, 37) <= input(4);
output(0, 38) <= input(5);
output(0, 39) <= input(6);
output(0, 40) <= input(7);
output(0, 41) <= input(8);
output(0, 42) <= input(9);
output(0, 43) <= input(10);
output(0, 44) <= input(11);
output(0, 45) <= input(12);
output(0, 46) <= input(13);
output(0, 47) <= input(14);
output(0, 48) <= input(33);
output(0, 49) <= input(16);
output(0, 50) <= input(17);
output(0, 51) <= input(18);
output(0, 52) <= input(19);
output(0, 53) <= input(20);
output(0, 54) <= input(21);
output(0, 55) <= input(22);
output(0, 56) <= input(23);
output(0, 57) <= input(24);
output(0, 58) <= input(25);
output(0, 59) <= input(26);
output(0, 60) <= input(27);
output(0, 61) <= input(28);
output(0, 62) <= input(29);
output(0, 63) <= input(30);
output(0, 64) <= input(34);
output(0, 65) <= input(32);
output(0, 66) <= input(0);
output(0, 67) <= input(1);
output(0, 68) <= input(2);
output(0, 69) <= input(3);
output(0, 70) <= input(4);
output(0, 71) <= input(5);
output(0, 72) <= input(6);
output(0, 73) <= input(7);
output(0, 74) <= input(8);
output(0, 75) <= input(9);
output(0, 76) <= input(10);
output(0, 77) <= input(11);
output(0, 78) <= input(12);
output(0, 79) <= input(13);
output(0, 80) <= input(35);
output(0, 81) <= input(33);
output(0, 82) <= input(16);
output(0, 83) <= input(17);
output(0, 84) <= input(18);
output(0, 85) <= input(19);
output(0, 86) <= input(20);
output(0, 87) <= input(21);
output(0, 88) <= input(22);
output(0, 89) <= input(23);
output(0, 90) <= input(24);
output(0, 91) <= input(25);
output(0, 92) <= input(26);
output(0, 93) <= input(27);
output(0, 94) <= input(28);
output(0, 95) <= input(29);
output(0, 96) <= input(36);
output(0, 97) <= input(34);
output(0, 98) <= input(32);
output(0, 99) <= input(0);
output(0, 100) <= input(1);
output(0, 101) <= input(2);
output(0, 102) <= input(3);
output(0, 103) <= input(4);
output(0, 104) <= input(5);
output(0, 105) <= input(6);
output(0, 106) <= input(7);
output(0, 107) <= input(8);
output(0, 108) <= input(9);
output(0, 109) <= input(10);
output(0, 110) <= input(11);
output(0, 111) <= input(12);
output(0, 112) <= input(37);
output(0, 113) <= input(35);
output(0, 114) <= input(33);
output(0, 115) <= input(16);
output(0, 116) <= input(17);
output(0, 117) <= input(18);
output(0, 118) <= input(19);
output(0, 119) <= input(20);
output(0, 120) <= input(21);
output(0, 121) <= input(22);
output(0, 122) <= input(23);
output(0, 123) <= input(24);
output(0, 124) <= input(25);
output(0, 125) <= input(26);
output(0, 126) <= input(27);
output(0, 127) <= input(28);
output(0, 128) <= input(38);
output(0, 129) <= input(37);
output(0, 130) <= input(35);
output(0, 131) <= input(33);
output(0, 132) <= input(16);
output(0, 133) <= input(17);
output(0, 134) <= input(18);
output(0, 135) <= input(19);
output(0, 136) <= input(20);
output(0, 137) <= input(21);
output(0, 138) <= input(22);
output(0, 139) <= input(23);
output(0, 140) <= input(24);
output(0, 141) <= input(25);
output(0, 142) <= input(26);
output(0, 143) <= input(27);
output(0, 144) <= input(39);
output(0, 145) <= input(40);
output(0, 146) <= input(36);
output(0, 147) <= input(34);
output(0, 148) <= input(32);
output(0, 149) <= input(0);
output(0, 150) <= input(1);
output(0, 151) <= input(2);
output(0, 152) <= input(3);
output(0, 153) <= input(4);
output(0, 154) <= input(5);
output(0, 155) <= input(6);
output(0, 156) <= input(7);
output(0, 157) <= input(8);
output(0, 158) <= input(9);
output(0, 159) <= input(10);
output(0, 160) <= input(41);
output(0, 161) <= input(38);
output(0, 162) <= input(37);
output(0, 163) <= input(35);
output(0, 164) <= input(33);
output(0, 165) <= input(16);
output(0, 166) <= input(17);
output(0, 167) <= input(18);
output(0, 168) <= input(19);
output(0, 169) <= input(20);
output(0, 170) <= input(21);
output(0, 171) <= input(22);
output(0, 172) <= input(23);
output(0, 173) <= input(24);
output(0, 174) <= input(25);
output(0, 175) <= input(26);
output(0, 176) <= input(42);
output(0, 177) <= input(39);
output(0, 178) <= input(40);
output(0, 179) <= input(36);
output(0, 180) <= input(34);
output(0, 181) <= input(32);
output(0, 182) <= input(0);
output(0, 183) <= input(1);
output(0, 184) <= input(2);
output(0, 185) <= input(3);
output(0, 186) <= input(4);
output(0, 187) <= input(5);
output(0, 188) <= input(6);
output(0, 189) <= input(7);
output(0, 190) <= input(8);
output(0, 191) <= input(9);
output(0, 192) <= input(43);
output(0, 193) <= input(41);
output(0, 194) <= input(38);
output(0, 195) <= input(37);
output(0, 196) <= input(35);
output(0, 197) <= input(33);
output(0, 198) <= input(16);
output(0, 199) <= input(17);
output(0, 200) <= input(18);
output(0, 201) <= input(19);
output(0, 202) <= input(20);
output(0, 203) <= input(21);
output(0, 204) <= input(22);
output(0, 205) <= input(23);
output(0, 206) <= input(24);
output(0, 207) <= input(25);
output(0, 208) <= input(44);
output(0, 209) <= input(42);
output(0, 210) <= input(39);
output(0, 211) <= input(40);
output(0, 212) <= input(36);
output(0, 213) <= input(34);
output(0, 214) <= input(32);
output(0, 215) <= input(0);
output(0, 216) <= input(1);
output(0, 217) <= input(2);
output(0, 218) <= input(3);
output(0, 219) <= input(4);
output(0, 220) <= input(5);
output(0, 221) <= input(6);
output(0, 222) <= input(7);
output(0, 223) <= input(8);
output(0, 224) <= input(45);
output(0, 225) <= input(43);
output(0, 226) <= input(41);
output(0, 227) <= input(38);
output(0, 228) <= input(37);
output(0, 229) <= input(35);
output(0, 230) <= input(33);
output(0, 231) <= input(16);
output(0, 232) <= input(17);
output(0, 233) <= input(18);
output(0, 234) <= input(19);
output(0, 235) <= input(20);
output(0, 236) <= input(21);
output(0, 237) <= input(22);
output(0, 238) <= input(23);
output(0, 239) <= input(24);
output(0, 240) <= input(46);
output(0, 241) <= input(44);
output(0, 242) <= input(42);
output(0, 243) <= input(39);
output(0, 244) <= input(40);
output(0, 245) <= input(36);
output(0, 246) <= input(34);
output(0, 247) <= input(32);
output(0, 248) <= input(0);
output(0, 249) <= input(1);
output(0, 250) <= input(2);
output(0, 251) <= input(3);
output(0, 252) <= input(4);
output(0, 253) <= input(5);
output(0, 254) <= input(6);
output(0, 255) <= input(7);
output(1, 0) <= input(17);
output(1, 1) <= input(47);
output(1, 2) <= input(48);
output(1, 3) <= input(49);
output(1, 4) <= input(50);
output(1, 5) <= input(51);
output(1, 6) <= input(52);
output(1, 7) <= input(25);
output(1, 8) <= input(26);
output(1, 9) <= input(27);
output(1, 10) <= input(28);
output(1, 11) <= input(29);
output(1, 12) <= input(30);
output(1, 13) <= input(31);
output(1, 14) <= input(53);
output(1, 15) <= input(54);
output(1, 16) <= input(0);
output(1, 17) <= input(55);
output(1, 18) <= input(56);
output(1, 19) <= input(57);
output(1, 20) <= input(58);
output(1, 21) <= input(59);
output(1, 22) <= input(60);
output(1, 23) <= input(8);
output(1, 24) <= input(9);
output(1, 25) <= input(10);
output(1, 26) <= input(11);
output(1, 27) <= input(12);
output(1, 28) <= input(13);
output(1, 29) <= input(14);
output(1, 30) <= input(15);
output(1, 31) <= input(61);
output(1, 32) <= input(16);
output(1, 33) <= input(17);
output(1, 34) <= input(47);
output(1, 35) <= input(48);
output(1, 36) <= input(49);
output(1, 37) <= input(50);
output(1, 38) <= input(51);
output(1, 39) <= input(52);
output(1, 40) <= input(25);
output(1, 41) <= input(26);
output(1, 42) <= input(27);
output(1, 43) <= input(28);
output(1, 44) <= input(29);
output(1, 45) <= input(30);
output(1, 46) <= input(31);
output(1, 47) <= input(53);
output(1, 48) <= input(32);
output(1, 49) <= input(0);
output(1, 50) <= input(55);
output(1, 51) <= input(56);
output(1, 52) <= input(57);
output(1, 53) <= input(58);
output(1, 54) <= input(59);
output(1, 55) <= input(60);
output(1, 56) <= input(8);
output(1, 57) <= input(9);
output(1, 58) <= input(10);
output(1, 59) <= input(11);
output(1, 60) <= input(12);
output(1, 61) <= input(13);
output(1, 62) <= input(14);
output(1, 63) <= input(15);
output(1, 64) <= input(62);
output(1, 65) <= input(16);
output(1, 66) <= input(17);
output(1, 67) <= input(47);
output(1, 68) <= input(48);
output(1, 69) <= input(49);
output(1, 70) <= input(50);
output(1, 71) <= input(51);
output(1, 72) <= input(52);
output(1, 73) <= input(25);
output(1, 74) <= input(26);
output(1, 75) <= input(27);
output(1, 76) <= input(28);
output(1, 77) <= input(29);
output(1, 78) <= input(30);
output(1, 79) <= input(31);
output(1, 80) <= input(63);
output(1, 81) <= input(32);
output(1, 82) <= input(0);
output(1, 83) <= input(55);
output(1, 84) <= input(56);
output(1, 85) <= input(57);
output(1, 86) <= input(58);
output(1, 87) <= input(59);
output(1, 88) <= input(60);
output(1, 89) <= input(8);
output(1, 90) <= input(9);
output(1, 91) <= input(10);
output(1, 92) <= input(11);
output(1, 93) <= input(12);
output(1, 94) <= input(13);
output(1, 95) <= input(14);
output(1, 96) <= input(64);
output(1, 97) <= input(62);
output(1, 98) <= input(16);
output(1, 99) <= input(17);
output(1, 100) <= input(47);
output(1, 101) <= input(48);
output(1, 102) <= input(49);
output(1, 103) <= input(50);
output(1, 104) <= input(51);
output(1, 105) <= input(52);
output(1, 106) <= input(25);
output(1, 107) <= input(26);
output(1, 108) <= input(27);
output(1, 109) <= input(28);
output(1, 110) <= input(29);
output(1, 111) <= input(30);
output(1, 112) <= input(65);
output(1, 113) <= input(63);
output(1, 114) <= input(32);
output(1, 115) <= input(0);
output(1, 116) <= input(55);
output(1, 117) <= input(56);
output(1, 118) <= input(57);
output(1, 119) <= input(58);
output(1, 120) <= input(59);
output(1, 121) <= input(60);
output(1, 122) <= input(8);
output(1, 123) <= input(9);
output(1, 124) <= input(10);
output(1, 125) <= input(11);
output(1, 126) <= input(12);
output(1, 127) <= input(13);
output(1, 128) <= input(66);
output(1, 129) <= input(64);
output(1, 130) <= input(62);
output(1, 131) <= input(16);
output(1, 132) <= input(17);
output(1, 133) <= input(47);
output(1, 134) <= input(48);
output(1, 135) <= input(49);
output(1, 136) <= input(50);
output(1, 137) <= input(51);
output(1, 138) <= input(52);
output(1, 139) <= input(25);
output(1, 140) <= input(26);
output(1, 141) <= input(27);
output(1, 142) <= input(28);
output(1, 143) <= input(29);
output(1, 144) <= input(67);
output(1, 145) <= input(65);
output(1, 146) <= input(63);
output(1, 147) <= input(32);
output(1, 148) <= input(0);
output(1, 149) <= input(55);
output(1, 150) <= input(56);
output(1, 151) <= input(57);
output(1, 152) <= input(58);
output(1, 153) <= input(59);
output(1, 154) <= input(60);
output(1, 155) <= input(8);
output(1, 156) <= input(9);
output(1, 157) <= input(10);
output(1, 158) <= input(11);
output(1, 159) <= input(12);
output(1, 160) <= input(68);
output(1, 161) <= input(66);
output(1, 162) <= input(64);
output(1, 163) <= input(62);
output(1, 164) <= input(16);
output(1, 165) <= input(17);
output(1, 166) <= input(47);
output(1, 167) <= input(48);
output(1, 168) <= input(49);
output(1, 169) <= input(50);
output(1, 170) <= input(51);
output(1, 171) <= input(52);
output(1, 172) <= input(25);
output(1, 173) <= input(26);
output(1, 174) <= input(27);
output(1, 175) <= input(28);
output(1, 176) <= input(69);
output(1, 177) <= input(67);
output(1, 178) <= input(65);
output(1, 179) <= input(63);
output(1, 180) <= input(32);
output(1, 181) <= input(0);
output(1, 182) <= input(55);
output(1, 183) <= input(56);
output(1, 184) <= input(57);
output(1, 185) <= input(58);
output(1, 186) <= input(59);
output(1, 187) <= input(60);
output(1, 188) <= input(8);
output(1, 189) <= input(9);
output(1, 190) <= input(10);
output(1, 191) <= input(11);
output(1, 192) <= input(70);
output(1, 193) <= input(68);
output(1, 194) <= input(66);
output(1, 195) <= input(64);
output(1, 196) <= input(62);
output(1, 197) <= input(16);
output(1, 198) <= input(17);
output(1, 199) <= input(47);
output(1, 200) <= input(48);
output(1, 201) <= input(49);
output(1, 202) <= input(50);
output(1, 203) <= input(51);
output(1, 204) <= input(52);
output(1, 205) <= input(25);
output(1, 206) <= input(26);
output(1, 207) <= input(27);
output(1, 208) <= input(71);
output(1, 209) <= input(69);
output(1, 210) <= input(67);
output(1, 211) <= input(65);
output(1, 212) <= input(63);
output(1, 213) <= input(32);
output(1, 214) <= input(0);
output(1, 215) <= input(55);
output(1, 216) <= input(56);
output(1, 217) <= input(57);
output(1, 218) <= input(58);
output(1, 219) <= input(59);
output(1, 220) <= input(60);
output(1, 221) <= input(8);
output(1, 222) <= input(9);
output(1, 223) <= input(10);
output(1, 224) <= input(72);
output(1, 225) <= input(70);
output(1, 226) <= input(68);
output(1, 227) <= input(66);
output(1, 228) <= input(64);
output(1, 229) <= input(62);
output(1, 230) <= input(16);
output(1, 231) <= input(17);
output(1, 232) <= input(47);
output(1, 233) <= input(48);
output(1, 234) <= input(49);
output(1, 235) <= input(50);
output(1, 236) <= input(51);
output(1, 237) <= input(52);
output(1, 238) <= input(25);
output(1, 239) <= input(26);
output(1, 240) <= input(73);
output(1, 241) <= input(71);
output(1, 242) <= input(69);
output(1, 243) <= input(67);
output(1, 244) <= input(65);
output(1, 245) <= input(63);
output(1, 246) <= input(32);
output(1, 247) <= input(0);
output(1, 248) <= input(55);
output(1, 249) <= input(56);
output(1, 250) <= input(57);
output(1, 251) <= input(58);
output(1, 252) <= input(59);
output(1, 253) <= input(60);
output(1, 254) <= input(8);
output(1, 255) <= input(9);
when "1011" =>
output(0, 0) <= input(0);
output(0, 1) <= input(1);
output(0, 2) <= input(2);
output(0, 3) <= input(3);
output(0, 4) <= input(4);
output(0, 5) <= input(5);
output(0, 6) <= input(6);
output(0, 7) <= input(7);
output(0, 8) <= input(8);
output(0, 9) <= input(9);
output(0, 10) <= input(10);
output(0, 11) <= input(11);
output(0, 12) <= input(12);
output(0, 13) <= input(13);
output(0, 14) <= input(14);
output(0, 15) <= input(15);
output(0, 16) <= input(16);
output(0, 17) <= input(17);
output(0, 18) <= input(18);
output(0, 19) <= input(19);
output(0, 20) <= input(20);
output(0, 21) <= input(21);
output(0, 22) <= input(22);
output(0, 23) <= input(23);
output(0, 24) <= input(24);
output(0, 25) <= input(25);
output(0, 26) <= input(26);
output(0, 27) <= input(27);
output(0, 28) <= input(28);
output(0, 29) <= input(29);
output(0, 30) <= input(30);
output(0, 31) <= input(31);
output(0, 32) <= input(32);
output(0, 33) <= input(0);
output(0, 34) <= input(1);
output(0, 35) <= input(2);
output(0, 36) <= input(3);
output(0, 37) <= input(4);
output(0, 38) <= input(5);
output(0, 39) <= input(6);
output(0, 40) <= input(7);
output(0, 41) <= input(8);
output(0, 42) <= input(9);
output(0, 43) <= input(10);
output(0, 44) <= input(11);
output(0, 45) <= input(12);
output(0, 46) <= input(13);
output(0, 47) <= input(14);
output(0, 48) <= input(33);
output(0, 49) <= input(16);
output(0, 50) <= input(17);
output(0, 51) <= input(18);
output(0, 52) <= input(19);
output(0, 53) <= input(20);
output(0, 54) <= input(21);
output(0, 55) <= input(22);
output(0, 56) <= input(23);
output(0, 57) <= input(24);
output(0, 58) <= input(25);
output(0, 59) <= input(26);
output(0, 60) <= input(27);
output(0, 61) <= input(28);
output(0, 62) <= input(29);
output(0, 63) <= input(30);
output(0, 64) <= input(34);
output(0, 65) <= input(32);
output(0, 66) <= input(0);
output(0, 67) <= input(1);
output(0, 68) <= input(2);
output(0, 69) <= input(3);
output(0, 70) <= input(4);
output(0, 71) <= input(5);
output(0, 72) <= input(6);
output(0, 73) <= input(7);
output(0, 74) <= input(8);
output(0, 75) <= input(9);
output(0, 76) <= input(10);
output(0, 77) <= input(11);
output(0, 78) <= input(12);
output(0, 79) <= input(13);
output(0, 80) <= input(35);
output(0, 81) <= input(33);
output(0, 82) <= input(16);
output(0, 83) <= input(17);
output(0, 84) <= input(18);
output(0, 85) <= input(19);
output(0, 86) <= input(20);
output(0, 87) <= input(21);
output(0, 88) <= input(22);
output(0, 89) <= input(23);
output(0, 90) <= input(24);
output(0, 91) <= input(25);
output(0, 92) <= input(26);
output(0, 93) <= input(27);
output(0, 94) <= input(28);
output(0, 95) <= input(29);
output(0, 96) <= input(36);
output(0, 97) <= input(34);
output(0, 98) <= input(32);
output(0, 99) <= input(0);
output(0, 100) <= input(1);
output(0, 101) <= input(2);
output(0, 102) <= input(3);
output(0, 103) <= input(4);
output(0, 104) <= input(5);
output(0, 105) <= input(6);
output(0, 106) <= input(7);
output(0, 107) <= input(8);
output(0, 108) <= input(9);
output(0, 109) <= input(10);
output(0, 110) <= input(11);
output(0, 111) <= input(12);
output(0, 112) <= input(36);
output(0, 113) <= input(34);
output(0, 114) <= input(32);
output(0, 115) <= input(0);
output(0, 116) <= input(1);
output(0, 117) <= input(2);
output(0, 118) <= input(3);
output(0, 119) <= input(4);
output(0, 120) <= input(5);
output(0, 121) <= input(6);
output(0, 122) <= input(7);
output(0, 123) <= input(8);
output(0, 124) <= input(9);
output(0, 125) <= input(10);
output(0, 126) <= input(11);
output(0, 127) <= input(12);
output(0, 128) <= input(37);
output(0, 129) <= input(35);
output(0, 130) <= input(33);
output(0, 131) <= input(16);
output(0, 132) <= input(17);
output(0, 133) <= input(18);
output(0, 134) <= input(19);
output(0, 135) <= input(20);
output(0, 136) <= input(21);
output(0, 137) <= input(22);
output(0, 138) <= input(23);
output(0, 139) <= input(24);
output(0, 140) <= input(25);
output(0, 141) <= input(26);
output(0, 142) <= input(27);
output(0, 143) <= input(28);
output(0, 144) <= input(38);
output(0, 145) <= input(36);
output(0, 146) <= input(34);
output(0, 147) <= input(32);
output(0, 148) <= input(0);
output(0, 149) <= input(1);
output(0, 150) <= input(2);
output(0, 151) <= input(3);
output(0, 152) <= input(4);
output(0, 153) <= input(5);
output(0, 154) <= input(6);
output(0, 155) <= input(7);
output(0, 156) <= input(8);
output(0, 157) <= input(9);
output(0, 158) <= input(10);
output(0, 159) <= input(11);
output(0, 160) <= input(39);
output(0, 161) <= input(37);
output(0, 162) <= input(35);
output(0, 163) <= input(33);
output(0, 164) <= input(16);
output(0, 165) <= input(17);
output(0, 166) <= input(18);
output(0, 167) <= input(19);
output(0, 168) <= input(20);
output(0, 169) <= input(21);
output(0, 170) <= input(22);
output(0, 171) <= input(23);
output(0, 172) <= input(24);
output(0, 173) <= input(25);
output(0, 174) <= input(26);
output(0, 175) <= input(27);
output(0, 176) <= input(40);
output(0, 177) <= input(38);
output(0, 178) <= input(36);
output(0, 179) <= input(34);
output(0, 180) <= input(32);
output(0, 181) <= input(0);
output(0, 182) <= input(1);
output(0, 183) <= input(2);
output(0, 184) <= input(3);
output(0, 185) <= input(4);
output(0, 186) <= input(5);
output(0, 187) <= input(6);
output(0, 188) <= input(7);
output(0, 189) <= input(8);
output(0, 190) <= input(9);
output(0, 191) <= input(10);
output(0, 192) <= input(41);
output(0, 193) <= input(39);
output(0, 194) <= input(37);
output(0, 195) <= input(35);
output(0, 196) <= input(33);
output(0, 197) <= input(16);
output(0, 198) <= input(17);
output(0, 199) <= input(18);
output(0, 200) <= input(19);
output(0, 201) <= input(20);
output(0, 202) <= input(21);
output(0, 203) <= input(22);
output(0, 204) <= input(23);
output(0, 205) <= input(24);
output(0, 206) <= input(25);
output(0, 207) <= input(26);
output(0, 208) <= input(42);
output(0, 209) <= input(40);
output(0, 210) <= input(38);
output(0, 211) <= input(36);
output(0, 212) <= input(34);
output(0, 213) <= input(32);
output(0, 214) <= input(0);
output(0, 215) <= input(1);
output(0, 216) <= input(2);
output(0, 217) <= input(3);
output(0, 218) <= input(4);
output(0, 219) <= input(5);
output(0, 220) <= input(6);
output(0, 221) <= input(7);
output(0, 222) <= input(8);
output(0, 223) <= input(9);
output(0, 224) <= input(43);
output(0, 225) <= input(41);
output(0, 226) <= input(39);
output(0, 227) <= input(37);
output(0, 228) <= input(35);
output(0, 229) <= input(33);
output(0, 230) <= input(16);
output(0, 231) <= input(17);
output(0, 232) <= input(18);
output(0, 233) <= input(19);
output(0, 234) <= input(20);
output(0, 235) <= input(21);
output(0, 236) <= input(22);
output(0, 237) <= input(23);
output(0, 238) <= input(24);
output(0, 239) <= input(25);
output(0, 240) <= input(43);
output(0, 241) <= input(41);
output(0, 242) <= input(39);
output(0, 243) <= input(37);
output(0, 244) <= input(35);
output(0, 245) <= input(33);
output(0, 246) <= input(16);
output(0, 247) <= input(17);
output(0, 248) <= input(18);
output(0, 249) <= input(19);
output(0, 250) <= input(20);
output(0, 251) <= input(21);
output(0, 252) <= input(22);
output(0, 253) <= input(23);
output(0, 254) <= input(24);
output(0, 255) <= input(25);
output(1, 0) <= input(44);
output(1, 1) <= input(45);
output(1, 2) <= input(46);
output(1, 3) <= input(47);
output(1, 4) <= input(48);
output(1, 5) <= input(49);
output(1, 6) <= input(50);
output(1, 7) <= input(8);
output(1, 8) <= input(9);
output(1, 9) <= input(10);
output(1, 10) <= input(11);
output(1, 11) <= input(12);
output(1, 12) <= input(13);
output(1, 13) <= input(14);
output(1, 14) <= input(15);
output(1, 15) <= input(51);
output(1, 16) <= input(52);
output(1, 17) <= input(53);
output(1, 18) <= input(54);
output(1, 19) <= input(55);
output(1, 20) <= input(56);
output(1, 21) <= input(57);
output(1, 22) <= input(58);
output(1, 23) <= input(24);
output(1, 24) <= input(25);
output(1, 25) <= input(26);
output(1, 26) <= input(27);
output(1, 27) <= input(28);
output(1, 28) <= input(29);
output(1, 29) <= input(30);
output(1, 30) <= input(31);
output(1, 31) <= input(59);
output(1, 32) <= input(60);
output(1, 33) <= input(44);
output(1, 34) <= input(45);
output(1, 35) <= input(46);
output(1, 36) <= input(47);
output(1, 37) <= input(48);
output(1, 38) <= input(49);
output(1, 39) <= input(50);
output(1, 40) <= input(8);
output(1, 41) <= input(9);
output(1, 42) <= input(10);
output(1, 43) <= input(11);
output(1, 44) <= input(12);
output(1, 45) <= input(13);
output(1, 46) <= input(14);
output(1, 47) <= input(15);
output(1, 48) <= input(60);
output(1, 49) <= input(44);
output(1, 50) <= input(45);
output(1, 51) <= input(46);
output(1, 52) <= input(47);
output(1, 53) <= input(48);
output(1, 54) <= input(49);
output(1, 55) <= input(50);
output(1, 56) <= input(8);
output(1, 57) <= input(9);
output(1, 58) <= input(10);
output(1, 59) <= input(11);
output(1, 60) <= input(12);
output(1, 61) <= input(13);
output(1, 62) <= input(14);
output(1, 63) <= input(15);
output(1, 64) <= input(61);
output(1, 65) <= input(52);
output(1, 66) <= input(53);
output(1, 67) <= input(54);
output(1, 68) <= input(55);
output(1, 69) <= input(56);
output(1, 70) <= input(57);
output(1, 71) <= input(58);
output(1, 72) <= input(24);
output(1, 73) <= input(25);
output(1, 74) <= input(26);
output(1, 75) <= input(27);
output(1, 76) <= input(28);
output(1, 77) <= input(29);
output(1, 78) <= input(30);
output(1, 79) <= input(31);
output(1, 80) <= input(62);
output(1, 81) <= input(60);
output(1, 82) <= input(44);
output(1, 83) <= input(45);
output(1, 84) <= input(46);
output(1, 85) <= input(47);
output(1, 86) <= input(48);
output(1, 87) <= input(49);
output(1, 88) <= input(50);
output(1, 89) <= input(8);
output(1, 90) <= input(9);
output(1, 91) <= input(10);
output(1, 92) <= input(11);
output(1, 93) <= input(12);
output(1, 94) <= input(13);
output(1, 95) <= input(14);
output(1, 96) <= input(63);
output(1, 97) <= input(61);
output(1, 98) <= input(52);
output(1, 99) <= input(53);
output(1, 100) <= input(54);
output(1, 101) <= input(55);
output(1, 102) <= input(56);
output(1, 103) <= input(57);
output(1, 104) <= input(58);
output(1, 105) <= input(24);
output(1, 106) <= input(25);
output(1, 107) <= input(26);
output(1, 108) <= input(27);
output(1, 109) <= input(28);
output(1, 110) <= input(29);
output(1, 111) <= input(30);
output(1, 112) <= input(63);
output(1, 113) <= input(61);
output(1, 114) <= input(52);
output(1, 115) <= input(53);
output(1, 116) <= input(54);
output(1, 117) <= input(55);
output(1, 118) <= input(56);
output(1, 119) <= input(57);
output(1, 120) <= input(58);
output(1, 121) <= input(24);
output(1, 122) <= input(25);
output(1, 123) <= input(26);
output(1, 124) <= input(27);
output(1, 125) <= input(28);
output(1, 126) <= input(29);
output(1, 127) <= input(30);
output(1, 128) <= input(64);
output(1, 129) <= input(62);
output(1, 130) <= input(60);
output(1, 131) <= input(44);
output(1, 132) <= input(45);
output(1, 133) <= input(46);
output(1, 134) <= input(47);
output(1, 135) <= input(48);
output(1, 136) <= input(49);
output(1, 137) <= input(50);
output(1, 138) <= input(8);
output(1, 139) <= input(9);
output(1, 140) <= input(10);
output(1, 141) <= input(11);
output(1, 142) <= input(12);
output(1, 143) <= input(13);
output(1, 144) <= input(65);
output(1, 145) <= input(63);
output(1, 146) <= input(61);
output(1, 147) <= input(52);
output(1, 148) <= input(53);
output(1, 149) <= input(54);
output(1, 150) <= input(55);
output(1, 151) <= input(56);
output(1, 152) <= input(57);
output(1, 153) <= input(58);
output(1, 154) <= input(24);
output(1, 155) <= input(25);
output(1, 156) <= input(26);
output(1, 157) <= input(27);
output(1, 158) <= input(28);
output(1, 159) <= input(29);
output(1, 160) <= input(66);
output(1, 161) <= input(64);
output(1, 162) <= input(62);
output(1, 163) <= input(60);
output(1, 164) <= input(44);
output(1, 165) <= input(45);
output(1, 166) <= input(46);
output(1, 167) <= input(47);
output(1, 168) <= input(48);
output(1, 169) <= input(49);
output(1, 170) <= input(50);
output(1, 171) <= input(8);
output(1, 172) <= input(9);
output(1, 173) <= input(10);
output(1, 174) <= input(11);
output(1, 175) <= input(12);
output(1, 176) <= input(66);
output(1, 177) <= input(64);
output(1, 178) <= input(62);
output(1, 179) <= input(60);
output(1, 180) <= input(44);
output(1, 181) <= input(45);
output(1, 182) <= input(46);
output(1, 183) <= input(47);
output(1, 184) <= input(48);
output(1, 185) <= input(49);
output(1, 186) <= input(50);
output(1, 187) <= input(8);
output(1, 188) <= input(9);
output(1, 189) <= input(10);
output(1, 190) <= input(11);
output(1, 191) <= input(12);
output(1, 192) <= input(67);
output(1, 193) <= input(65);
output(1, 194) <= input(63);
output(1, 195) <= input(61);
output(1, 196) <= input(52);
output(1, 197) <= input(53);
output(1, 198) <= input(54);
output(1, 199) <= input(55);
output(1, 200) <= input(56);
output(1, 201) <= input(57);
output(1, 202) <= input(58);
output(1, 203) <= input(24);
output(1, 204) <= input(25);
output(1, 205) <= input(26);
output(1, 206) <= input(27);
output(1, 207) <= input(28);
output(1, 208) <= input(68);
output(1, 209) <= input(66);
output(1, 210) <= input(64);
output(1, 211) <= input(62);
output(1, 212) <= input(60);
output(1, 213) <= input(44);
output(1, 214) <= input(45);
output(1, 215) <= input(46);
output(1, 216) <= input(47);
output(1, 217) <= input(48);
output(1, 218) <= input(49);
output(1, 219) <= input(50);
output(1, 220) <= input(8);
output(1, 221) <= input(9);
output(1, 222) <= input(10);
output(1, 223) <= input(11);
output(1, 224) <= input(69);
output(1, 225) <= input(67);
output(1, 226) <= input(65);
output(1, 227) <= input(63);
output(1, 228) <= input(61);
output(1, 229) <= input(52);
output(1, 230) <= input(53);
output(1, 231) <= input(54);
output(1, 232) <= input(55);
output(1, 233) <= input(56);
output(1, 234) <= input(57);
output(1, 235) <= input(58);
output(1, 236) <= input(24);
output(1, 237) <= input(25);
output(1, 238) <= input(26);
output(1, 239) <= input(27);
output(1, 240) <= input(69);
output(1, 241) <= input(67);
output(1, 242) <= input(65);
output(1, 243) <= input(63);
output(1, 244) <= input(61);
output(1, 245) <= input(52);
output(1, 246) <= input(53);
output(1, 247) <= input(54);
output(1, 248) <= input(55);
output(1, 249) <= input(56);
output(1, 250) <= input(57);
output(1, 251) <= input(58);
output(1, 252) <= input(24);
output(1, 253) <= input(25);
output(1, 254) <= input(26);
output(1, 255) <= input(27);
output(2, 0) <= input(70);
output(2, 1) <= input(71);
output(2, 2) <= input(72);
output(2, 3) <= input(73);
output(2, 4) <= input(74);
output(2, 5) <= input(50);
output(2, 6) <= input(8);
output(2, 7) <= input(9);
output(2, 8) <= input(10);
output(2, 9) <= input(11);
output(2, 10) <= input(12);
output(2, 11) <= input(13);
output(2, 12) <= input(14);
output(2, 13) <= input(15);
output(2, 14) <= input(51);
output(2, 15) <= input(75);
output(2, 16) <= input(76);
output(2, 17) <= input(77);
output(2, 18) <= input(78);
output(2, 19) <= input(79);
output(2, 20) <= input(80);
output(2, 21) <= input(58);
output(2, 22) <= input(24);
output(2, 23) <= input(25);
output(2, 24) <= input(26);
output(2, 25) <= input(27);
output(2, 26) <= input(28);
output(2, 27) <= input(29);
output(2, 28) <= input(30);
output(2, 29) <= input(31);
output(2, 30) <= input(59);
output(2, 31) <= input(81);
output(2, 32) <= input(76);
output(2, 33) <= input(77);
output(2, 34) <= input(78);
output(2, 35) <= input(79);
output(2, 36) <= input(80);
output(2, 37) <= input(58);
output(2, 38) <= input(24);
output(2, 39) <= input(25);
output(2, 40) <= input(26);
output(2, 41) <= input(27);
output(2, 42) <= input(28);
output(2, 43) <= input(29);
output(2, 44) <= input(30);
output(2, 45) <= input(31);
output(2, 46) <= input(59);
output(2, 47) <= input(81);
output(2, 48) <= input(82);
output(2, 49) <= input(70);
output(2, 50) <= input(71);
output(2, 51) <= input(72);
output(2, 52) <= input(73);
output(2, 53) <= input(74);
output(2, 54) <= input(50);
output(2, 55) <= input(8);
output(2, 56) <= input(9);
output(2, 57) <= input(10);
output(2, 58) <= input(11);
output(2, 59) <= input(12);
output(2, 60) <= input(13);
output(2, 61) <= input(14);
output(2, 62) <= input(15);
output(2, 63) <= input(51);
output(2, 64) <= input(83);
output(2, 65) <= input(76);
output(2, 66) <= input(77);
output(2, 67) <= input(78);
output(2, 68) <= input(79);
output(2, 69) <= input(80);
output(2, 70) <= input(58);
output(2, 71) <= input(24);
output(2, 72) <= input(25);
output(2, 73) <= input(26);
output(2, 74) <= input(27);
output(2, 75) <= input(28);
output(2, 76) <= input(29);
output(2, 77) <= input(30);
output(2, 78) <= input(31);
output(2, 79) <= input(59);
output(2, 80) <= input(83);
output(2, 81) <= input(76);
output(2, 82) <= input(77);
output(2, 83) <= input(78);
output(2, 84) <= input(79);
output(2, 85) <= input(80);
output(2, 86) <= input(58);
output(2, 87) <= input(24);
output(2, 88) <= input(25);
output(2, 89) <= input(26);
output(2, 90) <= input(27);
output(2, 91) <= input(28);
output(2, 92) <= input(29);
output(2, 93) <= input(30);
output(2, 94) <= input(31);
output(2, 95) <= input(59);
output(2, 96) <= input(84);
output(2, 97) <= input(82);
output(2, 98) <= input(70);
output(2, 99) <= input(71);
output(2, 100) <= input(72);
output(2, 101) <= input(73);
output(2, 102) <= input(74);
output(2, 103) <= input(50);
output(2, 104) <= input(8);
output(2, 105) <= input(9);
output(2, 106) <= input(10);
output(2, 107) <= input(11);
output(2, 108) <= input(12);
output(2, 109) <= input(13);
output(2, 110) <= input(14);
output(2, 111) <= input(15);
output(2, 112) <= input(84);
output(2, 113) <= input(82);
output(2, 114) <= input(70);
output(2, 115) <= input(71);
output(2, 116) <= input(72);
output(2, 117) <= input(73);
output(2, 118) <= input(74);
output(2, 119) <= input(50);
output(2, 120) <= input(8);
output(2, 121) <= input(9);
output(2, 122) <= input(10);
output(2, 123) <= input(11);
output(2, 124) <= input(12);
output(2, 125) <= input(13);
output(2, 126) <= input(14);
output(2, 127) <= input(15);
output(2, 128) <= input(85);
output(2, 129) <= input(83);
output(2, 130) <= input(76);
output(2, 131) <= input(77);
output(2, 132) <= input(78);
output(2, 133) <= input(79);
output(2, 134) <= input(80);
output(2, 135) <= input(58);
output(2, 136) <= input(24);
output(2, 137) <= input(25);
output(2, 138) <= input(26);
output(2, 139) <= input(27);
output(2, 140) <= input(28);
output(2, 141) <= input(29);
output(2, 142) <= input(30);
output(2, 143) <= input(31);
output(2, 144) <= input(86);
output(2, 145) <= input(84);
output(2, 146) <= input(82);
output(2, 147) <= input(70);
output(2, 148) <= input(71);
output(2, 149) <= input(72);
output(2, 150) <= input(73);
output(2, 151) <= input(74);
output(2, 152) <= input(50);
output(2, 153) <= input(8);
output(2, 154) <= input(9);
output(2, 155) <= input(10);
output(2, 156) <= input(11);
output(2, 157) <= input(12);
output(2, 158) <= input(13);
output(2, 159) <= input(14);
output(2, 160) <= input(86);
output(2, 161) <= input(84);
output(2, 162) <= input(82);
output(2, 163) <= input(70);
output(2, 164) <= input(71);
output(2, 165) <= input(72);
output(2, 166) <= input(73);
output(2, 167) <= input(74);
output(2, 168) <= input(50);
output(2, 169) <= input(8);
output(2, 170) <= input(9);
output(2, 171) <= input(10);
output(2, 172) <= input(11);
output(2, 173) <= input(12);
output(2, 174) <= input(13);
output(2, 175) <= input(14);
output(2, 176) <= input(87);
output(2, 177) <= input(85);
output(2, 178) <= input(83);
output(2, 179) <= input(76);
output(2, 180) <= input(77);
output(2, 181) <= input(78);
output(2, 182) <= input(79);
output(2, 183) <= input(80);
output(2, 184) <= input(58);
output(2, 185) <= input(24);
output(2, 186) <= input(25);
output(2, 187) <= input(26);
output(2, 188) <= input(27);
output(2, 189) <= input(28);
output(2, 190) <= input(29);
output(2, 191) <= input(30);
output(2, 192) <= input(88);
output(2, 193) <= input(86);
output(2, 194) <= input(84);
output(2, 195) <= input(82);
output(2, 196) <= input(70);
output(2, 197) <= input(71);
output(2, 198) <= input(72);
output(2, 199) <= input(73);
output(2, 200) <= input(74);
output(2, 201) <= input(50);
output(2, 202) <= input(8);
output(2, 203) <= input(9);
output(2, 204) <= input(10);
output(2, 205) <= input(11);
output(2, 206) <= input(12);
output(2, 207) <= input(13);
output(2, 208) <= input(88);
output(2, 209) <= input(86);
output(2, 210) <= input(84);
output(2, 211) <= input(82);
output(2, 212) <= input(70);
output(2, 213) <= input(71);
output(2, 214) <= input(72);
output(2, 215) <= input(73);
output(2, 216) <= input(74);
output(2, 217) <= input(50);
output(2, 218) <= input(8);
output(2, 219) <= input(9);
output(2, 220) <= input(10);
output(2, 221) <= input(11);
output(2, 222) <= input(12);
output(2, 223) <= input(13);
output(2, 224) <= input(89);
output(2, 225) <= input(87);
output(2, 226) <= input(85);
output(2, 227) <= input(83);
output(2, 228) <= input(76);
output(2, 229) <= input(77);
output(2, 230) <= input(78);
output(2, 231) <= input(79);
output(2, 232) <= input(80);
output(2, 233) <= input(58);
output(2, 234) <= input(24);
output(2, 235) <= input(25);
output(2, 236) <= input(26);
output(2, 237) <= input(27);
output(2, 238) <= input(28);
output(2, 239) <= input(29);
output(2, 240) <= input(89);
output(2, 241) <= input(87);
output(2, 242) <= input(85);
output(2, 243) <= input(83);
output(2, 244) <= input(76);
output(2, 245) <= input(77);
output(2, 246) <= input(78);
output(2, 247) <= input(79);
output(2, 248) <= input(80);
output(2, 249) <= input(58);
output(2, 250) <= input(24);
output(2, 251) <= input(25);
output(2, 252) <= input(26);
output(2, 253) <= input(27);
output(2, 254) <= input(28);
output(2, 255) <= input(29);
when "1100" =>
output(0, 0) <= input(0);
output(0, 1) <= input(1);
output(0, 2) <= input(2);
output(0, 3) <= input(3);
output(0, 4) <= input(4);
output(0, 5) <= input(5);
output(0, 6) <= input(6);
output(0, 7) <= input(7);
output(0, 8) <= input(8);
output(0, 9) <= input(9);
output(0, 10) <= input(10);
output(0, 11) <= input(11);
output(0, 12) <= input(12);
output(0, 13) <= input(13);
output(0, 14) <= input(14);
output(0, 15) <= input(15);
output(0, 16) <= input(0);
output(0, 17) <= input(1);
output(0, 18) <= input(2);
output(0, 19) <= input(3);
output(0, 20) <= input(4);
output(0, 21) <= input(5);
output(0, 22) <= input(6);
output(0, 23) <= input(7);
output(0, 24) <= input(8);
output(0, 25) <= input(9);
output(0, 26) <= input(10);
output(0, 27) <= input(11);
output(0, 28) <= input(12);
output(0, 29) <= input(13);
output(0, 30) <= input(14);
output(0, 31) <= input(15);
output(0, 32) <= input(16);
output(0, 33) <= input(17);
output(0, 34) <= input(18);
output(0, 35) <= input(19);
output(0, 36) <= input(20);
output(0, 37) <= input(21);
output(0, 38) <= input(22);
output(0, 39) <= input(23);
output(0, 40) <= input(24);
output(0, 41) <= input(25);
output(0, 42) <= input(26);
output(0, 43) <= input(27);
output(0, 44) <= input(28);
output(0, 45) <= input(29);
output(0, 46) <= input(30);
output(0, 47) <= input(31);
output(0, 48) <= input(16);
output(0, 49) <= input(17);
output(0, 50) <= input(18);
output(0, 51) <= input(19);
output(0, 52) <= input(20);
output(0, 53) <= input(21);
output(0, 54) <= input(22);
output(0, 55) <= input(23);
output(0, 56) <= input(24);
output(0, 57) <= input(25);
output(0, 58) <= input(26);
output(0, 59) <= input(27);
output(0, 60) <= input(28);
output(0, 61) <= input(29);
output(0, 62) <= input(30);
output(0, 63) <= input(31);
output(0, 64) <= input(32);
output(0, 65) <= input(0);
output(0, 66) <= input(1);
output(0, 67) <= input(2);
output(0, 68) <= input(3);
output(0, 69) <= input(4);
output(0, 70) <= input(5);
output(0, 71) <= input(6);
output(0, 72) <= input(7);
output(0, 73) <= input(8);
output(0, 74) <= input(9);
output(0, 75) <= input(10);
output(0, 76) <= input(11);
output(0, 77) <= input(12);
output(0, 78) <= input(13);
output(0, 79) <= input(14);
output(0, 80) <= input(32);
output(0, 81) <= input(0);
output(0, 82) <= input(1);
output(0, 83) <= input(2);
output(0, 84) <= input(3);
output(0, 85) <= input(4);
output(0, 86) <= input(5);
output(0, 87) <= input(6);
output(0, 88) <= input(7);
output(0, 89) <= input(8);
output(0, 90) <= input(9);
output(0, 91) <= input(10);
output(0, 92) <= input(11);
output(0, 93) <= input(12);
output(0, 94) <= input(13);
output(0, 95) <= input(14);
output(0, 96) <= input(33);
output(0, 97) <= input(16);
output(0, 98) <= input(17);
output(0, 99) <= input(18);
output(0, 100) <= input(19);
output(0, 101) <= input(20);
output(0, 102) <= input(21);
output(0, 103) <= input(22);
output(0, 104) <= input(23);
output(0, 105) <= input(24);
output(0, 106) <= input(25);
output(0, 107) <= input(26);
output(0, 108) <= input(27);
output(0, 109) <= input(28);
output(0, 110) <= input(29);
output(0, 111) <= input(30);
output(0, 112) <= input(33);
output(0, 113) <= input(16);
output(0, 114) <= input(17);
output(0, 115) <= input(18);
output(0, 116) <= input(19);
output(0, 117) <= input(20);
output(0, 118) <= input(21);
output(0, 119) <= input(22);
output(0, 120) <= input(23);
output(0, 121) <= input(24);
output(0, 122) <= input(25);
output(0, 123) <= input(26);
output(0, 124) <= input(27);
output(0, 125) <= input(28);
output(0, 126) <= input(29);
output(0, 127) <= input(30);
output(0, 128) <= input(34);
output(0, 129) <= input(32);
output(0, 130) <= input(0);
output(0, 131) <= input(1);
output(0, 132) <= input(2);
output(0, 133) <= input(3);
output(0, 134) <= input(4);
output(0, 135) <= input(5);
output(0, 136) <= input(6);
output(0, 137) <= input(7);
output(0, 138) <= input(8);
output(0, 139) <= input(9);
output(0, 140) <= input(10);
output(0, 141) <= input(11);
output(0, 142) <= input(12);
output(0, 143) <= input(13);
output(0, 144) <= input(34);
output(0, 145) <= input(32);
output(0, 146) <= input(0);
output(0, 147) <= input(1);
output(0, 148) <= input(2);
output(0, 149) <= input(3);
output(0, 150) <= input(4);
output(0, 151) <= input(5);
output(0, 152) <= input(6);
output(0, 153) <= input(7);
output(0, 154) <= input(8);
output(0, 155) <= input(9);
output(0, 156) <= input(10);
output(0, 157) <= input(11);
output(0, 158) <= input(12);
output(0, 159) <= input(13);
output(0, 160) <= input(35);
output(0, 161) <= input(33);
output(0, 162) <= input(16);
output(0, 163) <= input(17);
output(0, 164) <= input(18);
output(0, 165) <= input(19);
output(0, 166) <= input(20);
output(0, 167) <= input(21);
output(0, 168) <= input(22);
output(0, 169) <= input(23);
output(0, 170) <= input(24);
output(0, 171) <= input(25);
output(0, 172) <= input(26);
output(0, 173) <= input(27);
output(0, 174) <= input(28);
output(0, 175) <= input(29);
output(0, 176) <= input(35);
output(0, 177) <= input(33);
output(0, 178) <= input(16);
output(0, 179) <= input(17);
output(0, 180) <= input(18);
output(0, 181) <= input(19);
output(0, 182) <= input(20);
output(0, 183) <= input(21);
output(0, 184) <= input(22);
output(0, 185) <= input(23);
output(0, 186) <= input(24);
output(0, 187) <= input(25);
output(0, 188) <= input(26);
output(0, 189) <= input(27);
output(0, 190) <= input(28);
output(0, 191) <= input(29);
output(0, 192) <= input(36);
output(0, 193) <= input(34);
output(0, 194) <= input(32);
output(0, 195) <= input(0);
output(0, 196) <= input(1);
output(0, 197) <= input(2);
output(0, 198) <= input(3);
output(0, 199) <= input(4);
output(0, 200) <= input(5);
output(0, 201) <= input(6);
output(0, 202) <= input(7);
output(0, 203) <= input(8);
output(0, 204) <= input(9);
output(0, 205) <= input(10);
output(0, 206) <= input(11);
output(0, 207) <= input(12);
output(0, 208) <= input(36);
output(0, 209) <= input(34);
output(0, 210) <= input(32);
output(0, 211) <= input(0);
output(0, 212) <= input(1);
output(0, 213) <= input(2);
output(0, 214) <= input(3);
output(0, 215) <= input(4);
output(0, 216) <= input(5);
output(0, 217) <= input(6);
output(0, 218) <= input(7);
output(0, 219) <= input(8);
output(0, 220) <= input(9);
output(0, 221) <= input(10);
output(0, 222) <= input(11);
output(0, 223) <= input(12);
output(0, 224) <= input(37);
output(0, 225) <= input(35);
output(0, 226) <= input(33);
output(0, 227) <= input(16);
output(0, 228) <= input(17);
output(0, 229) <= input(18);
output(0, 230) <= input(19);
output(0, 231) <= input(20);
output(0, 232) <= input(21);
output(0, 233) <= input(22);
output(0, 234) <= input(23);
output(0, 235) <= input(24);
output(0, 236) <= input(25);
output(0, 237) <= input(26);
output(0, 238) <= input(27);
output(0, 239) <= input(28);
output(0, 240) <= input(37);
output(0, 241) <= input(35);
output(0, 242) <= input(33);
output(0, 243) <= input(16);
output(0, 244) <= input(17);
output(0, 245) <= input(18);
output(0, 246) <= input(19);
output(0, 247) <= input(20);
output(0, 248) <= input(21);
output(0, 249) <= input(22);
output(0, 250) <= input(23);
output(0, 251) <= input(24);
output(0, 252) <= input(25);
output(0, 253) <= input(26);
output(0, 254) <= input(27);
output(0, 255) <= input(28);
output(1, 0) <= input(38);
output(1, 1) <= input(39);
output(1, 2) <= input(40);
output(1, 3) <= input(41);
output(1, 4) <= input(5);
output(1, 5) <= input(6);
output(1, 6) <= input(7);
output(1, 7) <= input(8);
output(1, 8) <= input(9);
output(1, 9) <= input(10);
output(1, 10) <= input(11);
output(1, 11) <= input(12);
output(1, 12) <= input(13);
output(1, 13) <= input(14);
output(1, 14) <= input(15);
output(1, 15) <= input(42);
output(1, 16) <= input(38);
output(1, 17) <= input(39);
output(1, 18) <= input(40);
output(1, 19) <= input(41);
output(1, 20) <= input(5);
output(1, 21) <= input(6);
output(1, 22) <= input(7);
output(1, 23) <= input(8);
output(1, 24) <= input(9);
output(1, 25) <= input(10);
output(1, 26) <= input(11);
output(1, 27) <= input(12);
output(1, 28) <= input(13);
output(1, 29) <= input(14);
output(1, 30) <= input(15);
output(1, 31) <= input(42);
output(1, 32) <= input(43);
output(1, 33) <= input(44);
output(1, 34) <= input(45);
output(1, 35) <= input(46);
output(1, 36) <= input(21);
output(1, 37) <= input(22);
output(1, 38) <= input(23);
output(1, 39) <= input(24);
output(1, 40) <= input(25);
output(1, 41) <= input(26);
output(1, 42) <= input(27);
output(1, 43) <= input(28);
output(1, 44) <= input(29);
output(1, 45) <= input(30);
output(1, 46) <= input(31);
output(1, 47) <= input(47);
output(1, 48) <= input(43);
output(1, 49) <= input(44);
output(1, 50) <= input(45);
output(1, 51) <= input(46);
output(1, 52) <= input(21);
output(1, 53) <= input(22);
output(1, 54) <= input(23);
output(1, 55) <= input(24);
output(1, 56) <= input(25);
output(1, 57) <= input(26);
output(1, 58) <= input(27);
output(1, 59) <= input(28);
output(1, 60) <= input(29);
output(1, 61) <= input(30);
output(1, 62) <= input(31);
output(1, 63) <= input(47);
output(1, 64) <= input(43);
output(1, 65) <= input(44);
output(1, 66) <= input(45);
output(1, 67) <= input(46);
output(1, 68) <= input(21);
output(1, 69) <= input(22);
output(1, 70) <= input(23);
output(1, 71) <= input(24);
output(1, 72) <= input(25);
output(1, 73) <= input(26);
output(1, 74) <= input(27);
output(1, 75) <= input(28);
output(1, 76) <= input(29);
output(1, 77) <= input(30);
output(1, 78) <= input(31);
output(1, 79) <= input(47);
output(1, 80) <= input(48);
output(1, 81) <= input(38);
output(1, 82) <= input(39);
output(1, 83) <= input(40);
output(1, 84) <= input(41);
output(1, 85) <= input(5);
output(1, 86) <= input(6);
output(1, 87) <= input(7);
output(1, 88) <= input(8);
output(1, 89) <= input(9);
output(1, 90) <= input(10);
output(1, 91) <= input(11);
output(1, 92) <= input(12);
output(1, 93) <= input(13);
output(1, 94) <= input(14);
output(1, 95) <= input(15);
output(1, 96) <= input(48);
output(1, 97) <= input(38);
output(1, 98) <= input(39);
output(1, 99) <= input(40);
output(1, 100) <= input(41);
output(1, 101) <= input(5);
output(1, 102) <= input(6);
output(1, 103) <= input(7);
output(1, 104) <= input(8);
output(1, 105) <= input(9);
output(1, 106) <= input(10);
output(1, 107) <= input(11);
output(1, 108) <= input(12);
output(1, 109) <= input(13);
output(1, 110) <= input(14);
output(1, 111) <= input(15);
output(1, 112) <= input(48);
output(1, 113) <= input(38);
output(1, 114) <= input(39);
output(1, 115) <= input(40);
output(1, 116) <= input(41);
output(1, 117) <= input(5);
output(1, 118) <= input(6);
output(1, 119) <= input(7);
output(1, 120) <= input(8);
output(1, 121) <= input(9);
output(1, 122) <= input(10);
output(1, 123) <= input(11);
output(1, 124) <= input(12);
output(1, 125) <= input(13);
output(1, 126) <= input(14);
output(1, 127) <= input(15);
output(1, 128) <= input(49);
output(1, 129) <= input(43);
output(1, 130) <= input(44);
output(1, 131) <= input(45);
output(1, 132) <= input(46);
output(1, 133) <= input(21);
output(1, 134) <= input(22);
output(1, 135) <= input(23);
output(1, 136) <= input(24);
output(1, 137) <= input(25);
output(1, 138) <= input(26);
output(1, 139) <= input(27);
output(1, 140) <= input(28);
output(1, 141) <= input(29);
output(1, 142) <= input(30);
output(1, 143) <= input(31);
output(1, 144) <= input(49);
output(1, 145) <= input(43);
output(1, 146) <= input(44);
output(1, 147) <= input(45);
output(1, 148) <= input(46);
output(1, 149) <= input(21);
output(1, 150) <= input(22);
output(1, 151) <= input(23);
output(1, 152) <= input(24);
output(1, 153) <= input(25);
output(1, 154) <= input(26);
output(1, 155) <= input(27);
output(1, 156) <= input(28);
output(1, 157) <= input(29);
output(1, 158) <= input(30);
output(1, 159) <= input(31);
output(1, 160) <= input(50);
output(1, 161) <= input(48);
output(1, 162) <= input(38);
output(1, 163) <= input(39);
output(1, 164) <= input(40);
output(1, 165) <= input(41);
output(1, 166) <= input(5);
output(1, 167) <= input(6);
output(1, 168) <= input(7);
output(1, 169) <= input(8);
output(1, 170) <= input(9);
output(1, 171) <= input(10);
output(1, 172) <= input(11);
output(1, 173) <= input(12);
output(1, 174) <= input(13);
output(1, 175) <= input(14);
output(1, 176) <= input(50);
output(1, 177) <= input(48);
output(1, 178) <= input(38);
output(1, 179) <= input(39);
output(1, 180) <= input(40);
output(1, 181) <= input(41);
output(1, 182) <= input(5);
output(1, 183) <= input(6);
output(1, 184) <= input(7);
output(1, 185) <= input(8);
output(1, 186) <= input(9);
output(1, 187) <= input(10);
output(1, 188) <= input(11);
output(1, 189) <= input(12);
output(1, 190) <= input(13);
output(1, 191) <= input(14);
output(1, 192) <= input(50);
output(1, 193) <= input(48);
output(1, 194) <= input(38);
output(1, 195) <= input(39);
output(1, 196) <= input(40);
output(1, 197) <= input(41);
output(1, 198) <= input(5);
output(1, 199) <= input(6);
output(1, 200) <= input(7);
output(1, 201) <= input(8);
output(1, 202) <= input(9);
output(1, 203) <= input(10);
output(1, 204) <= input(11);
output(1, 205) <= input(12);
output(1, 206) <= input(13);
output(1, 207) <= input(14);
output(1, 208) <= input(51);
output(1, 209) <= input(49);
output(1, 210) <= input(43);
output(1, 211) <= input(44);
output(1, 212) <= input(45);
output(1, 213) <= input(46);
output(1, 214) <= input(21);
output(1, 215) <= input(22);
output(1, 216) <= input(23);
output(1, 217) <= input(24);
output(1, 218) <= input(25);
output(1, 219) <= input(26);
output(1, 220) <= input(27);
output(1, 221) <= input(28);
output(1, 222) <= input(29);
output(1, 223) <= input(30);
output(1, 224) <= input(51);
output(1, 225) <= input(49);
output(1, 226) <= input(43);
output(1, 227) <= input(44);
output(1, 228) <= input(45);
output(1, 229) <= input(46);
output(1, 230) <= input(21);
output(1, 231) <= input(22);
output(1, 232) <= input(23);
output(1, 233) <= input(24);
output(1, 234) <= input(25);
output(1, 235) <= input(26);
output(1, 236) <= input(27);
output(1, 237) <= input(28);
output(1, 238) <= input(29);
output(1, 239) <= input(30);
output(1, 240) <= input(51);
output(1, 241) <= input(49);
output(1, 242) <= input(43);
output(1, 243) <= input(44);
output(1, 244) <= input(45);
output(1, 245) <= input(46);
output(1, 246) <= input(21);
output(1, 247) <= input(22);
output(1, 248) <= input(23);
output(1, 249) <= input(24);
output(1, 250) <= input(25);
output(1, 251) <= input(26);
output(1, 252) <= input(27);
output(1, 253) <= input(28);
output(1, 254) <= input(29);
output(1, 255) <= input(30);
output(2, 0) <= input(52);
output(2, 1) <= input(53);
output(2, 2) <= input(54);
output(2, 3) <= input(5);
output(2, 4) <= input(6);
output(2, 5) <= input(7);
output(2, 6) <= input(8);
output(2, 7) <= input(9);
output(2, 8) <= input(10);
output(2, 9) <= input(11);
output(2, 10) <= input(12);
output(2, 11) <= input(13);
output(2, 12) <= input(14);
output(2, 13) <= input(15);
output(2, 14) <= input(42);
output(2, 15) <= input(55);
output(2, 16) <= input(52);
output(2, 17) <= input(53);
output(2, 18) <= input(54);
output(2, 19) <= input(5);
output(2, 20) <= input(6);
output(2, 21) <= input(7);
output(2, 22) <= input(8);
output(2, 23) <= input(9);
output(2, 24) <= input(10);
output(2, 25) <= input(11);
output(2, 26) <= input(12);
output(2, 27) <= input(13);
output(2, 28) <= input(14);
output(2, 29) <= input(15);
output(2, 30) <= input(42);
output(2, 31) <= input(55);
output(2, 32) <= input(52);
output(2, 33) <= input(53);
output(2, 34) <= input(54);
output(2, 35) <= input(5);
output(2, 36) <= input(6);
output(2, 37) <= input(7);
output(2, 38) <= input(8);
output(2, 39) <= input(9);
output(2, 40) <= input(10);
output(2, 41) <= input(11);
output(2, 42) <= input(12);
output(2, 43) <= input(13);
output(2, 44) <= input(14);
output(2, 45) <= input(15);
output(2, 46) <= input(42);
output(2, 47) <= input(55);
output(2, 48) <= input(52);
output(2, 49) <= input(53);
output(2, 50) <= input(54);
output(2, 51) <= input(5);
output(2, 52) <= input(6);
output(2, 53) <= input(7);
output(2, 54) <= input(8);
output(2, 55) <= input(9);
output(2, 56) <= input(10);
output(2, 57) <= input(11);
output(2, 58) <= input(12);
output(2, 59) <= input(13);
output(2, 60) <= input(14);
output(2, 61) <= input(15);
output(2, 62) <= input(42);
output(2, 63) <= input(55);
output(2, 64) <= input(56);
output(2, 65) <= input(57);
output(2, 66) <= input(58);
output(2, 67) <= input(21);
output(2, 68) <= input(22);
output(2, 69) <= input(23);
output(2, 70) <= input(24);
output(2, 71) <= input(25);
output(2, 72) <= input(26);
output(2, 73) <= input(27);
output(2, 74) <= input(28);
output(2, 75) <= input(29);
output(2, 76) <= input(30);
output(2, 77) <= input(31);
output(2, 78) <= input(47);
output(2, 79) <= input(59);
output(2, 80) <= input(56);
output(2, 81) <= input(57);
output(2, 82) <= input(58);
output(2, 83) <= input(21);
output(2, 84) <= input(22);
output(2, 85) <= input(23);
output(2, 86) <= input(24);
output(2, 87) <= input(25);
output(2, 88) <= input(26);
output(2, 89) <= input(27);
output(2, 90) <= input(28);
output(2, 91) <= input(29);
output(2, 92) <= input(30);
output(2, 93) <= input(31);
output(2, 94) <= input(47);
output(2, 95) <= input(59);
output(2, 96) <= input(56);
output(2, 97) <= input(57);
output(2, 98) <= input(58);
output(2, 99) <= input(21);
output(2, 100) <= input(22);
output(2, 101) <= input(23);
output(2, 102) <= input(24);
output(2, 103) <= input(25);
output(2, 104) <= input(26);
output(2, 105) <= input(27);
output(2, 106) <= input(28);
output(2, 107) <= input(29);
output(2, 108) <= input(30);
output(2, 109) <= input(31);
output(2, 110) <= input(47);
output(2, 111) <= input(59);
output(2, 112) <= input(56);
output(2, 113) <= input(57);
output(2, 114) <= input(58);
output(2, 115) <= input(21);
output(2, 116) <= input(22);
output(2, 117) <= input(23);
output(2, 118) <= input(24);
output(2, 119) <= input(25);
output(2, 120) <= input(26);
output(2, 121) <= input(27);
output(2, 122) <= input(28);
output(2, 123) <= input(29);
output(2, 124) <= input(30);
output(2, 125) <= input(31);
output(2, 126) <= input(47);
output(2, 127) <= input(59);
output(2, 128) <= input(60);
output(2, 129) <= input(52);
output(2, 130) <= input(53);
output(2, 131) <= input(54);
output(2, 132) <= input(5);
output(2, 133) <= input(6);
output(2, 134) <= input(7);
output(2, 135) <= input(8);
output(2, 136) <= input(9);
output(2, 137) <= input(10);
output(2, 138) <= input(11);
output(2, 139) <= input(12);
output(2, 140) <= input(13);
output(2, 141) <= input(14);
output(2, 142) <= input(15);
output(2, 143) <= input(42);
output(2, 144) <= input(60);
output(2, 145) <= input(52);
output(2, 146) <= input(53);
output(2, 147) <= input(54);
output(2, 148) <= input(5);
output(2, 149) <= input(6);
output(2, 150) <= input(7);
output(2, 151) <= input(8);
output(2, 152) <= input(9);
output(2, 153) <= input(10);
output(2, 154) <= input(11);
output(2, 155) <= input(12);
output(2, 156) <= input(13);
output(2, 157) <= input(14);
output(2, 158) <= input(15);
output(2, 159) <= input(42);
output(2, 160) <= input(60);
output(2, 161) <= input(52);
output(2, 162) <= input(53);
output(2, 163) <= input(54);
output(2, 164) <= input(5);
output(2, 165) <= input(6);
output(2, 166) <= input(7);
output(2, 167) <= input(8);
output(2, 168) <= input(9);
output(2, 169) <= input(10);
output(2, 170) <= input(11);
output(2, 171) <= input(12);
output(2, 172) <= input(13);
output(2, 173) <= input(14);
output(2, 174) <= input(15);
output(2, 175) <= input(42);
output(2, 176) <= input(60);
output(2, 177) <= input(52);
output(2, 178) <= input(53);
output(2, 179) <= input(54);
output(2, 180) <= input(5);
output(2, 181) <= input(6);
output(2, 182) <= input(7);
output(2, 183) <= input(8);
output(2, 184) <= input(9);
output(2, 185) <= input(10);
output(2, 186) <= input(11);
output(2, 187) <= input(12);
output(2, 188) <= input(13);
output(2, 189) <= input(14);
output(2, 190) <= input(15);
output(2, 191) <= input(42);
output(2, 192) <= input(61);
output(2, 193) <= input(56);
output(2, 194) <= input(57);
output(2, 195) <= input(58);
output(2, 196) <= input(21);
output(2, 197) <= input(22);
output(2, 198) <= input(23);
output(2, 199) <= input(24);
output(2, 200) <= input(25);
output(2, 201) <= input(26);
output(2, 202) <= input(27);
output(2, 203) <= input(28);
output(2, 204) <= input(29);
output(2, 205) <= input(30);
output(2, 206) <= input(31);
output(2, 207) <= input(47);
output(2, 208) <= input(61);
output(2, 209) <= input(56);
output(2, 210) <= input(57);
output(2, 211) <= input(58);
output(2, 212) <= input(21);
output(2, 213) <= input(22);
output(2, 214) <= input(23);
output(2, 215) <= input(24);
output(2, 216) <= input(25);
output(2, 217) <= input(26);
output(2, 218) <= input(27);
output(2, 219) <= input(28);
output(2, 220) <= input(29);
output(2, 221) <= input(30);
output(2, 222) <= input(31);
output(2, 223) <= input(47);
output(2, 224) <= input(61);
output(2, 225) <= input(56);
output(2, 226) <= input(57);
output(2, 227) <= input(58);
output(2, 228) <= input(21);
output(2, 229) <= input(22);
output(2, 230) <= input(23);
output(2, 231) <= input(24);
output(2, 232) <= input(25);
output(2, 233) <= input(26);
output(2, 234) <= input(27);
output(2, 235) <= input(28);
output(2, 236) <= input(29);
output(2, 237) <= input(30);
output(2, 238) <= input(31);
output(2, 239) <= input(47);
output(2, 240) <= input(61);
output(2, 241) <= input(56);
output(2, 242) <= input(57);
output(2, 243) <= input(58);
output(2, 244) <= input(21);
output(2, 245) <= input(22);
output(2, 246) <= input(23);
output(2, 247) <= input(24);
output(2, 248) <= input(25);
output(2, 249) <= input(26);
output(2, 250) <= input(27);
output(2, 251) <= input(28);
output(2, 252) <= input(29);
output(2, 253) <= input(30);
output(2, 254) <= input(31);
output(2, 255) <= input(47);
when "1101" =>
output(0, 0) <= input(0);
output(0, 1) <= input(1);
output(0, 2) <= input(2);
output(0, 3) <= input(3);
output(0, 4) <= input(4);
output(0, 5) <= input(5);
output(0, 6) <= input(6);
output(0, 7) <= input(7);
output(0, 8) <= input(8);
output(0, 9) <= input(9);
output(0, 10) <= input(10);
output(0, 11) <= input(11);
output(0, 12) <= input(12);
output(0, 13) <= input(13);
output(0, 14) <= input(14);
output(0, 15) <= input(15);
output(0, 16) <= input(0);
output(0, 17) <= input(1);
output(0, 18) <= input(2);
output(0, 19) <= input(3);
output(0, 20) <= input(4);
output(0, 21) <= input(5);
output(0, 22) <= input(6);
output(0, 23) <= input(7);
output(0, 24) <= input(8);
output(0, 25) <= input(9);
output(0, 26) <= input(10);
output(0, 27) <= input(11);
output(0, 28) <= input(12);
output(0, 29) <= input(13);
output(0, 30) <= input(14);
output(0, 31) <= input(15);
output(0, 32) <= input(0);
output(0, 33) <= input(1);
output(0, 34) <= input(2);
output(0, 35) <= input(3);
output(0, 36) <= input(4);
output(0, 37) <= input(5);
output(0, 38) <= input(6);
output(0, 39) <= input(7);
output(0, 40) <= input(8);
output(0, 41) <= input(9);
output(0, 42) <= input(10);
output(0, 43) <= input(11);
output(0, 44) <= input(12);
output(0, 45) <= input(13);
output(0, 46) <= input(14);
output(0, 47) <= input(15);
output(0, 48) <= input(0);
output(0, 49) <= input(1);
output(0, 50) <= input(2);
output(0, 51) <= input(3);
output(0, 52) <= input(4);
output(0, 53) <= input(5);
output(0, 54) <= input(6);
output(0, 55) <= input(7);
output(0, 56) <= input(8);
output(0, 57) <= input(9);
output(0, 58) <= input(10);
output(0, 59) <= input(11);
output(0, 60) <= input(12);
output(0, 61) <= input(13);
output(0, 62) <= input(14);
output(0, 63) <= input(15);
output(0, 64) <= input(0);
output(0, 65) <= input(1);
output(0, 66) <= input(2);
output(0, 67) <= input(3);
output(0, 68) <= input(4);
output(0, 69) <= input(5);
output(0, 70) <= input(6);
output(0, 71) <= input(7);
output(0, 72) <= input(8);
output(0, 73) <= input(9);
output(0, 74) <= input(10);
output(0, 75) <= input(11);
output(0, 76) <= input(12);
output(0, 77) <= input(13);
output(0, 78) <= input(14);
output(0, 79) <= input(15);
output(0, 80) <= input(16);
output(0, 81) <= input(17);
output(0, 82) <= input(18);
output(0, 83) <= input(19);
output(0, 84) <= input(20);
output(0, 85) <= input(21);
output(0, 86) <= input(22);
output(0, 87) <= input(23);
output(0, 88) <= input(24);
output(0, 89) <= input(25);
output(0, 90) <= input(26);
output(0, 91) <= input(27);
output(0, 92) <= input(28);
output(0, 93) <= input(29);
output(0, 94) <= input(30);
output(0, 95) <= input(31);
output(0, 96) <= input(16);
output(0, 97) <= input(17);
output(0, 98) <= input(18);
output(0, 99) <= input(19);
output(0, 100) <= input(20);
output(0, 101) <= input(21);
output(0, 102) <= input(22);
output(0, 103) <= input(23);
output(0, 104) <= input(24);
output(0, 105) <= input(25);
output(0, 106) <= input(26);
output(0, 107) <= input(27);
output(0, 108) <= input(28);
output(0, 109) <= input(29);
output(0, 110) <= input(30);
output(0, 111) <= input(31);
output(0, 112) <= input(16);
output(0, 113) <= input(17);
output(0, 114) <= input(18);
output(0, 115) <= input(19);
output(0, 116) <= input(20);
output(0, 117) <= input(21);
output(0, 118) <= input(22);
output(0, 119) <= input(23);
output(0, 120) <= input(24);
output(0, 121) <= input(25);
output(0, 122) <= input(26);
output(0, 123) <= input(27);
output(0, 124) <= input(28);
output(0, 125) <= input(29);
output(0, 126) <= input(30);
output(0, 127) <= input(31);
output(0, 128) <= input(16);
output(0, 129) <= input(17);
output(0, 130) <= input(18);
output(0, 131) <= input(19);
output(0, 132) <= input(20);
output(0, 133) <= input(21);
output(0, 134) <= input(22);
output(0, 135) <= input(23);
output(0, 136) <= input(24);
output(0, 137) <= input(25);
output(0, 138) <= input(26);
output(0, 139) <= input(27);
output(0, 140) <= input(28);
output(0, 141) <= input(29);
output(0, 142) <= input(30);
output(0, 143) <= input(31);
output(0, 144) <= input(16);
output(0, 145) <= input(17);
output(0, 146) <= input(18);
output(0, 147) <= input(19);
output(0, 148) <= input(20);
output(0, 149) <= input(21);
output(0, 150) <= input(22);
output(0, 151) <= input(23);
output(0, 152) <= input(24);
output(0, 153) <= input(25);
output(0, 154) <= input(26);
output(0, 155) <= input(27);
output(0, 156) <= input(28);
output(0, 157) <= input(29);
output(0, 158) <= input(30);
output(0, 159) <= input(31);
output(0, 160) <= input(32);
output(0, 161) <= input(0);
output(0, 162) <= input(1);
output(0, 163) <= input(2);
output(0, 164) <= input(3);
output(0, 165) <= input(4);
output(0, 166) <= input(5);
output(0, 167) <= input(6);
output(0, 168) <= input(7);
output(0, 169) <= input(8);
output(0, 170) <= input(9);
output(0, 171) <= input(10);
output(0, 172) <= input(11);
output(0, 173) <= input(12);
output(0, 174) <= input(13);
output(0, 175) <= input(14);
output(0, 176) <= input(32);
output(0, 177) <= input(0);
output(0, 178) <= input(1);
output(0, 179) <= input(2);
output(0, 180) <= input(3);
output(0, 181) <= input(4);
output(0, 182) <= input(5);
output(0, 183) <= input(6);
output(0, 184) <= input(7);
output(0, 185) <= input(8);
output(0, 186) <= input(9);
output(0, 187) <= input(10);
output(0, 188) <= input(11);
output(0, 189) <= input(12);
output(0, 190) <= input(13);
output(0, 191) <= input(14);
output(0, 192) <= input(32);
output(0, 193) <= input(0);
output(0, 194) <= input(1);
output(0, 195) <= input(2);
output(0, 196) <= input(3);
output(0, 197) <= input(4);
output(0, 198) <= input(5);
output(0, 199) <= input(6);
output(0, 200) <= input(7);
output(0, 201) <= input(8);
output(0, 202) <= input(9);
output(0, 203) <= input(10);
output(0, 204) <= input(11);
output(0, 205) <= input(12);
output(0, 206) <= input(13);
output(0, 207) <= input(14);
output(0, 208) <= input(32);
output(0, 209) <= input(0);
output(0, 210) <= input(1);
output(0, 211) <= input(2);
output(0, 212) <= input(3);
output(0, 213) <= input(4);
output(0, 214) <= input(5);
output(0, 215) <= input(6);
output(0, 216) <= input(7);
output(0, 217) <= input(8);
output(0, 218) <= input(9);
output(0, 219) <= input(10);
output(0, 220) <= input(11);
output(0, 221) <= input(12);
output(0, 222) <= input(13);
output(0, 223) <= input(14);
output(0, 224) <= input(32);
output(0, 225) <= input(0);
output(0, 226) <= input(1);
output(0, 227) <= input(2);
output(0, 228) <= input(3);
output(0, 229) <= input(4);
output(0, 230) <= input(5);
output(0, 231) <= input(6);
output(0, 232) <= input(7);
output(0, 233) <= input(8);
output(0, 234) <= input(9);
output(0, 235) <= input(10);
output(0, 236) <= input(11);
output(0, 237) <= input(12);
output(0, 238) <= input(13);
output(0, 239) <= input(14);
output(0, 240) <= input(32);
output(0, 241) <= input(0);
output(0, 242) <= input(1);
output(0, 243) <= input(2);
output(0, 244) <= input(3);
output(0, 245) <= input(4);
output(0, 246) <= input(5);
output(0, 247) <= input(6);
output(0, 248) <= input(7);
output(0, 249) <= input(8);
output(0, 250) <= input(9);
output(0, 251) <= input(10);
output(0, 252) <= input(11);
output(0, 253) <= input(12);
output(0, 254) <= input(13);
output(0, 255) <= input(14);
output(1, 0) <= input(33);
output(1, 1) <= input(34);
output(1, 2) <= input(19);
output(1, 3) <= input(20);
output(1, 4) <= input(21);
output(1, 5) <= input(22);
output(1, 6) <= input(23);
output(1, 7) <= input(24);
output(1, 8) <= input(25);
output(1, 9) <= input(26);
output(1, 10) <= input(27);
output(1, 11) <= input(28);
output(1, 12) <= input(29);
output(1, 13) <= input(30);
output(1, 14) <= input(31);
output(1, 15) <= input(35);
output(1, 16) <= input(33);
output(1, 17) <= input(34);
output(1, 18) <= input(19);
output(1, 19) <= input(20);
output(1, 20) <= input(21);
output(1, 21) <= input(22);
output(1, 22) <= input(23);
output(1, 23) <= input(24);
output(1, 24) <= input(25);
output(1, 25) <= input(26);
output(1, 26) <= input(27);
output(1, 27) <= input(28);
output(1, 28) <= input(29);
output(1, 29) <= input(30);
output(1, 30) <= input(31);
output(1, 31) <= input(35);
output(1, 32) <= input(33);
output(1, 33) <= input(34);
output(1, 34) <= input(19);
output(1, 35) <= input(20);
output(1, 36) <= input(21);
output(1, 37) <= input(22);
output(1, 38) <= input(23);
output(1, 39) <= input(24);
output(1, 40) <= input(25);
output(1, 41) <= input(26);
output(1, 42) <= input(27);
output(1, 43) <= input(28);
output(1, 44) <= input(29);
output(1, 45) <= input(30);
output(1, 46) <= input(31);
output(1, 47) <= input(35);
output(1, 48) <= input(33);
output(1, 49) <= input(34);
output(1, 50) <= input(19);
output(1, 51) <= input(20);
output(1, 52) <= input(21);
output(1, 53) <= input(22);
output(1, 54) <= input(23);
output(1, 55) <= input(24);
output(1, 56) <= input(25);
output(1, 57) <= input(26);
output(1, 58) <= input(27);
output(1, 59) <= input(28);
output(1, 60) <= input(29);
output(1, 61) <= input(30);
output(1, 62) <= input(31);
output(1, 63) <= input(35);
output(1, 64) <= input(33);
output(1, 65) <= input(34);
output(1, 66) <= input(19);
output(1, 67) <= input(20);
output(1, 68) <= input(21);
output(1, 69) <= input(22);
output(1, 70) <= input(23);
output(1, 71) <= input(24);
output(1, 72) <= input(25);
output(1, 73) <= input(26);
output(1, 74) <= input(27);
output(1, 75) <= input(28);
output(1, 76) <= input(29);
output(1, 77) <= input(30);
output(1, 78) <= input(31);
output(1, 79) <= input(35);
output(1, 80) <= input(33);
output(1, 81) <= input(34);
output(1, 82) <= input(19);
output(1, 83) <= input(20);
output(1, 84) <= input(21);
output(1, 85) <= input(22);
output(1, 86) <= input(23);
output(1, 87) <= input(24);
output(1, 88) <= input(25);
output(1, 89) <= input(26);
output(1, 90) <= input(27);
output(1, 91) <= input(28);
output(1, 92) <= input(29);
output(1, 93) <= input(30);
output(1, 94) <= input(31);
output(1, 95) <= input(35);
output(1, 96) <= input(33);
output(1, 97) <= input(34);
output(1, 98) <= input(19);
output(1, 99) <= input(20);
output(1, 100) <= input(21);
output(1, 101) <= input(22);
output(1, 102) <= input(23);
output(1, 103) <= input(24);
output(1, 104) <= input(25);
output(1, 105) <= input(26);
output(1, 106) <= input(27);
output(1, 107) <= input(28);
output(1, 108) <= input(29);
output(1, 109) <= input(30);
output(1, 110) <= input(31);
output(1, 111) <= input(35);
output(1, 112) <= input(33);
output(1, 113) <= input(34);
output(1, 114) <= input(19);
output(1, 115) <= input(20);
output(1, 116) <= input(21);
output(1, 117) <= input(22);
output(1, 118) <= input(23);
output(1, 119) <= input(24);
output(1, 120) <= input(25);
output(1, 121) <= input(26);
output(1, 122) <= input(27);
output(1, 123) <= input(28);
output(1, 124) <= input(29);
output(1, 125) <= input(30);
output(1, 126) <= input(31);
output(1, 127) <= input(35);
output(1, 128) <= input(36);
output(1, 129) <= input(37);
output(1, 130) <= input(2);
output(1, 131) <= input(3);
output(1, 132) <= input(4);
output(1, 133) <= input(5);
output(1, 134) <= input(6);
output(1, 135) <= input(7);
output(1, 136) <= input(8);
output(1, 137) <= input(9);
output(1, 138) <= input(10);
output(1, 139) <= input(11);
output(1, 140) <= input(12);
output(1, 141) <= input(13);
output(1, 142) <= input(14);
output(1, 143) <= input(15);
output(1, 144) <= input(36);
output(1, 145) <= input(37);
output(1, 146) <= input(2);
output(1, 147) <= input(3);
output(1, 148) <= input(4);
output(1, 149) <= input(5);
output(1, 150) <= input(6);
output(1, 151) <= input(7);
output(1, 152) <= input(8);
output(1, 153) <= input(9);
output(1, 154) <= input(10);
output(1, 155) <= input(11);
output(1, 156) <= input(12);
output(1, 157) <= input(13);
output(1, 158) <= input(14);
output(1, 159) <= input(15);
output(1, 160) <= input(36);
output(1, 161) <= input(37);
output(1, 162) <= input(2);
output(1, 163) <= input(3);
output(1, 164) <= input(4);
output(1, 165) <= input(5);
output(1, 166) <= input(6);
output(1, 167) <= input(7);
output(1, 168) <= input(8);
output(1, 169) <= input(9);
output(1, 170) <= input(10);
output(1, 171) <= input(11);
output(1, 172) <= input(12);
output(1, 173) <= input(13);
output(1, 174) <= input(14);
output(1, 175) <= input(15);
output(1, 176) <= input(36);
output(1, 177) <= input(37);
output(1, 178) <= input(2);
output(1, 179) <= input(3);
output(1, 180) <= input(4);
output(1, 181) <= input(5);
output(1, 182) <= input(6);
output(1, 183) <= input(7);
output(1, 184) <= input(8);
output(1, 185) <= input(9);
output(1, 186) <= input(10);
output(1, 187) <= input(11);
output(1, 188) <= input(12);
output(1, 189) <= input(13);
output(1, 190) <= input(14);
output(1, 191) <= input(15);
output(1, 192) <= input(36);
output(1, 193) <= input(37);
output(1, 194) <= input(2);
output(1, 195) <= input(3);
output(1, 196) <= input(4);
output(1, 197) <= input(5);
output(1, 198) <= input(6);
output(1, 199) <= input(7);
output(1, 200) <= input(8);
output(1, 201) <= input(9);
output(1, 202) <= input(10);
output(1, 203) <= input(11);
output(1, 204) <= input(12);
output(1, 205) <= input(13);
output(1, 206) <= input(14);
output(1, 207) <= input(15);
output(1, 208) <= input(36);
output(1, 209) <= input(37);
output(1, 210) <= input(2);
output(1, 211) <= input(3);
output(1, 212) <= input(4);
output(1, 213) <= input(5);
output(1, 214) <= input(6);
output(1, 215) <= input(7);
output(1, 216) <= input(8);
output(1, 217) <= input(9);
output(1, 218) <= input(10);
output(1, 219) <= input(11);
output(1, 220) <= input(12);
output(1, 221) <= input(13);
output(1, 222) <= input(14);
output(1, 223) <= input(15);
output(1, 224) <= input(36);
output(1, 225) <= input(37);
output(1, 226) <= input(2);
output(1, 227) <= input(3);
output(1, 228) <= input(4);
output(1, 229) <= input(5);
output(1, 230) <= input(6);
output(1, 231) <= input(7);
output(1, 232) <= input(8);
output(1, 233) <= input(9);
output(1, 234) <= input(10);
output(1, 235) <= input(11);
output(1, 236) <= input(12);
output(1, 237) <= input(13);
output(1, 238) <= input(14);
output(1, 239) <= input(15);
output(1, 240) <= input(36);
output(1, 241) <= input(37);
output(1, 242) <= input(2);
output(1, 243) <= input(3);
output(1, 244) <= input(4);
output(1, 245) <= input(5);
output(1, 246) <= input(6);
output(1, 247) <= input(7);
output(1, 248) <= input(8);
output(1, 249) <= input(9);
output(1, 250) <= input(10);
output(1, 251) <= input(11);
output(1, 252) <= input(12);
output(1, 253) <= input(13);
output(1, 254) <= input(14);
output(1, 255) <= input(15);
output(2, 0) <= input(38);
output(2, 1) <= input(2);
output(2, 2) <= input(3);
output(2, 3) <= input(4);
output(2, 4) <= input(5);
output(2, 5) <= input(6);
output(2, 6) <= input(7);
output(2, 7) <= input(8);
output(2, 8) <= input(9);
output(2, 9) <= input(10);
output(2, 10) <= input(11);
output(2, 11) <= input(12);
output(2, 12) <= input(13);
output(2, 13) <= input(14);
output(2, 14) <= input(15);
output(2, 15) <= input(39);
output(2, 16) <= input(38);
output(2, 17) <= input(2);
output(2, 18) <= input(3);
output(2, 19) <= input(4);
output(2, 20) <= input(5);
output(2, 21) <= input(6);
output(2, 22) <= input(7);
output(2, 23) <= input(8);
output(2, 24) <= input(9);
output(2, 25) <= input(10);
output(2, 26) <= input(11);
output(2, 27) <= input(12);
output(2, 28) <= input(13);
output(2, 29) <= input(14);
output(2, 30) <= input(15);
output(2, 31) <= input(39);
output(2, 32) <= input(38);
output(2, 33) <= input(2);
output(2, 34) <= input(3);
output(2, 35) <= input(4);
output(2, 36) <= input(5);
output(2, 37) <= input(6);
output(2, 38) <= input(7);
output(2, 39) <= input(8);
output(2, 40) <= input(9);
output(2, 41) <= input(10);
output(2, 42) <= input(11);
output(2, 43) <= input(12);
output(2, 44) <= input(13);
output(2, 45) <= input(14);
output(2, 46) <= input(15);
output(2, 47) <= input(39);
output(2, 48) <= input(38);
output(2, 49) <= input(2);
output(2, 50) <= input(3);
output(2, 51) <= input(4);
output(2, 52) <= input(5);
output(2, 53) <= input(6);
output(2, 54) <= input(7);
output(2, 55) <= input(8);
output(2, 56) <= input(9);
output(2, 57) <= input(10);
output(2, 58) <= input(11);
output(2, 59) <= input(12);
output(2, 60) <= input(13);
output(2, 61) <= input(14);
output(2, 62) <= input(15);
output(2, 63) <= input(39);
output(2, 64) <= input(38);
output(2, 65) <= input(2);
output(2, 66) <= input(3);
output(2, 67) <= input(4);
output(2, 68) <= input(5);
output(2, 69) <= input(6);
output(2, 70) <= input(7);
output(2, 71) <= input(8);
output(2, 72) <= input(9);
output(2, 73) <= input(10);
output(2, 74) <= input(11);
output(2, 75) <= input(12);
output(2, 76) <= input(13);
output(2, 77) <= input(14);
output(2, 78) <= input(15);
output(2, 79) <= input(39);
output(2, 80) <= input(38);
output(2, 81) <= input(2);
output(2, 82) <= input(3);
output(2, 83) <= input(4);
output(2, 84) <= input(5);
output(2, 85) <= input(6);
output(2, 86) <= input(7);
output(2, 87) <= input(8);
output(2, 88) <= input(9);
output(2, 89) <= input(10);
output(2, 90) <= input(11);
output(2, 91) <= input(12);
output(2, 92) <= input(13);
output(2, 93) <= input(14);
output(2, 94) <= input(15);
output(2, 95) <= input(39);
output(2, 96) <= input(38);
output(2, 97) <= input(2);
output(2, 98) <= input(3);
output(2, 99) <= input(4);
output(2, 100) <= input(5);
output(2, 101) <= input(6);
output(2, 102) <= input(7);
output(2, 103) <= input(8);
output(2, 104) <= input(9);
output(2, 105) <= input(10);
output(2, 106) <= input(11);
output(2, 107) <= input(12);
output(2, 108) <= input(13);
output(2, 109) <= input(14);
output(2, 110) <= input(15);
output(2, 111) <= input(39);
output(2, 112) <= input(38);
output(2, 113) <= input(2);
output(2, 114) <= input(3);
output(2, 115) <= input(4);
output(2, 116) <= input(5);
output(2, 117) <= input(6);
output(2, 118) <= input(7);
output(2, 119) <= input(8);
output(2, 120) <= input(9);
output(2, 121) <= input(10);
output(2, 122) <= input(11);
output(2, 123) <= input(12);
output(2, 124) <= input(13);
output(2, 125) <= input(14);
output(2, 126) <= input(15);
output(2, 127) <= input(39);
output(2, 128) <= input(38);
output(2, 129) <= input(2);
output(2, 130) <= input(3);
output(2, 131) <= input(4);
output(2, 132) <= input(5);
output(2, 133) <= input(6);
output(2, 134) <= input(7);
output(2, 135) <= input(8);
output(2, 136) <= input(9);
output(2, 137) <= input(10);
output(2, 138) <= input(11);
output(2, 139) <= input(12);
output(2, 140) <= input(13);
output(2, 141) <= input(14);
output(2, 142) <= input(15);
output(2, 143) <= input(39);
output(2, 144) <= input(38);
output(2, 145) <= input(2);
output(2, 146) <= input(3);
output(2, 147) <= input(4);
output(2, 148) <= input(5);
output(2, 149) <= input(6);
output(2, 150) <= input(7);
output(2, 151) <= input(8);
output(2, 152) <= input(9);
output(2, 153) <= input(10);
output(2, 154) <= input(11);
output(2, 155) <= input(12);
output(2, 156) <= input(13);
output(2, 157) <= input(14);
output(2, 158) <= input(15);
output(2, 159) <= input(39);
output(2, 160) <= input(38);
output(2, 161) <= input(2);
output(2, 162) <= input(3);
output(2, 163) <= input(4);
output(2, 164) <= input(5);
output(2, 165) <= input(6);
output(2, 166) <= input(7);
output(2, 167) <= input(8);
output(2, 168) <= input(9);
output(2, 169) <= input(10);
output(2, 170) <= input(11);
output(2, 171) <= input(12);
output(2, 172) <= input(13);
output(2, 173) <= input(14);
output(2, 174) <= input(15);
output(2, 175) <= input(39);
output(2, 176) <= input(38);
output(2, 177) <= input(2);
output(2, 178) <= input(3);
output(2, 179) <= input(4);
output(2, 180) <= input(5);
output(2, 181) <= input(6);
output(2, 182) <= input(7);
output(2, 183) <= input(8);
output(2, 184) <= input(9);
output(2, 185) <= input(10);
output(2, 186) <= input(11);
output(2, 187) <= input(12);
output(2, 188) <= input(13);
output(2, 189) <= input(14);
output(2, 190) <= input(15);
output(2, 191) <= input(39);
output(2, 192) <= input(38);
output(2, 193) <= input(2);
output(2, 194) <= input(3);
output(2, 195) <= input(4);
output(2, 196) <= input(5);
output(2, 197) <= input(6);
output(2, 198) <= input(7);
output(2, 199) <= input(8);
output(2, 200) <= input(9);
output(2, 201) <= input(10);
output(2, 202) <= input(11);
output(2, 203) <= input(12);
output(2, 204) <= input(13);
output(2, 205) <= input(14);
output(2, 206) <= input(15);
output(2, 207) <= input(39);
output(2, 208) <= input(38);
output(2, 209) <= input(2);
output(2, 210) <= input(3);
output(2, 211) <= input(4);
output(2, 212) <= input(5);
output(2, 213) <= input(6);
output(2, 214) <= input(7);
output(2, 215) <= input(8);
output(2, 216) <= input(9);
output(2, 217) <= input(10);
output(2, 218) <= input(11);
output(2, 219) <= input(12);
output(2, 220) <= input(13);
output(2, 221) <= input(14);
output(2, 222) <= input(15);
output(2, 223) <= input(39);
output(2, 224) <= input(38);
output(2, 225) <= input(2);
output(2, 226) <= input(3);
output(2, 227) <= input(4);
output(2, 228) <= input(5);
output(2, 229) <= input(6);
output(2, 230) <= input(7);
output(2, 231) <= input(8);
output(2, 232) <= input(9);
output(2, 233) <= input(10);
output(2, 234) <= input(11);
output(2, 235) <= input(12);
output(2, 236) <= input(13);
output(2, 237) <= input(14);
output(2, 238) <= input(15);
output(2, 239) <= input(39);
output(2, 240) <= input(38);
output(2, 241) <= input(2);
output(2, 242) <= input(3);
output(2, 243) <= input(4);
output(2, 244) <= input(5);
output(2, 245) <= input(6);
output(2, 246) <= input(7);
output(2, 247) <= input(8);
output(2, 248) <= input(9);
output(2, 249) <= input(10);
output(2, 250) <= input(11);
output(2, 251) <= input(12);
output(2, 252) <= input(13);
output(2, 253) <= input(14);
output(2, 254) <= input(15);
output(2, 255) <= input(39);
output(3, 0) <= input(2);
output(3, 1) <= input(3);
output(3, 2) <= input(4);
output(3, 3) <= input(5);
output(3, 4) <= input(6);
output(3, 5) <= input(7);
output(3, 6) <= input(8);
output(3, 7) <= input(9);
output(3, 8) <= input(10);
output(3, 9) <= input(11);
output(3, 10) <= input(12);
output(3, 11) <= input(13);
output(3, 12) <= input(14);
output(3, 13) <= input(15);
output(3, 14) <= input(39);
output(3, 15) <= input(40);
output(3, 16) <= input(2);
output(3, 17) <= input(3);
output(3, 18) <= input(4);
output(3, 19) <= input(5);
output(3, 20) <= input(6);
output(3, 21) <= input(7);
output(3, 22) <= input(8);
output(3, 23) <= input(9);
output(3, 24) <= input(10);
output(3, 25) <= input(11);
output(3, 26) <= input(12);
output(3, 27) <= input(13);
output(3, 28) <= input(14);
output(3, 29) <= input(15);
output(3, 30) <= input(39);
output(3, 31) <= input(40);
output(3, 32) <= input(2);
output(3, 33) <= input(3);
output(3, 34) <= input(4);
output(3, 35) <= input(5);
output(3, 36) <= input(6);
output(3, 37) <= input(7);
output(3, 38) <= input(8);
output(3, 39) <= input(9);
output(3, 40) <= input(10);
output(3, 41) <= input(11);
output(3, 42) <= input(12);
output(3, 43) <= input(13);
output(3, 44) <= input(14);
output(3, 45) <= input(15);
output(3, 46) <= input(39);
output(3, 47) <= input(40);
output(3, 48) <= input(2);
output(3, 49) <= input(3);
output(3, 50) <= input(4);
output(3, 51) <= input(5);
output(3, 52) <= input(6);
output(3, 53) <= input(7);
output(3, 54) <= input(8);
output(3, 55) <= input(9);
output(3, 56) <= input(10);
output(3, 57) <= input(11);
output(3, 58) <= input(12);
output(3, 59) <= input(13);
output(3, 60) <= input(14);
output(3, 61) <= input(15);
output(3, 62) <= input(39);
output(3, 63) <= input(40);
output(3, 64) <= input(2);
output(3, 65) <= input(3);
output(3, 66) <= input(4);
output(3, 67) <= input(5);
output(3, 68) <= input(6);
output(3, 69) <= input(7);
output(3, 70) <= input(8);
output(3, 71) <= input(9);
output(3, 72) <= input(10);
output(3, 73) <= input(11);
output(3, 74) <= input(12);
output(3, 75) <= input(13);
output(3, 76) <= input(14);
output(3, 77) <= input(15);
output(3, 78) <= input(39);
output(3, 79) <= input(40);
output(3, 80) <= input(2);
output(3, 81) <= input(3);
output(3, 82) <= input(4);
output(3, 83) <= input(5);
output(3, 84) <= input(6);
output(3, 85) <= input(7);
output(3, 86) <= input(8);
output(3, 87) <= input(9);
output(3, 88) <= input(10);
output(3, 89) <= input(11);
output(3, 90) <= input(12);
output(3, 91) <= input(13);
output(3, 92) <= input(14);
output(3, 93) <= input(15);
output(3, 94) <= input(39);
output(3, 95) <= input(40);
output(3, 96) <= input(2);
output(3, 97) <= input(3);
output(3, 98) <= input(4);
output(3, 99) <= input(5);
output(3, 100) <= input(6);
output(3, 101) <= input(7);
output(3, 102) <= input(8);
output(3, 103) <= input(9);
output(3, 104) <= input(10);
output(3, 105) <= input(11);
output(3, 106) <= input(12);
output(3, 107) <= input(13);
output(3, 108) <= input(14);
output(3, 109) <= input(15);
output(3, 110) <= input(39);
output(3, 111) <= input(40);
output(3, 112) <= input(2);
output(3, 113) <= input(3);
output(3, 114) <= input(4);
output(3, 115) <= input(5);
output(3, 116) <= input(6);
output(3, 117) <= input(7);
output(3, 118) <= input(8);
output(3, 119) <= input(9);
output(3, 120) <= input(10);
output(3, 121) <= input(11);
output(3, 122) <= input(12);
output(3, 123) <= input(13);
output(3, 124) <= input(14);
output(3, 125) <= input(15);
output(3, 126) <= input(39);
output(3, 127) <= input(40);
output(3, 128) <= input(2);
output(3, 129) <= input(3);
output(3, 130) <= input(4);
output(3, 131) <= input(5);
output(3, 132) <= input(6);
output(3, 133) <= input(7);
output(3, 134) <= input(8);
output(3, 135) <= input(9);
output(3, 136) <= input(10);
output(3, 137) <= input(11);
output(3, 138) <= input(12);
output(3, 139) <= input(13);
output(3, 140) <= input(14);
output(3, 141) <= input(15);
output(3, 142) <= input(39);
output(3, 143) <= input(40);
output(3, 144) <= input(2);
output(3, 145) <= input(3);
output(3, 146) <= input(4);
output(3, 147) <= input(5);
output(3, 148) <= input(6);
output(3, 149) <= input(7);
output(3, 150) <= input(8);
output(3, 151) <= input(9);
output(3, 152) <= input(10);
output(3, 153) <= input(11);
output(3, 154) <= input(12);
output(3, 155) <= input(13);
output(3, 156) <= input(14);
output(3, 157) <= input(15);
output(3, 158) <= input(39);
output(3, 159) <= input(40);
output(3, 160) <= input(2);
output(3, 161) <= input(3);
output(3, 162) <= input(4);
output(3, 163) <= input(5);
output(3, 164) <= input(6);
output(3, 165) <= input(7);
output(3, 166) <= input(8);
output(3, 167) <= input(9);
output(3, 168) <= input(10);
output(3, 169) <= input(11);
output(3, 170) <= input(12);
output(3, 171) <= input(13);
output(3, 172) <= input(14);
output(3, 173) <= input(15);
output(3, 174) <= input(39);
output(3, 175) <= input(40);
output(3, 176) <= input(2);
output(3, 177) <= input(3);
output(3, 178) <= input(4);
output(3, 179) <= input(5);
output(3, 180) <= input(6);
output(3, 181) <= input(7);
output(3, 182) <= input(8);
output(3, 183) <= input(9);
output(3, 184) <= input(10);
output(3, 185) <= input(11);
output(3, 186) <= input(12);
output(3, 187) <= input(13);
output(3, 188) <= input(14);
output(3, 189) <= input(15);
output(3, 190) <= input(39);
output(3, 191) <= input(40);
output(3, 192) <= input(2);
output(3, 193) <= input(3);
output(3, 194) <= input(4);
output(3, 195) <= input(5);
output(3, 196) <= input(6);
output(3, 197) <= input(7);
output(3, 198) <= input(8);
output(3, 199) <= input(9);
output(3, 200) <= input(10);
output(3, 201) <= input(11);
output(3, 202) <= input(12);
output(3, 203) <= input(13);
output(3, 204) <= input(14);
output(3, 205) <= input(15);
output(3, 206) <= input(39);
output(3, 207) <= input(40);
output(3, 208) <= input(2);
output(3, 209) <= input(3);
output(3, 210) <= input(4);
output(3, 211) <= input(5);
output(3, 212) <= input(6);
output(3, 213) <= input(7);
output(3, 214) <= input(8);
output(3, 215) <= input(9);
output(3, 216) <= input(10);
output(3, 217) <= input(11);
output(3, 218) <= input(12);
output(3, 219) <= input(13);
output(3, 220) <= input(14);
output(3, 221) <= input(15);
output(3, 222) <= input(39);
output(3, 223) <= input(40);
output(3, 224) <= input(2);
output(3, 225) <= input(3);
output(3, 226) <= input(4);
output(3, 227) <= input(5);
output(3, 228) <= input(6);
output(3, 229) <= input(7);
output(3, 230) <= input(8);
output(3, 231) <= input(9);
output(3, 232) <= input(10);
output(3, 233) <= input(11);
output(3, 234) <= input(12);
output(3, 235) <= input(13);
output(3, 236) <= input(14);
output(3, 237) <= input(15);
output(3, 238) <= input(39);
output(3, 239) <= input(40);
output(3, 240) <= input(2);
output(3, 241) <= input(3);
output(3, 242) <= input(4);
output(3, 243) <= input(5);
output(3, 244) <= input(6);
output(3, 245) <= input(7);
output(3, 246) <= input(8);
output(3, 247) <= input(9);
output(3, 248) <= input(10);
output(3, 249) <= input(11);
output(3, 250) <= input(12);
output(3, 251) <= input(13);
output(3, 252) <= input(14);
output(3, 253) <= input(15);
output(3, 254) <= input(39);
output(3, 255) <= input(40);
output(4, 0) <= input(19);
output(4, 1) <= input(20);
output(4, 2) <= input(21);
output(4, 3) <= input(22);
output(4, 4) <= input(23);
output(4, 5) <= input(24);
output(4, 6) <= input(25);
output(4, 7) <= input(26);
output(4, 8) <= input(27);
output(4, 9) <= input(28);
output(4, 10) <= input(29);
output(4, 11) <= input(30);
output(4, 12) <= input(31);
output(4, 13) <= input(35);
output(4, 14) <= input(41);
output(4, 15) <= input(42);
output(4, 16) <= input(19);
output(4, 17) <= input(20);
output(4, 18) <= input(21);
output(4, 19) <= input(22);
output(4, 20) <= input(23);
output(4, 21) <= input(24);
output(4, 22) <= input(25);
output(4, 23) <= input(26);
output(4, 24) <= input(27);
output(4, 25) <= input(28);
output(4, 26) <= input(29);
output(4, 27) <= input(30);
output(4, 28) <= input(31);
output(4, 29) <= input(35);
output(4, 30) <= input(41);
output(4, 31) <= input(42);
output(4, 32) <= input(19);
output(4, 33) <= input(20);
output(4, 34) <= input(21);
output(4, 35) <= input(22);
output(4, 36) <= input(23);
output(4, 37) <= input(24);
output(4, 38) <= input(25);
output(4, 39) <= input(26);
output(4, 40) <= input(27);
output(4, 41) <= input(28);
output(4, 42) <= input(29);
output(4, 43) <= input(30);
output(4, 44) <= input(31);
output(4, 45) <= input(35);
output(4, 46) <= input(41);
output(4, 47) <= input(42);
output(4, 48) <= input(19);
output(4, 49) <= input(20);
output(4, 50) <= input(21);
output(4, 51) <= input(22);
output(4, 52) <= input(23);
output(4, 53) <= input(24);
output(4, 54) <= input(25);
output(4, 55) <= input(26);
output(4, 56) <= input(27);
output(4, 57) <= input(28);
output(4, 58) <= input(29);
output(4, 59) <= input(30);
output(4, 60) <= input(31);
output(4, 61) <= input(35);
output(4, 62) <= input(41);
output(4, 63) <= input(42);
output(4, 64) <= input(19);
output(4, 65) <= input(20);
output(4, 66) <= input(21);
output(4, 67) <= input(22);
output(4, 68) <= input(23);
output(4, 69) <= input(24);
output(4, 70) <= input(25);
output(4, 71) <= input(26);
output(4, 72) <= input(27);
output(4, 73) <= input(28);
output(4, 74) <= input(29);
output(4, 75) <= input(30);
output(4, 76) <= input(31);
output(4, 77) <= input(35);
output(4, 78) <= input(41);
output(4, 79) <= input(42);
output(4, 80) <= input(19);
output(4, 81) <= input(20);
output(4, 82) <= input(21);
output(4, 83) <= input(22);
output(4, 84) <= input(23);
output(4, 85) <= input(24);
output(4, 86) <= input(25);
output(4, 87) <= input(26);
output(4, 88) <= input(27);
output(4, 89) <= input(28);
output(4, 90) <= input(29);
output(4, 91) <= input(30);
output(4, 92) <= input(31);
output(4, 93) <= input(35);
output(4, 94) <= input(41);
output(4, 95) <= input(42);
output(4, 96) <= input(19);
output(4, 97) <= input(20);
output(4, 98) <= input(21);
output(4, 99) <= input(22);
output(4, 100) <= input(23);
output(4, 101) <= input(24);
output(4, 102) <= input(25);
output(4, 103) <= input(26);
output(4, 104) <= input(27);
output(4, 105) <= input(28);
output(4, 106) <= input(29);
output(4, 107) <= input(30);
output(4, 108) <= input(31);
output(4, 109) <= input(35);
output(4, 110) <= input(41);
output(4, 111) <= input(42);
output(4, 112) <= input(19);
output(4, 113) <= input(20);
output(4, 114) <= input(21);
output(4, 115) <= input(22);
output(4, 116) <= input(23);
output(4, 117) <= input(24);
output(4, 118) <= input(25);
output(4, 119) <= input(26);
output(4, 120) <= input(27);
output(4, 121) <= input(28);
output(4, 122) <= input(29);
output(4, 123) <= input(30);
output(4, 124) <= input(31);
output(4, 125) <= input(35);
output(4, 126) <= input(41);
output(4, 127) <= input(42);
output(4, 128) <= input(19);
output(4, 129) <= input(20);
output(4, 130) <= input(21);
output(4, 131) <= input(22);
output(4, 132) <= input(23);
output(4, 133) <= input(24);
output(4, 134) <= input(25);
output(4, 135) <= input(26);
output(4, 136) <= input(27);
output(4, 137) <= input(28);
output(4, 138) <= input(29);
output(4, 139) <= input(30);
output(4, 140) <= input(31);
output(4, 141) <= input(35);
output(4, 142) <= input(41);
output(4, 143) <= input(42);
output(4, 144) <= input(19);
output(4, 145) <= input(20);
output(4, 146) <= input(21);
output(4, 147) <= input(22);
output(4, 148) <= input(23);
output(4, 149) <= input(24);
output(4, 150) <= input(25);
output(4, 151) <= input(26);
output(4, 152) <= input(27);
output(4, 153) <= input(28);
output(4, 154) <= input(29);
output(4, 155) <= input(30);
output(4, 156) <= input(31);
output(4, 157) <= input(35);
output(4, 158) <= input(41);
output(4, 159) <= input(42);
output(4, 160) <= input(19);
output(4, 161) <= input(20);
output(4, 162) <= input(21);
output(4, 163) <= input(22);
output(4, 164) <= input(23);
output(4, 165) <= input(24);
output(4, 166) <= input(25);
output(4, 167) <= input(26);
output(4, 168) <= input(27);
output(4, 169) <= input(28);
output(4, 170) <= input(29);
output(4, 171) <= input(30);
output(4, 172) <= input(31);
output(4, 173) <= input(35);
output(4, 174) <= input(41);
output(4, 175) <= input(42);
output(4, 176) <= input(19);
output(4, 177) <= input(20);
output(4, 178) <= input(21);
output(4, 179) <= input(22);
output(4, 180) <= input(23);
output(4, 181) <= input(24);
output(4, 182) <= input(25);
output(4, 183) <= input(26);
output(4, 184) <= input(27);
output(4, 185) <= input(28);
output(4, 186) <= input(29);
output(4, 187) <= input(30);
output(4, 188) <= input(31);
output(4, 189) <= input(35);
output(4, 190) <= input(41);
output(4, 191) <= input(42);
output(4, 192) <= input(19);
output(4, 193) <= input(20);
output(4, 194) <= input(21);
output(4, 195) <= input(22);
output(4, 196) <= input(23);
output(4, 197) <= input(24);
output(4, 198) <= input(25);
output(4, 199) <= input(26);
output(4, 200) <= input(27);
output(4, 201) <= input(28);
output(4, 202) <= input(29);
output(4, 203) <= input(30);
output(4, 204) <= input(31);
output(4, 205) <= input(35);
output(4, 206) <= input(41);
output(4, 207) <= input(42);
output(4, 208) <= input(19);
output(4, 209) <= input(20);
output(4, 210) <= input(21);
output(4, 211) <= input(22);
output(4, 212) <= input(23);
output(4, 213) <= input(24);
output(4, 214) <= input(25);
output(4, 215) <= input(26);
output(4, 216) <= input(27);
output(4, 217) <= input(28);
output(4, 218) <= input(29);
output(4, 219) <= input(30);
output(4, 220) <= input(31);
output(4, 221) <= input(35);
output(4, 222) <= input(41);
output(4, 223) <= input(42);
output(4, 224) <= input(19);
output(4, 225) <= input(20);
output(4, 226) <= input(21);
output(4, 227) <= input(22);
output(4, 228) <= input(23);
output(4, 229) <= input(24);
output(4, 230) <= input(25);
output(4, 231) <= input(26);
output(4, 232) <= input(27);
output(4, 233) <= input(28);
output(4, 234) <= input(29);
output(4, 235) <= input(30);
output(4, 236) <= input(31);
output(4, 237) <= input(35);
output(4, 238) <= input(41);
output(4, 239) <= input(42);
output(4, 240) <= input(3);
output(4, 241) <= input(4);
output(4, 242) <= input(5);
output(4, 243) <= input(6);
output(4, 244) <= input(7);
output(4, 245) <= input(8);
output(4, 246) <= input(9);
output(4, 247) <= input(10);
output(4, 248) <= input(11);
output(4, 249) <= input(12);
output(4, 250) <= input(13);
output(4, 251) <= input(14);
output(4, 252) <= input(15);
output(4, 253) <= input(39);
output(4, 254) <= input(40);
output(4, 255) <= input(43);
output(5, 0) <= input(3);
output(5, 1) <= input(4);
output(5, 2) <= input(5);
output(5, 3) <= input(6);
output(5, 4) <= input(7);
output(5, 5) <= input(8);
output(5, 6) <= input(9);
output(5, 7) <= input(10);
output(5, 8) <= input(11);
output(5, 9) <= input(12);
output(5, 10) <= input(13);
output(5, 11) <= input(14);
output(5, 12) <= input(15);
output(5, 13) <= input(39);
output(5, 14) <= input(40);
output(5, 15) <= input(43);
output(5, 16) <= input(3);
output(5, 17) <= input(4);
output(5, 18) <= input(5);
output(5, 19) <= input(6);
output(5, 20) <= input(7);
output(5, 21) <= input(8);
output(5, 22) <= input(9);
output(5, 23) <= input(10);
output(5, 24) <= input(11);
output(5, 25) <= input(12);
output(5, 26) <= input(13);
output(5, 27) <= input(14);
output(5, 28) <= input(15);
output(5, 29) <= input(39);
output(5, 30) <= input(40);
output(5, 31) <= input(43);
output(5, 32) <= input(3);
output(5, 33) <= input(4);
output(5, 34) <= input(5);
output(5, 35) <= input(6);
output(5, 36) <= input(7);
output(5, 37) <= input(8);
output(5, 38) <= input(9);
output(5, 39) <= input(10);
output(5, 40) <= input(11);
output(5, 41) <= input(12);
output(5, 42) <= input(13);
output(5, 43) <= input(14);
output(5, 44) <= input(15);
output(5, 45) <= input(39);
output(5, 46) <= input(40);
output(5, 47) <= input(43);
output(5, 48) <= input(3);
output(5, 49) <= input(4);
output(5, 50) <= input(5);
output(5, 51) <= input(6);
output(5, 52) <= input(7);
output(5, 53) <= input(8);
output(5, 54) <= input(9);
output(5, 55) <= input(10);
output(5, 56) <= input(11);
output(5, 57) <= input(12);
output(5, 58) <= input(13);
output(5, 59) <= input(14);
output(5, 60) <= input(15);
output(5, 61) <= input(39);
output(5, 62) <= input(40);
output(5, 63) <= input(43);
output(5, 64) <= input(3);
output(5, 65) <= input(4);
output(5, 66) <= input(5);
output(5, 67) <= input(6);
output(5, 68) <= input(7);
output(5, 69) <= input(8);
output(5, 70) <= input(9);
output(5, 71) <= input(10);
output(5, 72) <= input(11);
output(5, 73) <= input(12);
output(5, 74) <= input(13);
output(5, 75) <= input(14);
output(5, 76) <= input(15);
output(5, 77) <= input(39);
output(5, 78) <= input(40);
output(5, 79) <= input(43);
output(5, 80) <= input(3);
output(5, 81) <= input(4);
output(5, 82) <= input(5);
output(5, 83) <= input(6);
output(5, 84) <= input(7);
output(5, 85) <= input(8);
output(5, 86) <= input(9);
output(5, 87) <= input(10);
output(5, 88) <= input(11);
output(5, 89) <= input(12);
output(5, 90) <= input(13);
output(5, 91) <= input(14);
output(5, 92) <= input(15);
output(5, 93) <= input(39);
output(5, 94) <= input(40);
output(5, 95) <= input(43);
output(5, 96) <= input(3);
output(5, 97) <= input(4);
output(5, 98) <= input(5);
output(5, 99) <= input(6);
output(5, 100) <= input(7);
output(5, 101) <= input(8);
output(5, 102) <= input(9);
output(5, 103) <= input(10);
output(5, 104) <= input(11);
output(5, 105) <= input(12);
output(5, 106) <= input(13);
output(5, 107) <= input(14);
output(5, 108) <= input(15);
output(5, 109) <= input(39);
output(5, 110) <= input(40);
output(5, 111) <= input(43);
output(5, 112) <= input(20);
output(5, 113) <= input(21);
output(5, 114) <= input(22);
output(5, 115) <= input(23);
output(5, 116) <= input(24);
output(5, 117) <= input(25);
output(5, 118) <= input(26);
output(5, 119) <= input(27);
output(5, 120) <= input(28);
output(5, 121) <= input(29);
output(5, 122) <= input(30);
output(5, 123) <= input(31);
output(5, 124) <= input(35);
output(5, 125) <= input(41);
output(5, 126) <= input(42);
output(5, 127) <= input(44);
output(5, 128) <= input(20);
output(5, 129) <= input(21);
output(5, 130) <= input(22);
output(5, 131) <= input(23);
output(5, 132) <= input(24);
output(5, 133) <= input(25);
output(5, 134) <= input(26);
output(5, 135) <= input(27);
output(5, 136) <= input(28);
output(5, 137) <= input(29);
output(5, 138) <= input(30);
output(5, 139) <= input(31);
output(5, 140) <= input(35);
output(5, 141) <= input(41);
output(5, 142) <= input(42);
output(5, 143) <= input(44);
output(5, 144) <= input(20);
output(5, 145) <= input(21);
output(5, 146) <= input(22);
output(5, 147) <= input(23);
output(5, 148) <= input(24);
output(5, 149) <= input(25);
output(5, 150) <= input(26);
output(5, 151) <= input(27);
output(5, 152) <= input(28);
output(5, 153) <= input(29);
output(5, 154) <= input(30);
output(5, 155) <= input(31);
output(5, 156) <= input(35);
output(5, 157) <= input(41);
output(5, 158) <= input(42);
output(5, 159) <= input(44);
output(5, 160) <= input(20);
output(5, 161) <= input(21);
output(5, 162) <= input(22);
output(5, 163) <= input(23);
output(5, 164) <= input(24);
output(5, 165) <= input(25);
output(5, 166) <= input(26);
output(5, 167) <= input(27);
output(5, 168) <= input(28);
output(5, 169) <= input(29);
output(5, 170) <= input(30);
output(5, 171) <= input(31);
output(5, 172) <= input(35);
output(5, 173) <= input(41);
output(5, 174) <= input(42);
output(5, 175) <= input(44);
output(5, 176) <= input(20);
output(5, 177) <= input(21);
output(5, 178) <= input(22);
output(5, 179) <= input(23);
output(5, 180) <= input(24);
output(5, 181) <= input(25);
output(5, 182) <= input(26);
output(5, 183) <= input(27);
output(5, 184) <= input(28);
output(5, 185) <= input(29);
output(5, 186) <= input(30);
output(5, 187) <= input(31);
output(5, 188) <= input(35);
output(5, 189) <= input(41);
output(5, 190) <= input(42);
output(5, 191) <= input(44);
output(5, 192) <= input(20);
output(5, 193) <= input(21);
output(5, 194) <= input(22);
output(5, 195) <= input(23);
output(5, 196) <= input(24);
output(5, 197) <= input(25);
output(5, 198) <= input(26);
output(5, 199) <= input(27);
output(5, 200) <= input(28);
output(5, 201) <= input(29);
output(5, 202) <= input(30);
output(5, 203) <= input(31);
output(5, 204) <= input(35);
output(5, 205) <= input(41);
output(5, 206) <= input(42);
output(5, 207) <= input(44);
output(5, 208) <= input(20);
output(5, 209) <= input(21);
output(5, 210) <= input(22);
output(5, 211) <= input(23);
output(5, 212) <= input(24);
output(5, 213) <= input(25);
output(5, 214) <= input(26);
output(5, 215) <= input(27);
output(5, 216) <= input(28);
output(5, 217) <= input(29);
output(5, 218) <= input(30);
output(5, 219) <= input(31);
output(5, 220) <= input(35);
output(5, 221) <= input(41);
output(5, 222) <= input(42);
output(5, 223) <= input(44);
output(5, 224) <= input(20);
output(5, 225) <= input(21);
output(5, 226) <= input(22);
output(5, 227) <= input(23);
output(5, 228) <= input(24);
output(5, 229) <= input(25);
output(5, 230) <= input(26);
output(5, 231) <= input(27);
output(5, 232) <= input(28);
output(5, 233) <= input(29);
output(5, 234) <= input(30);
output(5, 235) <= input(31);
output(5, 236) <= input(35);
output(5, 237) <= input(41);
output(5, 238) <= input(42);
output(5, 239) <= input(44);
output(5, 240) <= input(4);
output(5, 241) <= input(5);
output(5, 242) <= input(6);
output(5, 243) <= input(7);
output(5, 244) <= input(8);
output(5, 245) <= input(9);
output(5, 246) <= input(10);
output(5, 247) <= input(11);
output(5, 248) <= input(12);
output(5, 249) <= input(13);
output(5, 250) <= input(14);
output(5, 251) <= input(15);
output(5, 252) <= input(39);
output(5, 253) <= input(40);
output(5, 254) <= input(43);
output(5, 255) <= input(45);
output(6, 0) <= input(20);
output(6, 1) <= input(21);
output(6, 2) <= input(22);
output(6, 3) <= input(23);
output(6, 4) <= input(24);
output(6, 5) <= input(25);
output(6, 6) <= input(26);
output(6, 7) <= input(27);
output(6, 8) <= input(28);
output(6, 9) <= input(29);
output(6, 10) <= input(30);
output(6, 11) <= input(31);
output(6, 12) <= input(35);
output(6, 13) <= input(41);
output(6, 14) <= input(42);
output(6, 15) <= input(44);
output(6, 16) <= input(20);
output(6, 17) <= input(21);
output(6, 18) <= input(22);
output(6, 19) <= input(23);
output(6, 20) <= input(24);
output(6, 21) <= input(25);
output(6, 22) <= input(26);
output(6, 23) <= input(27);
output(6, 24) <= input(28);
output(6, 25) <= input(29);
output(6, 26) <= input(30);
output(6, 27) <= input(31);
output(6, 28) <= input(35);
output(6, 29) <= input(41);
output(6, 30) <= input(42);
output(6, 31) <= input(44);
output(6, 32) <= input(20);
output(6, 33) <= input(21);
output(6, 34) <= input(22);
output(6, 35) <= input(23);
output(6, 36) <= input(24);
output(6, 37) <= input(25);
output(6, 38) <= input(26);
output(6, 39) <= input(27);
output(6, 40) <= input(28);
output(6, 41) <= input(29);
output(6, 42) <= input(30);
output(6, 43) <= input(31);
output(6, 44) <= input(35);
output(6, 45) <= input(41);
output(6, 46) <= input(42);
output(6, 47) <= input(44);
output(6, 48) <= input(20);
output(6, 49) <= input(21);
output(6, 50) <= input(22);
output(6, 51) <= input(23);
output(6, 52) <= input(24);
output(6, 53) <= input(25);
output(6, 54) <= input(26);
output(6, 55) <= input(27);
output(6, 56) <= input(28);
output(6, 57) <= input(29);
output(6, 58) <= input(30);
output(6, 59) <= input(31);
output(6, 60) <= input(35);
output(6, 61) <= input(41);
output(6, 62) <= input(42);
output(6, 63) <= input(44);
output(6, 64) <= input(20);
output(6, 65) <= input(21);
output(6, 66) <= input(22);
output(6, 67) <= input(23);
output(6, 68) <= input(24);
output(6, 69) <= input(25);
output(6, 70) <= input(26);
output(6, 71) <= input(27);
output(6, 72) <= input(28);
output(6, 73) <= input(29);
output(6, 74) <= input(30);
output(6, 75) <= input(31);
output(6, 76) <= input(35);
output(6, 77) <= input(41);
output(6, 78) <= input(42);
output(6, 79) <= input(44);
output(6, 80) <= input(4);
output(6, 81) <= input(5);
output(6, 82) <= input(6);
output(6, 83) <= input(7);
output(6, 84) <= input(8);
output(6, 85) <= input(9);
output(6, 86) <= input(10);
output(6, 87) <= input(11);
output(6, 88) <= input(12);
output(6, 89) <= input(13);
output(6, 90) <= input(14);
output(6, 91) <= input(15);
output(6, 92) <= input(39);
output(6, 93) <= input(40);
output(6, 94) <= input(43);
output(6, 95) <= input(45);
output(6, 96) <= input(4);
output(6, 97) <= input(5);
output(6, 98) <= input(6);
output(6, 99) <= input(7);
output(6, 100) <= input(8);
output(6, 101) <= input(9);
output(6, 102) <= input(10);
output(6, 103) <= input(11);
output(6, 104) <= input(12);
output(6, 105) <= input(13);
output(6, 106) <= input(14);
output(6, 107) <= input(15);
output(6, 108) <= input(39);
output(6, 109) <= input(40);
output(6, 110) <= input(43);
output(6, 111) <= input(45);
output(6, 112) <= input(4);
output(6, 113) <= input(5);
output(6, 114) <= input(6);
output(6, 115) <= input(7);
output(6, 116) <= input(8);
output(6, 117) <= input(9);
output(6, 118) <= input(10);
output(6, 119) <= input(11);
output(6, 120) <= input(12);
output(6, 121) <= input(13);
output(6, 122) <= input(14);
output(6, 123) <= input(15);
output(6, 124) <= input(39);
output(6, 125) <= input(40);
output(6, 126) <= input(43);
output(6, 127) <= input(45);
output(6, 128) <= input(4);
output(6, 129) <= input(5);
output(6, 130) <= input(6);
output(6, 131) <= input(7);
output(6, 132) <= input(8);
output(6, 133) <= input(9);
output(6, 134) <= input(10);
output(6, 135) <= input(11);
output(6, 136) <= input(12);
output(6, 137) <= input(13);
output(6, 138) <= input(14);
output(6, 139) <= input(15);
output(6, 140) <= input(39);
output(6, 141) <= input(40);
output(6, 142) <= input(43);
output(6, 143) <= input(45);
output(6, 144) <= input(4);
output(6, 145) <= input(5);
output(6, 146) <= input(6);
output(6, 147) <= input(7);
output(6, 148) <= input(8);
output(6, 149) <= input(9);
output(6, 150) <= input(10);
output(6, 151) <= input(11);
output(6, 152) <= input(12);
output(6, 153) <= input(13);
output(6, 154) <= input(14);
output(6, 155) <= input(15);
output(6, 156) <= input(39);
output(6, 157) <= input(40);
output(6, 158) <= input(43);
output(6, 159) <= input(45);
output(6, 160) <= input(21);
output(6, 161) <= input(22);
output(6, 162) <= input(23);
output(6, 163) <= input(24);
output(6, 164) <= input(25);
output(6, 165) <= input(26);
output(6, 166) <= input(27);
output(6, 167) <= input(28);
output(6, 168) <= input(29);
output(6, 169) <= input(30);
output(6, 170) <= input(31);
output(6, 171) <= input(35);
output(6, 172) <= input(41);
output(6, 173) <= input(42);
output(6, 174) <= input(44);
output(6, 175) <= input(46);
output(6, 176) <= input(21);
output(6, 177) <= input(22);
output(6, 178) <= input(23);
output(6, 179) <= input(24);
output(6, 180) <= input(25);
output(6, 181) <= input(26);
output(6, 182) <= input(27);
output(6, 183) <= input(28);
output(6, 184) <= input(29);
output(6, 185) <= input(30);
output(6, 186) <= input(31);
output(6, 187) <= input(35);
output(6, 188) <= input(41);
output(6, 189) <= input(42);
output(6, 190) <= input(44);
output(6, 191) <= input(46);
output(6, 192) <= input(21);
output(6, 193) <= input(22);
output(6, 194) <= input(23);
output(6, 195) <= input(24);
output(6, 196) <= input(25);
output(6, 197) <= input(26);
output(6, 198) <= input(27);
output(6, 199) <= input(28);
output(6, 200) <= input(29);
output(6, 201) <= input(30);
output(6, 202) <= input(31);
output(6, 203) <= input(35);
output(6, 204) <= input(41);
output(6, 205) <= input(42);
output(6, 206) <= input(44);
output(6, 207) <= input(46);
output(6, 208) <= input(21);
output(6, 209) <= input(22);
output(6, 210) <= input(23);
output(6, 211) <= input(24);
output(6, 212) <= input(25);
output(6, 213) <= input(26);
output(6, 214) <= input(27);
output(6, 215) <= input(28);
output(6, 216) <= input(29);
output(6, 217) <= input(30);
output(6, 218) <= input(31);
output(6, 219) <= input(35);
output(6, 220) <= input(41);
output(6, 221) <= input(42);
output(6, 222) <= input(44);
output(6, 223) <= input(46);
output(6, 224) <= input(21);
output(6, 225) <= input(22);
output(6, 226) <= input(23);
output(6, 227) <= input(24);
output(6, 228) <= input(25);
output(6, 229) <= input(26);
output(6, 230) <= input(27);
output(6, 231) <= input(28);
output(6, 232) <= input(29);
output(6, 233) <= input(30);
output(6, 234) <= input(31);
output(6, 235) <= input(35);
output(6, 236) <= input(41);
output(6, 237) <= input(42);
output(6, 238) <= input(44);
output(6, 239) <= input(46);
output(6, 240) <= input(5);
output(6, 241) <= input(6);
output(6, 242) <= input(7);
output(6, 243) <= input(8);
output(6, 244) <= input(9);
output(6, 245) <= input(10);
output(6, 246) <= input(11);
output(6, 247) <= input(12);
output(6, 248) <= input(13);
output(6, 249) <= input(14);
output(6, 250) <= input(15);
output(6, 251) <= input(39);
output(6, 252) <= input(40);
output(6, 253) <= input(43);
output(6, 254) <= input(45);
output(6, 255) <= input(47);
output(7, 0) <= input(4);
output(7, 1) <= input(5);
output(7, 2) <= input(6);
output(7, 3) <= input(7);
output(7, 4) <= input(8);
output(7, 5) <= input(9);
output(7, 6) <= input(10);
output(7, 7) <= input(11);
output(7, 8) <= input(12);
output(7, 9) <= input(13);
output(7, 10) <= input(14);
output(7, 11) <= input(15);
output(7, 12) <= input(39);
output(7, 13) <= input(40);
output(7, 14) <= input(43);
output(7, 15) <= input(45);
output(7, 16) <= input(4);
output(7, 17) <= input(5);
output(7, 18) <= input(6);
output(7, 19) <= input(7);
output(7, 20) <= input(8);
output(7, 21) <= input(9);
output(7, 22) <= input(10);
output(7, 23) <= input(11);
output(7, 24) <= input(12);
output(7, 25) <= input(13);
output(7, 26) <= input(14);
output(7, 27) <= input(15);
output(7, 28) <= input(39);
output(7, 29) <= input(40);
output(7, 30) <= input(43);
output(7, 31) <= input(45);
output(7, 32) <= input(4);
output(7, 33) <= input(5);
output(7, 34) <= input(6);
output(7, 35) <= input(7);
output(7, 36) <= input(8);
output(7, 37) <= input(9);
output(7, 38) <= input(10);
output(7, 39) <= input(11);
output(7, 40) <= input(12);
output(7, 41) <= input(13);
output(7, 42) <= input(14);
output(7, 43) <= input(15);
output(7, 44) <= input(39);
output(7, 45) <= input(40);
output(7, 46) <= input(43);
output(7, 47) <= input(45);
output(7, 48) <= input(21);
output(7, 49) <= input(22);
output(7, 50) <= input(23);
output(7, 51) <= input(24);
output(7, 52) <= input(25);
output(7, 53) <= input(26);
output(7, 54) <= input(27);
output(7, 55) <= input(28);
output(7, 56) <= input(29);
output(7, 57) <= input(30);
output(7, 58) <= input(31);
output(7, 59) <= input(35);
output(7, 60) <= input(41);
output(7, 61) <= input(42);
output(7, 62) <= input(44);
output(7, 63) <= input(46);
output(7, 64) <= input(21);
output(7, 65) <= input(22);
output(7, 66) <= input(23);
output(7, 67) <= input(24);
output(7, 68) <= input(25);
output(7, 69) <= input(26);
output(7, 70) <= input(27);
output(7, 71) <= input(28);
output(7, 72) <= input(29);
output(7, 73) <= input(30);
output(7, 74) <= input(31);
output(7, 75) <= input(35);
output(7, 76) <= input(41);
output(7, 77) <= input(42);
output(7, 78) <= input(44);
output(7, 79) <= input(46);
output(7, 80) <= input(21);
output(7, 81) <= input(22);
output(7, 82) <= input(23);
output(7, 83) <= input(24);
output(7, 84) <= input(25);
output(7, 85) <= input(26);
output(7, 86) <= input(27);
output(7, 87) <= input(28);
output(7, 88) <= input(29);
output(7, 89) <= input(30);
output(7, 90) <= input(31);
output(7, 91) <= input(35);
output(7, 92) <= input(41);
output(7, 93) <= input(42);
output(7, 94) <= input(44);
output(7, 95) <= input(46);
output(7, 96) <= input(21);
output(7, 97) <= input(22);
output(7, 98) <= input(23);
output(7, 99) <= input(24);
output(7, 100) <= input(25);
output(7, 101) <= input(26);
output(7, 102) <= input(27);
output(7, 103) <= input(28);
output(7, 104) <= input(29);
output(7, 105) <= input(30);
output(7, 106) <= input(31);
output(7, 107) <= input(35);
output(7, 108) <= input(41);
output(7, 109) <= input(42);
output(7, 110) <= input(44);
output(7, 111) <= input(46);
output(7, 112) <= input(5);
output(7, 113) <= input(6);
output(7, 114) <= input(7);
output(7, 115) <= input(8);
output(7, 116) <= input(9);
output(7, 117) <= input(10);
output(7, 118) <= input(11);
output(7, 119) <= input(12);
output(7, 120) <= input(13);
output(7, 121) <= input(14);
output(7, 122) <= input(15);
output(7, 123) <= input(39);
output(7, 124) <= input(40);
output(7, 125) <= input(43);
output(7, 126) <= input(45);
output(7, 127) <= input(47);
output(7, 128) <= input(5);
output(7, 129) <= input(6);
output(7, 130) <= input(7);
output(7, 131) <= input(8);
output(7, 132) <= input(9);
output(7, 133) <= input(10);
output(7, 134) <= input(11);
output(7, 135) <= input(12);
output(7, 136) <= input(13);
output(7, 137) <= input(14);
output(7, 138) <= input(15);
output(7, 139) <= input(39);
output(7, 140) <= input(40);
output(7, 141) <= input(43);
output(7, 142) <= input(45);
output(7, 143) <= input(47);
output(7, 144) <= input(5);
output(7, 145) <= input(6);
output(7, 146) <= input(7);
output(7, 147) <= input(8);
output(7, 148) <= input(9);
output(7, 149) <= input(10);
output(7, 150) <= input(11);
output(7, 151) <= input(12);
output(7, 152) <= input(13);
output(7, 153) <= input(14);
output(7, 154) <= input(15);
output(7, 155) <= input(39);
output(7, 156) <= input(40);
output(7, 157) <= input(43);
output(7, 158) <= input(45);
output(7, 159) <= input(47);
output(7, 160) <= input(5);
output(7, 161) <= input(6);
output(7, 162) <= input(7);
output(7, 163) <= input(8);
output(7, 164) <= input(9);
output(7, 165) <= input(10);
output(7, 166) <= input(11);
output(7, 167) <= input(12);
output(7, 168) <= input(13);
output(7, 169) <= input(14);
output(7, 170) <= input(15);
output(7, 171) <= input(39);
output(7, 172) <= input(40);
output(7, 173) <= input(43);
output(7, 174) <= input(45);
output(7, 175) <= input(47);
output(7, 176) <= input(22);
output(7, 177) <= input(23);
output(7, 178) <= input(24);
output(7, 179) <= input(25);
output(7, 180) <= input(26);
output(7, 181) <= input(27);
output(7, 182) <= input(28);
output(7, 183) <= input(29);
output(7, 184) <= input(30);
output(7, 185) <= input(31);
output(7, 186) <= input(35);
output(7, 187) <= input(41);
output(7, 188) <= input(42);
output(7, 189) <= input(44);
output(7, 190) <= input(46);
output(7, 191) <= input(48);
output(7, 192) <= input(22);
output(7, 193) <= input(23);
output(7, 194) <= input(24);
output(7, 195) <= input(25);
output(7, 196) <= input(26);
output(7, 197) <= input(27);
output(7, 198) <= input(28);
output(7, 199) <= input(29);
output(7, 200) <= input(30);
output(7, 201) <= input(31);
output(7, 202) <= input(35);
output(7, 203) <= input(41);
output(7, 204) <= input(42);
output(7, 205) <= input(44);
output(7, 206) <= input(46);
output(7, 207) <= input(48);
output(7, 208) <= input(22);
output(7, 209) <= input(23);
output(7, 210) <= input(24);
output(7, 211) <= input(25);
output(7, 212) <= input(26);
output(7, 213) <= input(27);
output(7, 214) <= input(28);
output(7, 215) <= input(29);
output(7, 216) <= input(30);
output(7, 217) <= input(31);
output(7, 218) <= input(35);
output(7, 219) <= input(41);
output(7, 220) <= input(42);
output(7, 221) <= input(44);
output(7, 222) <= input(46);
output(7, 223) <= input(48);
output(7, 224) <= input(22);
output(7, 225) <= input(23);
output(7, 226) <= input(24);
output(7, 227) <= input(25);
output(7, 228) <= input(26);
output(7, 229) <= input(27);
output(7, 230) <= input(28);
output(7, 231) <= input(29);
output(7, 232) <= input(30);
output(7, 233) <= input(31);
output(7, 234) <= input(35);
output(7, 235) <= input(41);
output(7, 236) <= input(42);
output(7, 237) <= input(44);
output(7, 238) <= input(46);
output(7, 239) <= input(48);
output(7, 240) <= input(6);
output(7, 241) <= input(7);
output(7, 242) <= input(8);
output(7, 243) <= input(9);
output(7, 244) <= input(10);
output(7, 245) <= input(11);
output(7, 246) <= input(12);
output(7, 247) <= input(13);
output(7, 248) <= input(14);
output(7, 249) <= input(15);
output(7, 250) <= input(39);
output(7, 251) <= input(40);
output(7, 252) <= input(43);
output(7, 253) <= input(45);
output(7, 254) <= input(47);
output(7, 255) <= input(49);
when "1110" =>
output(0, 0) <= input(0);
output(0, 1) <= input(1);
output(0, 2) <= input(2);
output(0, 3) <= input(3);
output(0, 4) <= input(4);
output(0, 5) <= input(5);
output(0, 6) <= input(6);
output(0, 7) <= input(7);
output(0, 8) <= input(8);
output(0, 9) <= input(9);
output(0, 10) <= input(10);
output(0, 11) <= input(11);
output(0, 12) <= input(12);
output(0, 13) <= input(13);
output(0, 14) <= input(14);
output(0, 15) <= input(15);
output(0, 16) <= input(0);
output(0, 17) <= input(1);
output(0, 18) <= input(2);
output(0, 19) <= input(3);
output(0, 20) <= input(4);
output(0, 21) <= input(5);
output(0, 22) <= input(6);
output(0, 23) <= input(7);
output(0, 24) <= input(8);
output(0, 25) <= input(9);
output(0, 26) <= input(10);
output(0, 27) <= input(11);
output(0, 28) <= input(12);
output(0, 29) <= input(13);
output(0, 30) <= input(14);
output(0, 31) <= input(15);
output(0, 32) <= input(16);
output(0, 33) <= input(17);
output(0, 34) <= input(18);
output(0, 35) <= input(19);
output(0, 36) <= input(20);
output(0, 37) <= input(21);
output(0, 38) <= input(22);
output(0, 39) <= input(23);
output(0, 40) <= input(24);
output(0, 41) <= input(25);
output(0, 42) <= input(26);
output(0, 43) <= input(27);
output(0, 44) <= input(28);
output(0, 45) <= input(29);
output(0, 46) <= input(30);
output(0, 47) <= input(31);
output(0, 48) <= input(16);
output(0, 49) <= input(17);
output(0, 50) <= input(18);
output(0, 51) <= input(19);
output(0, 52) <= input(20);
output(0, 53) <= input(21);
output(0, 54) <= input(22);
output(0, 55) <= input(23);
output(0, 56) <= input(24);
output(0, 57) <= input(25);
output(0, 58) <= input(26);
output(0, 59) <= input(27);
output(0, 60) <= input(28);
output(0, 61) <= input(29);
output(0, 62) <= input(30);
output(0, 63) <= input(31);
output(0, 64) <= input(16);
output(0, 65) <= input(17);
output(0, 66) <= input(18);
output(0, 67) <= input(19);
output(0, 68) <= input(20);
output(0, 69) <= input(21);
output(0, 70) <= input(22);
output(0, 71) <= input(23);
output(0, 72) <= input(24);
output(0, 73) <= input(25);
output(0, 74) <= input(26);
output(0, 75) <= input(27);
output(0, 76) <= input(28);
output(0, 77) <= input(29);
output(0, 78) <= input(30);
output(0, 79) <= input(31);
output(0, 80) <= input(1);
output(0, 81) <= input(2);
output(0, 82) <= input(3);
output(0, 83) <= input(4);
output(0, 84) <= input(5);
output(0, 85) <= input(6);
output(0, 86) <= input(7);
output(0, 87) <= input(8);
output(0, 88) <= input(9);
output(0, 89) <= input(10);
output(0, 90) <= input(11);
output(0, 91) <= input(12);
output(0, 92) <= input(13);
output(0, 93) <= input(14);
output(0, 94) <= input(15);
output(0, 95) <= input(32);
output(0, 96) <= input(1);
output(0, 97) <= input(2);
output(0, 98) <= input(3);
output(0, 99) <= input(4);
output(0, 100) <= input(5);
output(0, 101) <= input(6);
output(0, 102) <= input(7);
output(0, 103) <= input(8);
output(0, 104) <= input(9);
output(0, 105) <= input(10);
output(0, 106) <= input(11);
output(0, 107) <= input(12);
output(0, 108) <= input(13);
output(0, 109) <= input(14);
output(0, 110) <= input(15);
output(0, 111) <= input(32);
output(0, 112) <= input(17);
output(0, 113) <= input(18);
output(0, 114) <= input(19);
output(0, 115) <= input(20);
output(0, 116) <= input(21);
output(0, 117) <= input(22);
output(0, 118) <= input(23);
output(0, 119) <= input(24);
output(0, 120) <= input(25);
output(0, 121) <= input(26);
output(0, 122) <= input(27);
output(0, 123) <= input(28);
output(0, 124) <= input(29);
output(0, 125) <= input(30);
output(0, 126) <= input(31);
output(0, 127) <= input(33);
output(0, 128) <= input(17);
output(0, 129) <= input(18);
output(0, 130) <= input(19);
output(0, 131) <= input(20);
output(0, 132) <= input(21);
output(0, 133) <= input(22);
output(0, 134) <= input(23);
output(0, 135) <= input(24);
output(0, 136) <= input(25);
output(0, 137) <= input(26);
output(0, 138) <= input(27);
output(0, 139) <= input(28);
output(0, 140) <= input(29);
output(0, 141) <= input(30);
output(0, 142) <= input(31);
output(0, 143) <= input(33);
output(0, 144) <= input(17);
output(0, 145) <= input(18);
output(0, 146) <= input(19);
output(0, 147) <= input(20);
output(0, 148) <= input(21);
output(0, 149) <= input(22);
output(0, 150) <= input(23);
output(0, 151) <= input(24);
output(0, 152) <= input(25);
output(0, 153) <= input(26);
output(0, 154) <= input(27);
output(0, 155) <= input(28);
output(0, 156) <= input(29);
output(0, 157) <= input(30);
output(0, 158) <= input(31);
output(0, 159) <= input(33);
output(0, 160) <= input(2);
output(0, 161) <= input(3);
output(0, 162) <= input(4);
output(0, 163) <= input(5);
output(0, 164) <= input(6);
output(0, 165) <= input(7);
output(0, 166) <= input(8);
output(0, 167) <= input(9);
output(0, 168) <= input(10);
output(0, 169) <= input(11);
output(0, 170) <= input(12);
output(0, 171) <= input(13);
output(0, 172) <= input(14);
output(0, 173) <= input(15);
output(0, 174) <= input(32);
output(0, 175) <= input(34);
output(0, 176) <= input(2);
output(0, 177) <= input(3);
output(0, 178) <= input(4);
output(0, 179) <= input(5);
output(0, 180) <= input(6);
output(0, 181) <= input(7);
output(0, 182) <= input(8);
output(0, 183) <= input(9);
output(0, 184) <= input(10);
output(0, 185) <= input(11);
output(0, 186) <= input(12);
output(0, 187) <= input(13);
output(0, 188) <= input(14);
output(0, 189) <= input(15);
output(0, 190) <= input(32);
output(0, 191) <= input(34);
output(0, 192) <= input(2);
output(0, 193) <= input(3);
output(0, 194) <= input(4);
output(0, 195) <= input(5);
output(0, 196) <= input(6);
output(0, 197) <= input(7);
output(0, 198) <= input(8);
output(0, 199) <= input(9);
output(0, 200) <= input(10);
output(0, 201) <= input(11);
output(0, 202) <= input(12);
output(0, 203) <= input(13);
output(0, 204) <= input(14);
output(0, 205) <= input(15);
output(0, 206) <= input(32);
output(0, 207) <= input(34);
output(0, 208) <= input(18);
output(0, 209) <= input(19);
output(0, 210) <= input(20);
output(0, 211) <= input(21);
output(0, 212) <= input(22);
output(0, 213) <= input(23);
output(0, 214) <= input(24);
output(0, 215) <= input(25);
output(0, 216) <= input(26);
output(0, 217) <= input(27);
output(0, 218) <= input(28);
output(0, 219) <= input(29);
output(0, 220) <= input(30);
output(0, 221) <= input(31);
output(0, 222) <= input(33);
output(0, 223) <= input(35);
output(0, 224) <= input(18);
output(0, 225) <= input(19);
output(0, 226) <= input(20);
output(0, 227) <= input(21);
output(0, 228) <= input(22);
output(0, 229) <= input(23);
output(0, 230) <= input(24);
output(0, 231) <= input(25);
output(0, 232) <= input(26);
output(0, 233) <= input(27);
output(0, 234) <= input(28);
output(0, 235) <= input(29);
output(0, 236) <= input(30);
output(0, 237) <= input(31);
output(0, 238) <= input(33);
output(0, 239) <= input(35);
output(0, 240) <= input(3);
output(0, 241) <= input(4);
output(0, 242) <= input(5);
output(0, 243) <= input(6);
output(0, 244) <= input(7);
output(0, 245) <= input(8);
output(0, 246) <= input(9);
output(0, 247) <= input(10);
output(0, 248) <= input(11);
output(0, 249) <= input(12);
output(0, 250) <= input(13);
output(0, 251) <= input(14);
output(0, 252) <= input(15);
output(0, 253) <= input(32);
output(0, 254) <= input(34);
output(0, 255) <= input(36);
output(1, 0) <= input(1);
output(1, 1) <= input(2);
output(1, 2) <= input(3);
output(1, 3) <= input(4);
output(1, 4) <= input(5);
output(1, 5) <= input(6);
output(1, 6) <= input(7);
output(1, 7) <= input(8);
output(1, 8) <= input(9);
output(1, 9) <= input(10);
output(1, 10) <= input(11);
output(1, 11) <= input(12);
output(1, 12) <= input(13);
output(1, 13) <= input(14);
output(1, 14) <= input(15);
output(1, 15) <= input(32);
output(1, 16) <= input(17);
output(1, 17) <= input(18);
output(1, 18) <= input(19);
output(1, 19) <= input(20);
output(1, 20) <= input(21);
output(1, 21) <= input(22);
output(1, 22) <= input(23);
output(1, 23) <= input(24);
output(1, 24) <= input(25);
output(1, 25) <= input(26);
output(1, 26) <= input(27);
output(1, 27) <= input(28);
output(1, 28) <= input(29);
output(1, 29) <= input(30);
output(1, 30) <= input(31);
output(1, 31) <= input(33);
output(1, 32) <= input(17);
output(1, 33) <= input(18);
output(1, 34) <= input(19);
output(1, 35) <= input(20);
output(1, 36) <= input(21);
output(1, 37) <= input(22);
output(1, 38) <= input(23);
output(1, 39) <= input(24);
output(1, 40) <= input(25);
output(1, 41) <= input(26);
output(1, 42) <= input(27);
output(1, 43) <= input(28);
output(1, 44) <= input(29);
output(1, 45) <= input(30);
output(1, 46) <= input(31);
output(1, 47) <= input(33);
output(1, 48) <= input(2);
output(1, 49) <= input(3);
output(1, 50) <= input(4);
output(1, 51) <= input(5);
output(1, 52) <= input(6);
output(1, 53) <= input(7);
output(1, 54) <= input(8);
output(1, 55) <= input(9);
output(1, 56) <= input(10);
output(1, 57) <= input(11);
output(1, 58) <= input(12);
output(1, 59) <= input(13);
output(1, 60) <= input(14);
output(1, 61) <= input(15);
output(1, 62) <= input(32);
output(1, 63) <= input(34);
output(1, 64) <= input(2);
output(1, 65) <= input(3);
output(1, 66) <= input(4);
output(1, 67) <= input(5);
output(1, 68) <= input(6);
output(1, 69) <= input(7);
output(1, 70) <= input(8);
output(1, 71) <= input(9);
output(1, 72) <= input(10);
output(1, 73) <= input(11);
output(1, 74) <= input(12);
output(1, 75) <= input(13);
output(1, 76) <= input(14);
output(1, 77) <= input(15);
output(1, 78) <= input(32);
output(1, 79) <= input(34);
output(1, 80) <= input(18);
output(1, 81) <= input(19);
output(1, 82) <= input(20);
output(1, 83) <= input(21);
output(1, 84) <= input(22);
output(1, 85) <= input(23);
output(1, 86) <= input(24);
output(1, 87) <= input(25);
output(1, 88) <= input(26);
output(1, 89) <= input(27);
output(1, 90) <= input(28);
output(1, 91) <= input(29);
output(1, 92) <= input(30);
output(1, 93) <= input(31);
output(1, 94) <= input(33);
output(1, 95) <= input(35);
output(1, 96) <= input(18);
output(1, 97) <= input(19);
output(1, 98) <= input(20);
output(1, 99) <= input(21);
output(1, 100) <= input(22);
output(1, 101) <= input(23);
output(1, 102) <= input(24);
output(1, 103) <= input(25);
output(1, 104) <= input(26);
output(1, 105) <= input(27);
output(1, 106) <= input(28);
output(1, 107) <= input(29);
output(1, 108) <= input(30);
output(1, 109) <= input(31);
output(1, 110) <= input(33);
output(1, 111) <= input(35);
output(1, 112) <= input(3);
output(1, 113) <= input(4);
output(1, 114) <= input(5);
output(1, 115) <= input(6);
output(1, 116) <= input(7);
output(1, 117) <= input(8);
output(1, 118) <= input(9);
output(1, 119) <= input(10);
output(1, 120) <= input(11);
output(1, 121) <= input(12);
output(1, 122) <= input(13);
output(1, 123) <= input(14);
output(1, 124) <= input(15);
output(1, 125) <= input(32);
output(1, 126) <= input(34);
output(1, 127) <= input(36);
output(1, 128) <= input(3);
output(1, 129) <= input(4);
output(1, 130) <= input(5);
output(1, 131) <= input(6);
output(1, 132) <= input(7);
output(1, 133) <= input(8);
output(1, 134) <= input(9);
output(1, 135) <= input(10);
output(1, 136) <= input(11);
output(1, 137) <= input(12);
output(1, 138) <= input(13);
output(1, 139) <= input(14);
output(1, 140) <= input(15);
output(1, 141) <= input(32);
output(1, 142) <= input(34);
output(1, 143) <= input(36);
output(1, 144) <= input(19);
output(1, 145) <= input(20);
output(1, 146) <= input(21);
output(1, 147) <= input(22);
output(1, 148) <= input(23);
output(1, 149) <= input(24);
output(1, 150) <= input(25);
output(1, 151) <= input(26);
output(1, 152) <= input(27);
output(1, 153) <= input(28);
output(1, 154) <= input(29);
output(1, 155) <= input(30);
output(1, 156) <= input(31);
output(1, 157) <= input(33);
output(1, 158) <= input(35);
output(1, 159) <= input(37);
output(1, 160) <= input(19);
output(1, 161) <= input(20);
output(1, 162) <= input(21);
output(1, 163) <= input(22);
output(1, 164) <= input(23);
output(1, 165) <= input(24);
output(1, 166) <= input(25);
output(1, 167) <= input(26);
output(1, 168) <= input(27);
output(1, 169) <= input(28);
output(1, 170) <= input(29);
output(1, 171) <= input(30);
output(1, 172) <= input(31);
output(1, 173) <= input(33);
output(1, 174) <= input(35);
output(1, 175) <= input(37);
output(1, 176) <= input(4);
output(1, 177) <= input(5);
output(1, 178) <= input(6);
output(1, 179) <= input(7);
output(1, 180) <= input(8);
output(1, 181) <= input(9);
output(1, 182) <= input(10);
output(1, 183) <= input(11);
output(1, 184) <= input(12);
output(1, 185) <= input(13);
output(1, 186) <= input(14);
output(1, 187) <= input(15);
output(1, 188) <= input(32);
output(1, 189) <= input(34);
output(1, 190) <= input(36);
output(1, 191) <= input(38);
output(1, 192) <= input(4);
output(1, 193) <= input(5);
output(1, 194) <= input(6);
output(1, 195) <= input(7);
output(1, 196) <= input(8);
output(1, 197) <= input(9);
output(1, 198) <= input(10);
output(1, 199) <= input(11);
output(1, 200) <= input(12);
output(1, 201) <= input(13);
output(1, 202) <= input(14);
output(1, 203) <= input(15);
output(1, 204) <= input(32);
output(1, 205) <= input(34);
output(1, 206) <= input(36);
output(1, 207) <= input(38);
output(1, 208) <= input(20);
output(1, 209) <= input(21);
output(1, 210) <= input(22);
output(1, 211) <= input(23);
output(1, 212) <= input(24);
output(1, 213) <= input(25);
output(1, 214) <= input(26);
output(1, 215) <= input(27);
output(1, 216) <= input(28);
output(1, 217) <= input(29);
output(1, 218) <= input(30);
output(1, 219) <= input(31);
output(1, 220) <= input(33);
output(1, 221) <= input(35);
output(1, 222) <= input(37);
output(1, 223) <= input(39);
output(1, 224) <= input(20);
output(1, 225) <= input(21);
output(1, 226) <= input(22);
output(1, 227) <= input(23);
output(1, 228) <= input(24);
output(1, 229) <= input(25);
output(1, 230) <= input(26);
output(1, 231) <= input(27);
output(1, 232) <= input(28);
output(1, 233) <= input(29);
output(1, 234) <= input(30);
output(1, 235) <= input(31);
output(1, 236) <= input(33);
output(1, 237) <= input(35);
output(1, 238) <= input(37);
output(1, 239) <= input(39);
output(1, 240) <= input(5);
output(1, 241) <= input(6);
output(1, 242) <= input(7);
output(1, 243) <= input(8);
output(1, 244) <= input(9);
output(1, 245) <= input(10);
output(1, 246) <= input(11);
output(1, 247) <= input(12);
output(1, 248) <= input(13);
output(1, 249) <= input(14);
output(1, 250) <= input(15);
output(1, 251) <= input(32);
output(1, 252) <= input(34);
output(1, 253) <= input(36);
output(1, 254) <= input(38);
output(1, 255) <= input(40);
output(2, 0) <= input(2);
output(2, 1) <= input(3);
output(2, 2) <= input(4);
output(2, 3) <= input(5);
output(2, 4) <= input(6);
output(2, 5) <= input(7);
output(2, 6) <= input(8);
output(2, 7) <= input(9);
output(2, 8) <= input(10);
output(2, 9) <= input(11);
output(2, 10) <= input(12);
output(2, 11) <= input(13);
output(2, 12) <= input(14);
output(2, 13) <= input(15);
output(2, 14) <= input(32);
output(2, 15) <= input(34);
output(2, 16) <= input(18);
output(2, 17) <= input(19);
output(2, 18) <= input(20);
output(2, 19) <= input(21);
output(2, 20) <= input(22);
output(2, 21) <= input(23);
output(2, 22) <= input(24);
output(2, 23) <= input(25);
output(2, 24) <= input(26);
output(2, 25) <= input(27);
output(2, 26) <= input(28);
output(2, 27) <= input(29);
output(2, 28) <= input(30);
output(2, 29) <= input(31);
output(2, 30) <= input(33);
output(2, 31) <= input(35);
output(2, 32) <= input(18);
output(2, 33) <= input(19);
output(2, 34) <= input(20);
output(2, 35) <= input(21);
output(2, 36) <= input(22);
output(2, 37) <= input(23);
output(2, 38) <= input(24);
output(2, 39) <= input(25);
output(2, 40) <= input(26);
output(2, 41) <= input(27);
output(2, 42) <= input(28);
output(2, 43) <= input(29);
output(2, 44) <= input(30);
output(2, 45) <= input(31);
output(2, 46) <= input(33);
output(2, 47) <= input(35);
output(2, 48) <= input(3);
output(2, 49) <= input(4);
output(2, 50) <= input(5);
output(2, 51) <= input(6);
output(2, 52) <= input(7);
output(2, 53) <= input(8);
output(2, 54) <= input(9);
output(2, 55) <= input(10);
output(2, 56) <= input(11);
output(2, 57) <= input(12);
output(2, 58) <= input(13);
output(2, 59) <= input(14);
output(2, 60) <= input(15);
output(2, 61) <= input(32);
output(2, 62) <= input(34);
output(2, 63) <= input(36);
output(2, 64) <= input(19);
output(2, 65) <= input(20);
output(2, 66) <= input(21);
output(2, 67) <= input(22);
output(2, 68) <= input(23);
output(2, 69) <= input(24);
output(2, 70) <= input(25);
output(2, 71) <= input(26);
output(2, 72) <= input(27);
output(2, 73) <= input(28);
output(2, 74) <= input(29);
output(2, 75) <= input(30);
output(2, 76) <= input(31);
output(2, 77) <= input(33);
output(2, 78) <= input(35);
output(2, 79) <= input(37);
output(2, 80) <= input(19);
output(2, 81) <= input(20);
output(2, 82) <= input(21);
output(2, 83) <= input(22);
output(2, 84) <= input(23);
output(2, 85) <= input(24);
output(2, 86) <= input(25);
output(2, 87) <= input(26);
output(2, 88) <= input(27);
output(2, 89) <= input(28);
output(2, 90) <= input(29);
output(2, 91) <= input(30);
output(2, 92) <= input(31);
output(2, 93) <= input(33);
output(2, 94) <= input(35);
output(2, 95) <= input(37);
output(2, 96) <= input(4);
output(2, 97) <= input(5);
output(2, 98) <= input(6);
output(2, 99) <= input(7);
output(2, 100) <= input(8);
output(2, 101) <= input(9);
output(2, 102) <= input(10);
output(2, 103) <= input(11);
output(2, 104) <= input(12);
output(2, 105) <= input(13);
output(2, 106) <= input(14);
output(2, 107) <= input(15);
output(2, 108) <= input(32);
output(2, 109) <= input(34);
output(2, 110) <= input(36);
output(2, 111) <= input(38);
output(2, 112) <= input(20);
output(2, 113) <= input(21);
output(2, 114) <= input(22);
output(2, 115) <= input(23);
output(2, 116) <= input(24);
output(2, 117) <= input(25);
output(2, 118) <= input(26);
output(2, 119) <= input(27);
output(2, 120) <= input(28);
output(2, 121) <= input(29);
output(2, 122) <= input(30);
output(2, 123) <= input(31);
output(2, 124) <= input(33);
output(2, 125) <= input(35);
output(2, 126) <= input(37);
output(2, 127) <= input(39);
output(2, 128) <= input(20);
output(2, 129) <= input(21);
output(2, 130) <= input(22);
output(2, 131) <= input(23);
output(2, 132) <= input(24);
output(2, 133) <= input(25);
output(2, 134) <= input(26);
output(2, 135) <= input(27);
output(2, 136) <= input(28);
output(2, 137) <= input(29);
output(2, 138) <= input(30);
output(2, 139) <= input(31);
output(2, 140) <= input(33);
output(2, 141) <= input(35);
output(2, 142) <= input(37);
output(2, 143) <= input(39);
output(2, 144) <= input(5);
output(2, 145) <= input(6);
output(2, 146) <= input(7);
output(2, 147) <= input(8);
output(2, 148) <= input(9);
output(2, 149) <= input(10);
output(2, 150) <= input(11);
output(2, 151) <= input(12);
output(2, 152) <= input(13);
output(2, 153) <= input(14);
output(2, 154) <= input(15);
output(2, 155) <= input(32);
output(2, 156) <= input(34);
output(2, 157) <= input(36);
output(2, 158) <= input(38);
output(2, 159) <= input(40);
output(2, 160) <= input(5);
output(2, 161) <= input(6);
output(2, 162) <= input(7);
output(2, 163) <= input(8);
output(2, 164) <= input(9);
output(2, 165) <= input(10);
output(2, 166) <= input(11);
output(2, 167) <= input(12);
output(2, 168) <= input(13);
output(2, 169) <= input(14);
output(2, 170) <= input(15);
output(2, 171) <= input(32);
output(2, 172) <= input(34);
output(2, 173) <= input(36);
output(2, 174) <= input(38);
output(2, 175) <= input(40);
output(2, 176) <= input(21);
output(2, 177) <= input(22);
output(2, 178) <= input(23);
output(2, 179) <= input(24);
output(2, 180) <= input(25);
output(2, 181) <= input(26);
output(2, 182) <= input(27);
output(2, 183) <= input(28);
output(2, 184) <= input(29);
output(2, 185) <= input(30);
output(2, 186) <= input(31);
output(2, 187) <= input(33);
output(2, 188) <= input(35);
output(2, 189) <= input(37);
output(2, 190) <= input(39);
output(2, 191) <= input(41);
output(2, 192) <= input(6);
output(2, 193) <= input(7);
output(2, 194) <= input(8);
output(2, 195) <= input(9);
output(2, 196) <= input(10);
output(2, 197) <= input(11);
output(2, 198) <= input(12);
output(2, 199) <= input(13);
output(2, 200) <= input(14);
output(2, 201) <= input(15);
output(2, 202) <= input(32);
output(2, 203) <= input(34);
output(2, 204) <= input(36);
output(2, 205) <= input(38);
output(2, 206) <= input(40);
output(2, 207) <= input(42);
output(2, 208) <= input(6);
output(2, 209) <= input(7);
output(2, 210) <= input(8);
output(2, 211) <= input(9);
output(2, 212) <= input(10);
output(2, 213) <= input(11);
output(2, 214) <= input(12);
output(2, 215) <= input(13);
output(2, 216) <= input(14);
output(2, 217) <= input(15);
output(2, 218) <= input(32);
output(2, 219) <= input(34);
output(2, 220) <= input(36);
output(2, 221) <= input(38);
output(2, 222) <= input(40);
output(2, 223) <= input(42);
output(2, 224) <= input(22);
output(2, 225) <= input(23);
output(2, 226) <= input(24);
output(2, 227) <= input(25);
output(2, 228) <= input(26);
output(2, 229) <= input(27);
output(2, 230) <= input(28);
output(2, 231) <= input(29);
output(2, 232) <= input(30);
output(2, 233) <= input(31);
output(2, 234) <= input(33);
output(2, 235) <= input(35);
output(2, 236) <= input(37);
output(2, 237) <= input(39);
output(2, 238) <= input(41);
output(2, 239) <= input(43);
output(2, 240) <= input(7);
output(2, 241) <= input(8);
output(2, 242) <= input(9);
output(2, 243) <= input(10);
output(2, 244) <= input(11);
output(2, 245) <= input(12);
output(2, 246) <= input(13);
output(2, 247) <= input(14);
output(2, 248) <= input(15);
output(2, 249) <= input(32);
output(2, 250) <= input(34);
output(2, 251) <= input(36);
output(2, 252) <= input(38);
output(2, 253) <= input(40);
output(2, 254) <= input(42);
output(2, 255) <= input(44);
output(3, 0) <= input(3);
output(3, 1) <= input(4);
output(3, 2) <= input(5);
output(3, 3) <= input(6);
output(3, 4) <= input(7);
output(3, 5) <= input(8);
output(3, 6) <= input(9);
output(3, 7) <= input(10);
output(3, 8) <= input(11);
output(3, 9) <= input(12);
output(3, 10) <= input(13);
output(3, 11) <= input(14);
output(3, 12) <= input(15);
output(3, 13) <= input(32);
output(3, 14) <= input(34);
output(3, 15) <= input(36);
output(3, 16) <= input(19);
output(3, 17) <= input(20);
output(3, 18) <= input(21);
output(3, 19) <= input(22);
output(3, 20) <= input(23);
output(3, 21) <= input(24);
output(3, 22) <= input(25);
output(3, 23) <= input(26);
output(3, 24) <= input(27);
output(3, 25) <= input(28);
output(3, 26) <= input(29);
output(3, 27) <= input(30);
output(3, 28) <= input(31);
output(3, 29) <= input(33);
output(3, 30) <= input(35);
output(3, 31) <= input(37);
output(3, 32) <= input(4);
output(3, 33) <= input(5);
output(3, 34) <= input(6);
output(3, 35) <= input(7);
output(3, 36) <= input(8);
output(3, 37) <= input(9);
output(3, 38) <= input(10);
output(3, 39) <= input(11);
output(3, 40) <= input(12);
output(3, 41) <= input(13);
output(3, 42) <= input(14);
output(3, 43) <= input(15);
output(3, 44) <= input(32);
output(3, 45) <= input(34);
output(3, 46) <= input(36);
output(3, 47) <= input(38);
output(3, 48) <= input(20);
output(3, 49) <= input(21);
output(3, 50) <= input(22);
output(3, 51) <= input(23);
output(3, 52) <= input(24);
output(3, 53) <= input(25);
output(3, 54) <= input(26);
output(3, 55) <= input(27);
output(3, 56) <= input(28);
output(3, 57) <= input(29);
output(3, 58) <= input(30);
output(3, 59) <= input(31);
output(3, 60) <= input(33);
output(3, 61) <= input(35);
output(3, 62) <= input(37);
output(3, 63) <= input(39);
output(3, 64) <= input(20);
output(3, 65) <= input(21);
output(3, 66) <= input(22);
output(3, 67) <= input(23);
output(3, 68) <= input(24);
output(3, 69) <= input(25);
output(3, 70) <= input(26);
output(3, 71) <= input(27);
output(3, 72) <= input(28);
output(3, 73) <= input(29);
output(3, 74) <= input(30);
output(3, 75) <= input(31);
output(3, 76) <= input(33);
output(3, 77) <= input(35);
output(3, 78) <= input(37);
output(3, 79) <= input(39);
output(3, 80) <= input(5);
output(3, 81) <= input(6);
output(3, 82) <= input(7);
output(3, 83) <= input(8);
output(3, 84) <= input(9);
output(3, 85) <= input(10);
output(3, 86) <= input(11);
output(3, 87) <= input(12);
output(3, 88) <= input(13);
output(3, 89) <= input(14);
output(3, 90) <= input(15);
output(3, 91) <= input(32);
output(3, 92) <= input(34);
output(3, 93) <= input(36);
output(3, 94) <= input(38);
output(3, 95) <= input(40);
output(3, 96) <= input(21);
output(3, 97) <= input(22);
output(3, 98) <= input(23);
output(3, 99) <= input(24);
output(3, 100) <= input(25);
output(3, 101) <= input(26);
output(3, 102) <= input(27);
output(3, 103) <= input(28);
output(3, 104) <= input(29);
output(3, 105) <= input(30);
output(3, 106) <= input(31);
output(3, 107) <= input(33);
output(3, 108) <= input(35);
output(3, 109) <= input(37);
output(3, 110) <= input(39);
output(3, 111) <= input(41);
output(3, 112) <= input(6);
output(3, 113) <= input(7);
output(3, 114) <= input(8);
output(3, 115) <= input(9);
output(3, 116) <= input(10);
output(3, 117) <= input(11);
output(3, 118) <= input(12);
output(3, 119) <= input(13);
output(3, 120) <= input(14);
output(3, 121) <= input(15);
output(3, 122) <= input(32);
output(3, 123) <= input(34);
output(3, 124) <= input(36);
output(3, 125) <= input(38);
output(3, 126) <= input(40);
output(3, 127) <= input(42);
output(3, 128) <= input(6);
output(3, 129) <= input(7);
output(3, 130) <= input(8);
output(3, 131) <= input(9);
output(3, 132) <= input(10);
output(3, 133) <= input(11);
output(3, 134) <= input(12);
output(3, 135) <= input(13);
output(3, 136) <= input(14);
output(3, 137) <= input(15);
output(3, 138) <= input(32);
output(3, 139) <= input(34);
output(3, 140) <= input(36);
output(3, 141) <= input(38);
output(3, 142) <= input(40);
output(3, 143) <= input(42);
output(3, 144) <= input(22);
output(3, 145) <= input(23);
output(3, 146) <= input(24);
output(3, 147) <= input(25);
output(3, 148) <= input(26);
output(3, 149) <= input(27);
output(3, 150) <= input(28);
output(3, 151) <= input(29);
output(3, 152) <= input(30);
output(3, 153) <= input(31);
output(3, 154) <= input(33);
output(3, 155) <= input(35);
output(3, 156) <= input(37);
output(3, 157) <= input(39);
output(3, 158) <= input(41);
output(3, 159) <= input(43);
output(3, 160) <= input(7);
output(3, 161) <= input(8);
output(3, 162) <= input(9);
output(3, 163) <= input(10);
output(3, 164) <= input(11);
output(3, 165) <= input(12);
output(3, 166) <= input(13);
output(3, 167) <= input(14);
output(3, 168) <= input(15);
output(3, 169) <= input(32);
output(3, 170) <= input(34);
output(3, 171) <= input(36);
output(3, 172) <= input(38);
output(3, 173) <= input(40);
output(3, 174) <= input(42);
output(3, 175) <= input(44);
output(3, 176) <= input(23);
output(3, 177) <= input(24);
output(3, 178) <= input(25);
output(3, 179) <= input(26);
output(3, 180) <= input(27);
output(3, 181) <= input(28);
output(3, 182) <= input(29);
output(3, 183) <= input(30);
output(3, 184) <= input(31);
output(3, 185) <= input(33);
output(3, 186) <= input(35);
output(3, 187) <= input(37);
output(3, 188) <= input(39);
output(3, 189) <= input(41);
output(3, 190) <= input(43);
output(3, 191) <= input(45);
output(3, 192) <= input(23);
output(3, 193) <= input(24);
output(3, 194) <= input(25);
output(3, 195) <= input(26);
output(3, 196) <= input(27);
output(3, 197) <= input(28);
output(3, 198) <= input(29);
output(3, 199) <= input(30);
output(3, 200) <= input(31);
output(3, 201) <= input(33);
output(3, 202) <= input(35);
output(3, 203) <= input(37);
output(3, 204) <= input(39);
output(3, 205) <= input(41);
output(3, 206) <= input(43);
output(3, 207) <= input(45);
output(3, 208) <= input(8);
output(3, 209) <= input(9);
output(3, 210) <= input(10);
output(3, 211) <= input(11);
output(3, 212) <= input(12);
output(3, 213) <= input(13);
output(3, 214) <= input(14);
output(3, 215) <= input(15);
output(3, 216) <= input(32);
output(3, 217) <= input(34);
output(3, 218) <= input(36);
output(3, 219) <= input(38);
output(3, 220) <= input(40);
output(3, 221) <= input(42);
output(3, 222) <= input(44);
output(3, 223) <= input(46);
output(3, 224) <= input(24);
output(3, 225) <= input(25);
output(3, 226) <= input(26);
output(3, 227) <= input(27);
output(3, 228) <= input(28);
output(3, 229) <= input(29);
output(3, 230) <= input(30);
output(3, 231) <= input(31);
output(3, 232) <= input(33);
output(3, 233) <= input(35);
output(3, 234) <= input(37);
output(3, 235) <= input(39);
output(3, 236) <= input(41);
output(3, 237) <= input(43);
output(3, 238) <= input(45);
output(3, 239) <= input(47);
output(3, 240) <= input(9);
output(3, 241) <= input(10);
output(3, 242) <= input(11);
output(3, 243) <= input(12);
output(3, 244) <= input(13);
output(3, 245) <= input(14);
output(3, 246) <= input(15);
output(3, 247) <= input(32);
output(3, 248) <= input(34);
output(3, 249) <= input(36);
output(3, 250) <= input(38);
output(3, 251) <= input(40);
output(3, 252) <= input(42);
output(3, 253) <= input(44);
output(3, 254) <= input(46);
output(3, 255) <= input(48);
output(4, 0) <= input(4);
output(4, 1) <= input(5);
output(4, 2) <= input(6);
output(4, 3) <= input(7);
output(4, 4) <= input(8);
output(4, 5) <= input(9);
output(4, 6) <= input(10);
output(4, 7) <= input(11);
output(4, 8) <= input(12);
output(4, 9) <= input(13);
output(4, 10) <= input(14);
output(4, 11) <= input(15);
output(4, 12) <= input(32);
output(4, 13) <= input(34);
output(4, 14) <= input(36);
output(4, 15) <= input(38);
output(4, 16) <= input(20);
output(4, 17) <= input(21);
output(4, 18) <= input(22);
output(4, 19) <= input(23);
output(4, 20) <= input(24);
output(4, 21) <= input(25);
output(4, 22) <= input(26);
output(4, 23) <= input(27);
output(4, 24) <= input(28);
output(4, 25) <= input(29);
output(4, 26) <= input(30);
output(4, 27) <= input(31);
output(4, 28) <= input(33);
output(4, 29) <= input(35);
output(4, 30) <= input(37);
output(4, 31) <= input(39);
output(4, 32) <= input(5);
output(4, 33) <= input(6);
output(4, 34) <= input(7);
output(4, 35) <= input(8);
output(4, 36) <= input(9);
output(4, 37) <= input(10);
output(4, 38) <= input(11);
output(4, 39) <= input(12);
output(4, 40) <= input(13);
output(4, 41) <= input(14);
output(4, 42) <= input(15);
output(4, 43) <= input(32);
output(4, 44) <= input(34);
output(4, 45) <= input(36);
output(4, 46) <= input(38);
output(4, 47) <= input(40);
output(4, 48) <= input(21);
output(4, 49) <= input(22);
output(4, 50) <= input(23);
output(4, 51) <= input(24);
output(4, 52) <= input(25);
output(4, 53) <= input(26);
output(4, 54) <= input(27);
output(4, 55) <= input(28);
output(4, 56) <= input(29);
output(4, 57) <= input(30);
output(4, 58) <= input(31);
output(4, 59) <= input(33);
output(4, 60) <= input(35);
output(4, 61) <= input(37);
output(4, 62) <= input(39);
output(4, 63) <= input(41);
output(4, 64) <= input(6);
output(4, 65) <= input(7);
output(4, 66) <= input(8);
output(4, 67) <= input(9);
output(4, 68) <= input(10);
output(4, 69) <= input(11);
output(4, 70) <= input(12);
output(4, 71) <= input(13);
output(4, 72) <= input(14);
output(4, 73) <= input(15);
output(4, 74) <= input(32);
output(4, 75) <= input(34);
output(4, 76) <= input(36);
output(4, 77) <= input(38);
output(4, 78) <= input(40);
output(4, 79) <= input(42);
output(4, 80) <= input(22);
output(4, 81) <= input(23);
output(4, 82) <= input(24);
output(4, 83) <= input(25);
output(4, 84) <= input(26);
output(4, 85) <= input(27);
output(4, 86) <= input(28);
output(4, 87) <= input(29);
output(4, 88) <= input(30);
output(4, 89) <= input(31);
output(4, 90) <= input(33);
output(4, 91) <= input(35);
output(4, 92) <= input(37);
output(4, 93) <= input(39);
output(4, 94) <= input(41);
output(4, 95) <= input(43);
output(4, 96) <= input(7);
output(4, 97) <= input(8);
output(4, 98) <= input(9);
output(4, 99) <= input(10);
output(4, 100) <= input(11);
output(4, 101) <= input(12);
output(4, 102) <= input(13);
output(4, 103) <= input(14);
output(4, 104) <= input(15);
output(4, 105) <= input(32);
output(4, 106) <= input(34);
output(4, 107) <= input(36);
output(4, 108) <= input(38);
output(4, 109) <= input(40);
output(4, 110) <= input(42);
output(4, 111) <= input(44);
output(4, 112) <= input(23);
output(4, 113) <= input(24);
output(4, 114) <= input(25);
output(4, 115) <= input(26);
output(4, 116) <= input(27);
output(4, 117) <= input(28);
output(4, 118) <= input(29);
output(4, 119) <= input(30);
output(4, 120) <= input(31);
output(4, 121) <= input(33);
output(4, 122) <= input(35);
output(4, 123) <= input(37);
output(4, 124) <= input(39);
output(4, 125) <= input(41);
output(4, 126) <= input(43);
output(4, 127) <= input(45);
output(4, 128) <= input(23);
output(4, 129) <= input(24);
output(4, 130) <= input(25);
output(4, 131) <= input(26);
output(4, 132) <= input(27);
output(4, 133) <= input(28);
output(4, 134) <= input(29);
output(4, 135) <= input(30);
output(4, 136) <= input(31);
output(4, 137) <= input(33);
output(4, 138) <= input(35);
output(4, 139) <= input(37);
output(4, 140) <= input(39);
output(4, 141) <= input(41);
output(4, 142) <= input(43);
output(4, 143) <= input(45);
output(4, 144) <= input(8);
output(4, 145) <= input(9);
output(4, 146) <= input(10);
output(4, 147) <= input(11);
output(4, 148) <= input(12);
output(4, 149) <= input(13);
output(4, 150) <= input(14);
output(4, 151) <= input(15);
output(4, 152) <= input(32);
output(4, 153) <= input(34);
output(4, 154) <= input(36);
output(4, 155) <= input(38);
output(4, 156) <= input(40);
output(4, 157) <= input(42);
output(4, 158) <= input(44);
output(4, 159) <= input(46);
output(4, 160) <= input(24);
output(4, 161) <= input(25);
output(4, 162) <= input(26);
output(4, 163) <= input(27);
output(4, 164) <= input(28);
output(4, 165) <= input(29);
output(4, 166) <= input(30);
output(4, 167) <= input(31);
output(4, 168) <= input(33);
output(4, 169) <= input(35);
output(4, 170) <= input(37);
output(4, 171) <= input(39);
output(4, 172) <= input(41);
output(4, 173) <= input(43);
output(4, 174) <= input(45);
output(4, 175) <= input(47);
output(4, 176) <= input(9);
output(4, 177) <= input(10);
output(4, 178) <= input(11);
output(4, 179) <= input(12);
output(4, 180) <= input(13);
output(4, 181) <= input(14);
output(4, 182) <= input(15);
output(4, 183) <= input(32);
output(4, 184) <= input(34);
output(4, 185) <= input(36);
output(4, 186) <= input(38);
output(4, 187) <= input(40);
output(4, 188) <= input(42);
output(4, 189) <= input(44);
output(4, 190) <= input(46);
output(4, 191) <= input(48);
output(4, 192) <= input(25);
output(4, 193) <= input(26);
output(4, 194) <= input(27);
output(4, 195) <= input(28);
output(4, 196) <= input(29);
output(4, 197) <= input(30);
output(4, 198) <= input(31);
output(4, 199) <= input(33);
output(4, 200) <= input(35);
output(4, 201) <= input(37);
output(4, 202) <= input(39);
output(4, 203) <= input(41);
output(4, 204) <= input(43);
output(4, 205) <= input(45);
output(4, 206) <= input(47);
output(4, 207) <= input(49);
output(4, 208) <= input(10);
output(4, 209) <= input(11);
output(4, 210) <= input(12);
output(4, 211) <= input(13);
output(4, 212) <= input(14);
output(4, 213) <= input(15);
output(4, 214) <= input(32);
output(4, 215) <= input(34);
output(4, 216) <= input(36);
output(4, 217) <= input(38);
output(4, 218) <= input(40);
output(4, 219) <= input(42);
output(4, 220) <= input(44);
output(4, 221) <= input(46);
output(4, 222) <= input(48);
output(4, 223) <= input(50);
output(4, 224) <= input(26);
output(4, 225) <= input(27);
output(4, 226) <= input(28);
output(4, 227) <= input(29);
output(4, 228) <= input(30);
output(4, 229) <= input(31);
output(4, 230) <= input(33);
output(4, 231) <= input(35);
output(4, 232) <= input(37);
output(4, 233) <= input(39);
output(4, 234) <= input(41);
output(4, 235) <= input(43);
output(4, 236) <= input(45);
output(4, 237) <= input(47);
output(4, 238) <= input(49);
output(4, 239) <= input(51);
output(4, 240) <= input(11);
output(4, 241) <= input(12);
output(4, 242) <= input(13);
output(4, 243) <= input(14);
output(4, 244) <= input(15);
output(4, 245) <= input(32);
output(4, 246) <= input(34);
output(4, 247) <= input(36);
output(4, 248) <= input(38);
output(4, 249) <= input(40);
output(4, 250) <= input(42);
output(4, 251) <= input(44);
output(4, 252) <= input(46);
output(4, 253) <= input(48);
output(4, 254) <= input(50);
output(4, 255) <= input(52);
output(5, 0) <= input(21);
output(5, 1) <= input(22);
output(5, 2) <= input(23);
output(5, 3) <= input(24);
output(5, 4) <= input(25);
output(5, 5) <= input(26);
output(5, 6) <= input(27);
output(5, 7) <= input(28);
output(5, 8) <= input(29);
output(5, 9) <= input(30);
output(5, 10) <= input(31);
output(5, 11) <= input(33);
output(5, 12) <= input(35);
output(5, 13) <= input(37);
output(5, 14) <= input(39);
output(5, 15) <= input(41);
output(5, 16) <= input(6);
output(5, 17) <= input(7);
output(5, 18) <= input(8);
output(5, 19) <= input(9);
output(5, 20) <= input(10);
output(5, 21) <= input(11);
output(5, 22) <= input(12);
output(5, 23) <= input(13);
output(5, 24) <= input(14);
output(5, 25) <= input(15);
output(5, 26) <= input(32);
output(5, 27) <= input(34);
output(5, 28) <= input(36);
output(5, 29) <= input(38);
output(5, 30) <= input(40);
output(5, 31) <= input(42);
output(5, 32) <= input(22);
output(5, 33) <= input(23);
output(5, 34) <= input(24);
output(5, 35) <= input(25);
output(5, 36) <= input(26);
output(5, 37) <= input(27);
output(5, 38) <= input(28);
output(5, 39) <= input(29);
output(5, 40) <= input(30);
output(5, 41) <= input(31);
output(5, 42) <= input(33);
output(5, 43) <= input(35);
output(5, 44) <= input(37);
output(5, 45) <= input(39);
output(5, 46) <= input(41);
output(5, 47) <= input(43);
output(5, 48) <= input(7);
output(5, 49) <= input(8);
output(5, 50) <= input(9);
output(5, 51) <= input(10);
output(5, 52) <= input(11);
output(5, 53) <= input(12);
output(5, 54) <= input(13);
output(5, 55) <= input(14);
output(5, 56) <= input(15);
output(5, 57) <= input(32);
output(5, 58) <= input(34);
output(5, 59) <= input(36);
output(5, 60) <= input(38);
output(5, 61) <= input(40);
output(5, 62) <= input(42);
output(5, 63) <= input(44);
output(5, 64) <= input(23);
output(5, 65) <= input(24);
output(5, 66) <= input(25);
output(5, 67) <= input(26);
output(5, 68) <= input(27);
output(5, 69) <= input(28);
output(5, 70) <= input(29);
output(5, 71) <= input(30);
output(5, 72) <= input(31);
output(5, 73) <= input(33);
output(5, 74) <= input(35);
output(5, 75) <= input(37);
output(5, 76) <= input(39);
output(5, 77) <= input(41);
output(5, 78) <= input(43);
output(5, 79) <= input(45);
output(5, 80) <= input(8);
output(5, 81) <= input(9);
output(5, 82) <= input(10);
output(5, 83) <= input(11);
output(5, 84) <= input(12);
output(5, 85) <= input(13);
output(5, 86) <= input(14);
output(5, 87) <= input(15);
output(5, 88) <= input(32);
output(5, 89) <= input(34);
output(5, 90) <= input(36);
output(5, 91) <= input(38);
output(5, 92) <= input(40);
output(5, 93) <= input(42);
output(5, 94) <= input(44);
output(5, 95) <= input(46);
output(5, 96) <= input(24);
output(5, 97) <= input(25);
output(5, 98) <= input(26);
output(5, 99) <= input(27);
output(5, 100) <= input(28);
output(5, 101) <= input(29);
output(5, 102) <= input(30);
output(5, 103) <= input(31);
output(5, 104) <= input(33);
output(5, 105) <= input(35);
output(5, 106) <= input(37);
output(5, 107) <= input(39);
output(5, 108) <= input(41);
output(5, 109) <= input(43);
output(5, 110) <= input(45);
output(5, 111) <= input(47);
output(5, 112) <= input(9);
output(5, 113) <= input(10);
output(5, 114) <= input(11);
output(5, 115) <= input(12);
output(5, 116) <= input(13);
output(5, 117) <= input(14);
output(5, 118) <= input(15);
output(5, 119) <= input(32);
output(5, 120) <= input(34);
output(5, 121) <= input(36);
output(5, 122) <= input(38);
output(5, 123) <= input(40);
output(5, 124) <= input(42);
output(5, 125) <= input(44);
output(5, 126) <= input(46);
output(5, 127) <= input(48);
output(5, 128) <= input(25);
output(5, 129) <= input(26);
output(5, 130) <= input(27);
output(5, 131) <= input(28);
output(5, 132) <= input(29);
output(5, 133) <= input(30);
output(5, 134) <= input(31);
output(5, 135) <= input(33);
output(5, 136) <= input(35);
output(5, 137) <= input(37);
output(5, 138) <= input(39);
output(5, 139) <= input(41);
output(5, 140) <= input(43);
output(5, 141) <= input(45);
output(5, 142) <= input(47);
output(5, 143) <= input(49);
output(5, 144) <= input(10);
output(5, 145) <= input(11);
output(5, 146) <= input(12);
output(5, 147) <= input(13);
output(5, 148) <= input(14);
output(5, 149) <= input(15);
output(5, 150) <= input(32);
output(5, 151) <= input(34);
output(5, 152) <= input(36);
output(5, 153) <= input(38);
output(5, 154) <= input(40);
output(5, 155) <= input(42);
output(5, 156) <= input(44);
output(5, 157) <= input(46);
output(5, 158) <= input(48);
output(5, 159) <= input(50);
output(5, 160) <= input(26);
output(5, 161) <= input(27);
output(5, 162) <= input(28);
output(5, 163) <= input(29);
output(5, 164) <= input(30);
output(5, 165) <= input(31);
output(5, 166) <= input(33);
output(5, 167) <= input(35);
output(5, 168) <= input(37);
output(5, 169) <= input(39);
output(5, 170) <= input(41);
output(5, 171) <= input(43);
output(5, 172) <= input(45);
output(5, 173) <= input(47);
output(5, 174) <= input(49);
output(5, 175) <= input(51);
output(5, 176) <= input(11);
output(5, 177) <= input(12);
output(5, 178) <= input(13);
output(5, 179) <= input(14);
output(5, 180) <= input(15);
output(5, 181) <= input(32);
output(5, 182) <= input(34);
output(5, 183) <= input(36);
output(5, 184) <= input(38);
output(5, 185) <= input(40);
output(5, 186) <= input(42);
output(5, 187) <= input(44);
output(5, 188) <= input(46);
output(5, 189) <= input(48);
output(5, 190) <= input(50);
output(5, 191) <= input(52);
output(5, 192) <= input(27);
output(5, 193) <= input(28);
output(5, 194) <= input(29);
output(5, 195) <= input(30);
output(5, 196) <= input(31);
output(5, 197) <= input(33);
output(5, 198) <= input(35);
output(5, 199) <= input(37);
output(5, 200) <= input(39);
output(5, 201) <= input(41);
output(5, 202) <= input(43);
output(5, 203) <= input(45);
output(5, 204) <= input(47);
output(5, 205) <= input(49);
output(5, 206) <= input(51);
output(5, 207) <= input(53);
output(5, 208) <= input(12);
output(5, 209) <= input(13);
output(5, 210) <= input(14);
output(5, 211) <= input(15);
output(5, 212) <= input(32);
output(5, 213) <= input(34);
output(5, 214) <= input(36);
output(5, 215) <= input(38);
output(5, 216) <= input(40);
output(5, 217) <= input(42);
output(5, 218) <= input(44);
output(5, 219) <= input(46);
output(5, 220) <= input(48);
output(5, 221) <= input(50);
output(5, 222) <= input(52);
output(5, 223) <= input(54);
output(5, 224) <= input(28);
output(5, 225) <= input(29);
output(5, 226) <= input(30);
output(5, 227) <= input(31);
output(5, 228) <= input(33);
output(5, 229) <= input(35);
output(5, 230) <= input(37);
output(5, 231) <= input(39);
output(5, 232) <= input(41);
output(5, 233) <= input(43);
output(5, 234) <= input(45);
output(5, 235) <= input(47);
output(5, 236) <= input(49);
output(5, 237) <= input(51);
output(5, 238) <= input(53);
output(5, 239) <= input(55);
output(5, 240) <= input(13);
output(5, 241) <= input(14);
output(5, 242) <= input(15);
output(5, 243) <= input(32);
output(5, 244) <= input(34);
output(5, 245) <= input(36);
output(5, 246) <= input(38);
output(5, 247) <= input(40);
output(5, 248) <= input(42);
output(5, 249) <= input(44);
output(5, 250) <= input(46);
output(5, 251) <= input(48);
output(5, 252) <= input(50);
output(5, 253) <= input(52);
output(5, 254) <= input(54);
output(5, 255) <= input(56);
when "1111" =>
output(0, 0) <= input(0);
output(0, 1) <= input(1);
output(0, 2) <= input(2);
output(0, 3) <= input(3);
output(0, 4) <= input(4);
output(0, 5) <= input(5);
output(0, 6) <= input(6);
output(0, 7) <= input(7);
output(0, 8) <= input(8);
output(0, 9) <= input(9);
output(0, 10) <= input(10);
output(0, 11) <= input(11);
output(0, 12) <= input(12);
output(0, 13) <= input(13);
output(0, 14) <= input(14);
output(0, 15) <= input(15);
output(0, 16) <= input(16);
output(0, 17) <= input(17);
output(0, 18) <= input(18);
output(0, 19) <= input(19);
output(0, 20) <= input(20);
output(0, 21) <= input(21);
output(0, 22) <= input(22);
output(0, 23) <= input(23);
output(0, 24) <= input(24);
output(0, 25) <= input(25);
output(0, 26) <= input(26);
output(0, 27) <= input(27);
output(0, 28) <= input(28);
output(0, 29) <= input(29);
output(0, 30) <= input(30);
output(0, 31) <= input(31);
output(0, 32) <= input(1);
output(0, 33) <= input(2);
output(0, 34) <= input(3);
output(0, 35) <= input(4);
output(0, 36) <= input(5);
output(0, 37) <= input(6);
output(0, 38) <= input(7);
output(0, 39) <= input(8);
output(0, 40) <= input(9);
output(0, 41) <= input(10);
output(0, 42) <= input(11);
output(0, 43) <= input(12);
output(0, 44) <= input(13);
output(0, 45) <= input(14);
output(0, 46) <= input(15);
output(0, 47) <= input(32);
output(0, 48) <= input(17);
output(0, 49) <= input(18);
output(0, 50) <= input(19);
output(0, 51) <= input(20);
output(0, 52) <= input(21);
output(0, 53) <= input(22);
output(0, 54) <= input(23);
output(0, 55) <= input(24);
output(0, 56) <= input(25);
output(0, 57) <= input(26);
output(0, 58) <= input(27);
output(0, 59) <= input(28);
output(0, 60) <= input(29);
output(0, 61) <= input(30);
output(0, 62) <= input(31);
output(0, 63) <= input(33);
output(0, 64) <= input(2);
output(0, 65) <= input(3);
output(0, 66) <= input(4);
output(0, 67) <= input(5);
output(0, 68) <= input(6);
output(0, 69) <= input(7);
output(0, 70) <= input(8);
output(0, 71) <= input(9);
output(0, 72) <= input(10);
output(0, 73) <= input(11);
output(0, 74) <= input(12);
output(0, 75) <= input(13);
output(0, 76) <= input(14);
output(0, 77) <= input(15);
output(0, 78) <= input(32);
output(0, 79) <= input(34);
output(0, 80) <= input(18);
output(0, 81) <= input(19);
output(0, 82) <= input(20);
output(0, 83) <= input(21);
output(0, 84) <= input(22);
output(0, 85) <= input(23);
output(0, 86) <= input(24);
output(0, 87) <= input(25);
output(0, 88) <= input(26);
output(0, 89) <= input(27);
output(0, 90) <= input(28);
output(0, 91) <= input(29);
output(0, 92) <= input(30);
output(0, 93) <= input(31);
output(0, 94) <= input(33);
output(0, 95) <= input(35);
output(0, 96) <= input(3);
output(0, 97) <= input(4);
output(0, 98) <= input(5);
output(0, 99) <= input(6);
output(0, 100) <= input(7);
output(0, 101) <= input(8);
output(0, 102) <= input(9);
output(0, 103) <= input(10);
output(0, 104) <= input(11);
output(0, 105) <= input(12);
output(0, 106) <= input(13);
output(0, 107) <= input(14);
output(0, 108) <= input(15);
output(0, 109) <= input(32);
output(0, 110) <= input(34);
output(0, 111) <= input(36);
output(0, 112) <= input(4);
output(0, 113) <= input(5);
output(0, 114) <= input(6);
output(0, 115) <= input(7);
output(0, 116) <= input(8);
output(0, 117) <= input(9);
output(0, 118) <= input(10);
output(0, 119) <= input(11);
output(0, 120) <= input(12);
output(0, 121) <= input(13);
output(0, 122) <= input(14);
output(0, 123) <= input(15);
output(0, 124) <= input(32);
output(0, 125) <= input(34);
output(0, 126) <= input(36);
output(0, 127) <= input(37);
output(0, 128) <= input(20);
output(0, 129) <= input(21);
output(0, 130) <= input(22);
output(0, 131) <= input(23);
output(0, 132) <= input(24);
output(0, 133) <= input(25);
output(0, 134) <= input(26);
output(0, 135) <= input(27);
output(0, 136) <= input(28);
output(0, 137) <= input(29);
output(0, 138) <= input(30);
output(0, 139) <= input(31);
output(0, 140) <= input(33);
output(0, 141) <= input(35);
output(0, 142) <= input(38);
output(0, 143) <= input(39);
output(0, 144) <= input(5);
output(0, 145) <= input(6);
output(0, 146) <= input(7);
output(0, 147) <= input(8);
output(0, 148) <= input(9);
output(0, 149) <= input(10);
output(0, 150) <= input(11);
output(0, 151) <= input(12);
output(0, 152) <= input(13);
output(0, 153) <= input(14);
output(0, 154) <= input(15);
output(0, 155) <= input(32);
output(0, 156) <= input(34);
output(0, 157) <= input(36);
output(0, 158) <= input(37);
output(0, 159) <= input(40);
output(0, 160) <= input(21);
output(0, 161) <= input(22);
output(0, 162) <= input(23);
output(0, 163) <= input(24);
output(0, 164) <= input(25);
output(0, 165) <= input(26);
output(0, 166) <= input(27);
output(0, 167) <= input(28);
output(0, 168) <= input(29);
output(0, 169) <= input(30);
output(0, 170) <= input(31);
output(0, 171) <= input(33);
output(0, 172) <= input(35);
output(0, 173) <= input(38);
output(0, 174) <= input(39);
output(0, 175) <= input(41);
output(0, 176) <= input(6);
output(0, 177) <= input(7);
output(0, 178) <= input(8);
output(0, 179) <= input(9);
output(0, 180) <= input(10);
output(0, 181) <= input(11);
output(0, 182) <= input(12);
output(0, 183) <= input(13);
output(0, 184) <= input(14);
output(0, 185) <= input(15);
output(0, 186) <= input(32);
output(0, 187) <= input(34);
output(0, 188) <= input(36);
output(0, 189) <= input(37);
output(0, 190) <= input(40);
output(0, 191) <= input(42);
output(0, 192) <= input(22);
output(0, 193) <= input(23);
output(0, 194) <= input(24);
output(0, 195) <= input(25);
output(0, 196) <= input(26);
output(0, 197) <= input(27);
output(0, 198) <= input(28);
output(0, 199) <= input(29);
output(0, 200) <= input(30);
output(0, 201) <= input(31);
output(0, 202) <= input(33);
output(0, 203) <= input(35);
output(0, 204) <= input(38);
output(0, 205) <= input(39);
output(0, 206) <= input(41);
output(0, 207) <= input(43);
output(0, 208) <= input(7);
output(0, 209) <= input(8);
output(0, 210) <= input(9);
output(0, 211) <= input(10);
output(0, 212) <= input(11);
output(0, 213) <= input(12);
output(0, 214) <= input(13);
output(0, 215) <= input(14);
output(0, 216) <= input(15);
output(0, 217) <= input(32);
output(0, 218) <= input(34);
output(0, 219) <= input(36);
output(0, 220) <= input(37);
output(0, 221) <= input(40);
output(0, 222) <= input(42);
output(0, 223) <= input(44);
output(0, 224) <= input(23);
output(0, 225) <= input(24);
output(0, 226) <= input(25);
output(0, 227) <= input(26);
output(0, 228) <= input(27);
output(0, 229) <= input(28);
output(0, 230) <= input(29);
output(0, 231) <= input(30);
output(0, 232) <= input(31);
output(0, 233) <= input(33);
output(0, 234) <= input(35);
output(0, 235) <= input(38);
output(0, 236) <= input(39);
output(0, 237) <= input(41);
output(0, 238) <= input(43);
output(0, 239) <= input(45);
output(0, 240) <= input(24);
output(0, 241) <= input(25);
output(0, 242) <= input(26);
output(0, 243) <= input(27);
output(0, 244) <= input(28);
output(0, 245) <= input(29);
output(0, 246) <= input(30);
output(0, 247) <= input(31);
output(0, 248) <= input(33);
output(0, 249) <= input(35);
output(0, 250) <= input(38);
output(0, 251) <= input(39);
output(0, 252) <= input(41);
output(0, 253) <= input(43);
output(0, 254) <= input(45);
output(0, 255) <= input(46);
output(1, 0) <= input(1);
output(1, 1) <= input(2);
output(1, 2) <= input(3);
output(1, 3) <= input(4);
output(1, 4) <= input(5);
output(1, 5) <= input(6);
output(1, 6) <= input(7);
output(1, 7) <= input(8);
output(1, 8) <= input(9);
output(1, 9) <= input(10);
output(1, 10) <= input(11);
output(1, 11) <= input(12);
output(1, 12) <= input(13);
output(1, 13) <= input(14);
output(1, 14) <= input(15);
output(1, 15) <= input(32);
output(1, 16) <= input(17);
output(1, 17) <= input(18);
output(1, 18) <= input(19);
output(1, 19) <= input(20);
output(1, 20) <= input(21);
output(1, 21) <= input(22);
output(1, 22) <= input(23);
output(1, 23) <= input(24);
output(1, 24) <= input(25);
output(1, 25) <= input(26);
output(1, 26) <= input(27);
output(1, 27) <= input(28);
output(1, 28) <= input(29);
output(1, 29) <= input(30);
output(1, 30) <= input(31);
output(1, 31) <= input(33);
output(1, 32) <= input(2);
output(1, 33) <= input(3);
output(1, 34) <= input(4);
output(1, 35) <= input(5);
output(1, 36) <= input(6);
output(1, 37) <= input(7);
output(1, 38) <= input(8);
output(1, 39) <= input(9);
output(1, 40) <= input(10);
output(1, 41) <= input(11);
output(1, 42) <= input(12);
output(1, 43) <= input(13);
output(1, 44) <= input(14);
output(1, 45) <= input(15);
output(1, 46) <= input(32);
output(1, 47) <= input(34);
output(1, 48) <= input(3);
output(1, 49) <= input(4);
output(1, 50) <= input(5);
output(1, 51) <= input(6);
output(1, 52) <= input(7);
output(1, 53) <= input(8);
output(1, 54) <= input(9);
output(1, 55) <= input(10);
output(1, 56) <= input(11);
output(1, 57) <= input(12);
output(1, 58) <= input(13);
output(1, 59) <= input(14);
output(1, 60) <= input(15);
output(1, 61) <= input(32);
output(1, 62) <= input(34);
output(1, 63) <= input(36);
output(1, 64) <= input(19);
output(1, 65) <= input(20);
output(1, 66) <= input(21);
output(1, 67) <= input(22);
output(1, 68) <= input(23);
output(1, 69) <= input(24);
output(1, 70) <= input(25);
output(1, 71) <= input(26);
output(1, 72) <= input(27);
output(1, 73) <= input(28);
output(1, 74) <= input(29);
output(1, 75) <= input(30);
output(1, 76) <= input(31);
output(1, 77) <= input(33);
output(1, 78) <= input(35);
output(1, 79) <= input(38);
output(1, 80) <= input(4);
output(1, 81) <= input(5);
output(1, 82) <= input(6);
output(1, 83) <= input(7);
output(1, 84) <= input(8);
output(1, 85) <= input(9);
output(1, 86) <= input(10);
output(1, 87) <= input(11);
output(1, 88) <= input(12);
output(1, 89) <= input(13);
output(1, 90) <= input(14);
output(1, 91) <= input(15);
output(1, 92) <= input(32);
output(1, 93) <= input(34);
output(1, 94) <= input(36);
output(1, 95) <= input(37);
output(1, 96) <= input(20);
output(1, 97) <= input(21);
output(1, 98) <= input(22);
output(1, 99) <= input(23);
output(1, 100) <= input(24);
output(1, 101) <= input(25);
output(1, 102) <= input(26);
output(1, 103) <= input(27);
output(1, 104) <= input(28);
output(1, 105) <= input(29);
output(1, 106) <= input(30);
output(1, 107) <= input(31);
output(1, 108) <= input(33);
output(1, 109) <= input(35);
output(1, 110) <= input(38);
output(1, 111) <= input(39);
output(1, 112) <= input(21);
output(1, 113) <= input(22);
output(1, 114) <= input(23);
output(1, 115) <= input(24);
output(1, 116) <= input(25);
output(1, 117) <= input(26);
output(1, 118) <= input(27);
output(1, 119) <= input(28);
output(1, 120) <= input(29);
output(1, 121) <= input(30);
output(1, 122) <= input(31);
output(1, 123) <= input(33);
output(1, 124) <= input(35);
output(1, 125) <= input(38);
output(1, 126) <= input(39);
output(1, 127) <= input(41);
output(1, 128) <= input(6);
output(1, 129) <= input(7);
output(1, 130) <= input(8);
output(1, 131) <= input(9);
output(1, 132) <= input(10);
output(1, 133) <= input(11);
output(1, 134) <= input(12);
output(1, 135) <= input(13);
output(1, 136) <= input(14);
output(1, 137) <= input(15);
output(1, 138) <= input(32);
output(1, 139) <= input(34);
output(1, 140) <= input(36);
output(1, 141) <= input(37);
output(1, 142) <= input(40);
output(1, 143) <= input(42);
output(1, 144) <= input(22);
output(1, 145) <= input(23);
output(1, 146) <= input(24);
output(1, 147) <= input(25);
output(1, 148) <= input(26);
output(1, 149) <= input(27);
output(1, 150) <= input(28);
output(1, 151) <= input(29);
output(1, 152) <= input(30);
output(1, 153) <= input(31);
output(1, 154) <= input(33);
output(1, 155) <= input(35);
output(1, 156) <= input(38);
output(1, 157) <= input(39);
output(1, 158) <= input(41);
output(1, 159) <= input(43);
output(1, 160) <= input(7);
output(1, 161) <= input(8);
output(1, 162) <= input(9);
output(1, 163) <= input(10);
output(1, 164) <= input(11);
output(1, 165) <= input(12);
output(1, 166) <= input(13);
output(1, 167) <= input(14);
output(1, 168) <= input(15);
output(1, 169) <= input(32);
output(1, 170) <= input(34);
output(1, 171) <= input(36);
output(1, 172) <= input(37);
output(1, 173) <= input(40);
output(1, 174) <= input(42);
output(1, 175) <= input(44);
output(1, 176) <= input(8);
output(1, 177) <= input(9);
output(1, 178) <= input(10);
output(1, 179) <= input(11);
output(1, 180) <= input(12);
output(1, 181) <= input(13);
output(1, 182) <= input(14);
output(1, 183) <= input(15);
output(1, 184) <= input(32);
output(1, 185) <= input(34);
output(1, 186) <= input(36);
output(1, 187) <= input(37);
output(1, 188) <= input(40);
output(1, 189) <= input(42);
output(1, 190) <= input(44);
output(1, 191) <= input(47);
output(1, 192) <= input(24);
output(1, 193) <= input(25);
output(1, 194) <= input(26);
output(1, 195) <= input(27);
output(1, 196) <= input(28);
output(1, 197) <= input(29);
output(1, 198) <= input(30);
output(1, 199) <= input(31);
output(1, 200) <= input(33);
output(1, 201) <= input(35);
output(1, 202) <= input(38);
output(1, 203) <= input(39);
output(1, 204) <= input(41);
output(1, 205) <= input(43);
output(1, 206) <= input(45);
output(1, 207) <= input(46);
output(1, 208) <= input(9);
output(1, 209) <= input(10);
output(1, 210) <= input(11);
output(1, 211) <= input(12);
output(1, 212) <= input(13);
output(1, 213) <= input(14);
output(1, 214) <= input(15);
output(1, 215) <= input(32);
output(1, 216) <= input(34);
output(1, 217) <= input(36);
output(1, 218) <= input(37);
output(1, 219) <= input(40);
output(1, 220) <= input(42);
output(1, 221) <= input(44);
output(1, 222) <= input(47);
output(1, 223) <= input(48);
output(1, 224) <= input(25);
output(1, 225) <= input(26);
output(1, 226) <= input(27);
output(1, 227) <= input(28);
output(1, 228) <= input(29);
output(1, 229) <= input(30);
output(1, 230) <= input(31);
output(1, 231) <= input(33);
output(1, 232) <= input(35);
output(1, 233) <= input(38);
output(1, 234) <= input(39);
output(1, 235) <= input(41);
output(1, 236) <= input(43);
output(1, 237) <= input(45);
output(1, 238) <= input(46);
output(1, 239) <= input(49);
output(1, 240) <= input(26);
output(1, 241) <= input(27);
output(1, 242) <= input(28);
output(1, 243) <= input(29);
output(1, 244) <= input(30);
output(1, 245) <= input(31);
output(1, 246) <= input(33);
output(1, 247) <= input(35);
output(1, 248) <= input(38);
output(1, 249) <= input(39);
output(1, 250) <= input(41);
output(1, 251) <= input(43);
output(1, 252) <= input(45);
output(1, 253) <= input(46);
output(1, 254) <= input(49);
output(1, 255) <= input(50);
output(2, 0) <= input(18);
output(2, 1) <= input(19);
output(2, 2) <= input(20);
output(2, 3) <= input(21);
output(2, 4) <= input(22);
output(2, 5) <= input(23);
output(2, 6) <= input(24);
output(2, 7) <= input(25);
output(2, 8) <= input(26);
output(2, 9) <= input(27);
output(2, 10) <= input(28);
output(2, 11) <= input(29);
output(2, 12) <= input(30);
output(2, 13) <= input(31);
output(2, 14) <= input(33);
output(2, 15) <= input(35);
output(2, 16) <= input(3);
output(2, 17) <= input(4);
output(2, 18) <= input(5);
output(2, 19) <= input(6);
output(2, 20) <= input(7);
output(2, 21) <= input(8);
output(2, 22) <= input(9);
output(2, 23) <= input(10);
output(2, 24) <= input(11);
output(2, 25) <= input(12);
output(2, 26) <= input(13);
output(2, 27) <= input(14);
output(2, 28) <= input(15);
output(2, 29) <= input(32);
output(2, 30) <= input(34);
output(2, 31) <= input(36);
output(2, 32) <= input(4);
output(2, 33) <= input(5);
output(2, 34) <= input(6);
output(2, 35) <= input(7);
output(2, 36) <= input(8);
output(2, 37) <= input(9);
output(2, 38) <= input(10);
output(2, 39) <= input(11);
output(2, 40) <= input(12);
output(2, 41) <= input(13);
output(2, 42) <= input(14);
output(2, 43) <= input(15);
output(2, 44) <= input(32);
output(2, 45) <= input(34);
output(2, 46) <= input(36);
output(2, 47) <= input(37);
output(2, 48) <= input(20);
output(2, 49) <= input(21);
output(2, 50) <= input(22);
output(2, 51) <= input(23);
output(2, 52) <= input(24);
output(2, 53) <= input(25);
output(2, 54) <= input(26);
output(2, 55) <= input(27);
output(2, 56) <= input(28);
output(2, 57) <= input(29);
output(2, 58) <= input(30);
output(2, 59) <= input(31);
output(2, 60) <= input(33);
output(2, 61) <= input(35);
output(2, 62) <= input(38);
output(2, 63) <= input(39);
output(2, 64) <= input(21);
output(2, 65) <= input(22);
output(2, 66) <= input(23);
output(2, 67) <= input(24);
output(2, 68) <= input(25);
output(2, 69) <= input(26);
output(2, 70) <= input(27);
output(2, 71) <= input(28);
output(2, 72) <= input(29);
output(2, 73) <= input(30);
output(2, 74) <= input(31);
output(2, 75) <= input(33);
output(2, 76) <= input(35);
output(2, 77) <= input(38);
output(2, 78) <= input(39);
output(2, 79) <= input(41);
output(2, 80) <= input(6);
output(2, 81) <= input(7);
output(2, 82) <= input(8);
output(2, 83) <= input(9);
output(2, 84) <= input(10);
output(2, 85) <= input(11);
output(2, 86) <= input(12);
output(2, 87) <= input(13);
output(2, 88) <= input(14);
output(2, 89) <= input(15);
output(2, 90) <= input(32);
output(2, 91) <= input(34);
output(2, 92) <= input(36);
output(2, 93) <= input(37);
output(2, 94) <= input(40);
output(2, 95) <= input(42);
output(2, 96) <= input(7);
output(2, 97) <= input(8);
output(2, 98) <= input(9);
output(2, 99) <= input(10);
output(2, 100) <= input(11);
output(2, 101) <= input(12);
output(2, 102) <= input(13);
output(2, 103) <= input(14);
output(2, 104) <= input(15);
output(2, 105) <= input(32);
output(2, 106) <= input(34);
output(2, 107) <= input(36);
output(2, 108) <= input(37);
output(2, 109) <= input(40);
output(2, 110) <= input(42);
output(2, 111) <= input(44);
output(2, 112) <= input(23);
output(2, 113) <= input(24);
output(2, 114) <= input(25);
output(2, 115) <= input(26);
output(2, 116) <= input(27);
output(2, 117) <= input(28);
output(2, 118) <= input(29);
output(2, 119) <= input(30);
output(2, 120) <= input(31);
output(2, 121) <= input(33);
output(2, 122) <= input(35);
output(2, 123) <= input(38);
output(2, 124) <= input(39);
output(2, 125) <= input(41);
output(2, 126) <= input(43);
output(2, 127) <= input(45);
output(2, 128) <= input(8);
output(2, 129) <= input(9);
output(2, 130) <= input(10);
output(2, 131) <= input(11);
output(2, 132) <= input(12);
output(2, 133) <= input(13);
output(2, 134) <= input(14);
output(2, 135) <= input(15);
output(2, 136) <= input(32);
output(2, 137) <= input(34);
output(2, 138) <= input(36);
output(2, 139) <= input(37);
output(2, 140) <= input(40);
output(2, 141) <= input(42);
output(2, 142) <= input(44);
output(2, 143) <= input(47);
output(2, 144) <= input(9);
output(2, 145) <= input(10);
output(2, 146) <= input(11);
output(2, 147) <= input(12);
output(2, 148) <= input(13);
output(2, 149) <= input(14);
output(2, 150) <= input(15);
output(2, 151) <= input(32);
output(2, 152) <= input(34);
output(2, 153) <= input(36);
output(2, 154) <= input(37);
output(2, 155) <= input(40);
output(2, 156) <= input(42);
output(2, 157) <= input(44);
output(2, 158) <= input(47);
output(2, 159) <= input(48);
output(2, 160) <= input(25);
output(2, 161) <= input(26);
output(2, 162) <= input(27);
output(2, 163) <= input(28);
output(2, 164) <= input(29);
output(2, 165) <= input(30);
output(2, 166) <= input(31);
output(2, 167) <= input(33);
output(2, 168) <= input(35);
output(2, 169) <= input(38);
output(2, 170) <= input(39);
output(2, 171) <= input(41);
output(2, 172) <= input(43);
output(2, 173) <= input(45);
output(2, 174) <= input(46);
output(2, 175) <= input(49);
output(2, 176) <= input(26);
output(2, 177) <= input(27);
output(2, 178) <= input(28);
output(2, 179) <= input(29);
output(2, 180) <= input(30);
output(2, 181) <= input(31);
output(2, 182) <= input(33);
output(2, 183) <= input(35);
output(2, 184) <= input(38);
output(2, 185) <= input(39);
output(2, 186) <= input(41);
output(2, 187) <= input(43);
output(2, 188) <= input(45);
output(2, 189) <= input(46);
output(2, 190) <= input(49);
output(2, 191) <= input(50);
output(2, 192) <= input(11);
output(2, 193) <= input(12);
output(2, 194) <= input(13);
output(2, 195) <= input(14);
output(2, 196) <= input(15);
output(2, 197) <= input(32);
output(2, 198) <= input(34);
output(2, 199) <= input(36);
output(2, 200) <= input(37);
output(2, 201) <= input(40);
output(2, 202) <= input(42);
output(2, 203) <= input(44);
output(2, 204) <= input(47);
output(2, 205) <= input(48);
output(2, 206) <= input(51);
output(2, 207) <= input(52);
output(2, 208) <= input(12);
output(2, 209) <= input(13);
output(2, 210) <= input(14);
output(2, 211) <= input(15);
output(2, 212) <= input(32);
output(2, 213) <= input(34);
output(2, 214) <= input(36);
output(2, 215) <= input(37);
output(2, 216) <= input(40);
output(2, 217) <= input(42);
output(2, 218) <= input(44);
output(2, 219) <= input(47);
output(2, 220) <= input(48);
output(2, 221) <= input(51);
output(2, 222) <= input(52);
output(2, 223) <= input(53);
output(2, 224) <= input(28);
output(2, 225) <= input(29);
output(2, 226) <= input(30);
output(2, 227) <= input(31);
output(2, 228) <= input(33);
output(2, 229) <= input(35);
output(2, 230) <= input(38);
output(2, 231) <= input(39);
output(2, 232) <= input(41);
output(2, 233) <= input(43);
output(2, 234) <= input(45);
output(2, 235) <= input(46);
output(2, 236) <= input(49);
output(2, 237) <= input(50);
output(2, 238) <= input(54);
output(2, 239) <= input(55);
output(2, 240) <= input(29);
output(2, 241) <= input(30);
output(2, 242) <= input(31);
output(2, 243) <= input(33);
output(2, 244) <= input(35);
output(2, 245) <= input(38);
output(2, 246) <= input(39);
output(2, 247) <= input(41);
output(2, 248) <= input(43);
output(2, 249) <= input(45);
output(2, 250) <= input(46);
output(2, 251) <= input(49);
output(2, 252) <= input(50);
output(2, 253) <= input(54);
output(2, 254) <= input(55);
output(2, 255) <= input(56);
output(3, 0) <= input(4);
output(3, 1) <= input(5);
output(3, 2) <= input(6);
output(3, 3) <= input(7);
output(3, 4) <= input(8);
output(3, 5) <= input(9);
output(3, 6) <= input(10);
output(3, 7) <= input(11);
output(3, 8) <= input(12);
output(3, 9) <= input(13);
output(3, 10) <= input(14);
output(3, 11) <= input(15);
output(3, 12) <= input(32);
output(3, 13) <= input(34);
output(3, 14) <= input(36);
output(3, 15) <= input(37);
output(3, 16) <= input(5);
output(3, 17) <= input(6);
output(3, 18) <= input(7);
output(3, 19) <= input(8);
output(3, 20) <= input(9);
output(3, 21) <= input(10);
output(3, 22) <= input(11);
output(3, 23) <= input(12);
output(3, 24) <= input(13);
output(3, 25) <= input(14);
output(3, 26) <= input(15);
output(3, 27) <= input(32);
output(3, 28) <= input(34);
output(3, 29) <= input(36);
output(3, 30) <= input(37);
output(3, 31) <= input(40);
output(3, 32) <= input(21);
output(3, 33) <= input(22);
output(3, 34) <= input(23);
output(3, 35) <= input(24);
output(3, 36) <= input(25);
output(3, 37) <= input(26);
output(3, 38) <= input(27);
output(3, 39) <= input(28);
output(3, 40) <= input(29);
output(3, 41) <= input(30);
output(3, 42) <= input(31);
output(3, 43) <= input(33);
output(3, 44) <= input(35);
output(3, 45) <= input(38);
output(3, 46) <= input(39);
output(3, 47) <= input(41);
output(3, 48) <= input(22);
output(3, 49) <= input(23);
output(3, 50) <= input(24);
output(3, 51) <= input(25);
output(3, 52) <= input(26);
output(3, 53) <= input(27);
output(3, 54) <= input(28);
output(3, 55) <= input(29);
output(3, 56) <= input(30);
output(3, 57) <= input(31);
output(3, 58) <= input(33);
output(3, 59) <= input(35);
output(3, 60) <= input(38);
output(3, 61) <= input(39);
output(3, 62) <= input(41);
output(3, 63) <= input(43);
output(3, 64) <= input(23);
output(3, 65) <= input(24);
output(3, 66) <= input(25);
output(3, 67) <= input(26);
output(3, 68) <= input(27);
output(3, 69) <= input(28);
output(3, 70) <= input(29);
output(3, 71) <= input(30);
output(3, 72) <= input(31);
output(3, 73) <= input(33);
output(3, 74) <= input(35);
output(3, 75) <= input(38);
output(3, 76) <= input(39);
output(3, 77) <= input(41);
output(3, 78) <= input(43);
output(3, 79) <= input(45);
output(3, 80) <= input(8);
output(3, 81) <= input(9);
output(3, 82) <= input(10);
output(3, 83) <= input(11);
output(3, 84) <= input(12);
output(3, 85) <= input(13);
output(3, 86) <= input(14);
output(3, 87) <= input(15);
output(3, 88) <= input(32);
output(3, 89) <= input(34);
output(3, 90) <= input(36);
output(3, 91) <= input(37);
output(3, 92) <= input(40);
output(3, 93) <= input(42);
output(3, 94) <= input(44);
output(3, 95) <= input(47);
output(3, 96) <= input(9);
output(3, 97) <= input(10);
output(3, 98) <= input(11);
output(3, 99) <= input(12);
output(3, 100) <= input(13);
output(3, 101) <= input(14);
output(3, 102) <= input(15);
output(3, 103) <= input(32);
output(3, 104) <= input(34);
output(3, 105) <= input(36);
output(3, 106) <= input(37);
output(3, 107) <= input(40);
output(3, 108) <= input(42);
output(3, 109) <= input(44);
output(3, 110) <= input(47);
output(3, 111) <= input(48);
output(3, 112) <= input(10);
output(3, 113) <= input(11);
output(3, 114) <= input(12);
output(3, 115) <= input(13);
output(3, 116) <= input(14);
output(3, 117) <= input(15);
output(3, 118) <= input(32);
output(3, 119) <= input(34);
output(3, 120) <= input(36);
output(3, 121) <= input(37);
output(3, 122) <= input(40);
output(3, 123) <= input(42);
output(3, 124) <= input(44);
output(3, 125) <= input(47);
output(3, 126) <= input(48);
output(3, 127) <= input(51);
output(3, 128) <= input(26);
output(3, 129) <= input(27);
output(3, 130) <= input(28);
output(3, 131) <= input(29);
output(3, 132) <= input(30);
output(3, 133) <= input(31);
output(3, 134) <= input(33);
output(3, 135) <= input(35);
output(3, 136) <= input(38);
output(3, 137) <= input(39);
output(3, 138) <= input(41);
output(3, 139) <= input(43);
output(3, 140) <= input(45);
output(3, 141) <= input(46);
output(3, 142) <= input(49);
output(3, 143) <= input(50);
output(3, 144) <= input(27);
output(3, 145) <= input(28);
output(3, 146) <= input(29);
output(3, 147) <= input(30);
output(3, 148) <= input(31);
output(3, 149) <= input(33);
output(3, 150) <= input(35);
output(3, 151) <= input(38);
output(3, 152) <= input(39);
output(3, 153) <= input(41);
output(3, 154) <= input(43);
output(3, 155) <= input(45);
output(3, 156) <= input(46);
output(3, 157) <= input(49);
output(3, 158) <= input(50);
output(3, 159) <= input(54);
output(3, 160) <= input(12);
output(3, 161) <= input(13);
output(3, 162) <= input(14);
output(3, 163) <= input(15);
output(3, 164) <= input(32);
output(3, 165) <= input(34);
output(3, 166) <= input(36);
output(3, 167) <= input(37);
output(3, 168) <= input(40);
output(3, 169) <= input(42);
output(3, 170) <= input(44);
output(3, 171) <= input(47);
output(3, 172) <= input(48);
output(3, 173) <= input(51);
output(3, 174) <= input(52);
output(3, 175) <= input(53);
output(3, 176) <= input(13);
output(3, 177) <= input(14);
output(3, 178) <= input(15);
output(3, 179) <= input(32);
output(3, 180) <= input(34);
output(3, 181) <= input(36);
output(3, 182) <= input(37);
output(3, 183) <= input(40);
output(3, 184) <= input(42);
output(3, 185) <= input(44);
output(3, 186) <= input(47);
output(3, 187) <= input(48);
output(3, 188) <= input(51);
output(3, 189) <= input(52);
output(3, 190) <= input(53);
output(3, 191) <= input(57);
output(3, 192) <= input(14);
output(3, 193) <= input(15);
output(3, 194) <= input(32);
output(3, 195) <= input(34);
output(3, 196) <= input(36);
output(3, 197) <= input(37);
output(3, 198) <= input(40);
output(3, 199) <= input(42);
output(3, 200) <= input(44);
output(3, 201) <= input(47);
output(3, 202) <= input(48);
output(3, 203) <= input(51);
output(3, 204) <= input(52);
output(3, 205) <= input(53);
output(3, 206) <= input(57);
output(3, 207) <= input(58);
output(3, 208) <= input(30);
output(3, 209) <= input(31);
output(3, 210) <= input(33);
output(3, 211) <= input(35);
output(3, 212) <= input(38);
output(3, 213) <= input(39);
output(3, 214) <= input(41);
output(3, 215) <= input(43);
output(3, 216) <= input(45);
output(3, 217) <= input(46);
output(3, 218) <= input(49);
output(3, 219) <= input(50);
output(3, 220) <= input(54);
output(3, 221) <= input(55);
output(3, 222) <= input(56);
output(3, 223) <= input(59);
output(3, 224) <= input(31);
output(3, 225) <= input(33);
output(3, 226) <= input(35);
output(3, 227) <= input(38);
output(3, 228) <= input(39);
output(3, 229) <= input(41);
output(3, 230) <= input(43);
output(3, 231) <= input(45);
output(3, 232) <= input(46);
output(3, 233) <= input(49);
output(3, 234) <= input(50);
output(3, 235) <= input(54);
output(3, 236) <= input(55);
output(3, 237) <= input(56);
output(3, 238) <= input(59);
output(3, 239) <= input(60);
output(3, 240) <= input(33);
output(3, 241) <= input(35);
output(3, 242) <= input(38);
output(3, 243) <= input(39);
output(3, 244) <= input(41);
output(3, 245) <= input(43);
output(3, 246) <= input(45);
output(3, 247) <= input(46);
output(3, 248) <= input(49);
output(3, 249) <= input(50);
output(3, 250) <= input(54);
output(3, 251) <= input(55);
output(3, 252) <= input(56);
output(3, 253) <= input(59);
output(3, 254) <= input(60);
output(3, 255) <= input(61);
output(4, 0) <= input(21);
output(4, 1) <= input(22);
output(4, 2) <= input(23);
output(4, 3) <= input(24);
output(4, 4) <= input(25);
output(4, 5) <= input(26);
output(4, 6) <= input(27);
output(4, 7) <= input(28);
output(4, 8) <= input(29);
output(4, 9) <= input(30);
output(4, 10) <= input(31);
output(4, 11) <= input(33);
output(4, 12) <= input(35);
output(4, 13) <= input(38);
output(4, 14) <= input(39);
output(4, 15) <= input(41);
output(4, 16) <= input(22);
output(4, 17) <= input(23);
output(4, 18) <= input(24);
output(4, 19) <= input(25);
output(4, 20) <= input(26);
output(4, 21) <= input(27);
output(4, 22) <= input(28);
output(4, 23) <= input(29);
output(4, 24) <= input(30);
output(4, 25) <= input(31);
output(4, 26) <= input(33);
output(4, 27) <= input(35);
output(4, 28) <= input(38);
output(4, 29) <= input(39);
output(4, 30) <= input(41);
output(4, 31) <= input(43);
output(4, 32) <= input(23);
output(4, 33) <= input(24);
output(4, 34) <= input(25);
output(4, 35) <= input(26);
output(4, 36) <= input(27);
output(4, 37) <= input(28);
output(4, 38) <= input(29);
output(4, 39) <= input(30);
output(4, 40) <= input(31);
output(4, 41) <= input(33);
output(4, 42) <= input(35);
output(4, 43) <= input(38);
output(4, 44) <= input(39);
output(4, 45) <= input(41);
output(4, 46) <= input(43);
output(4, 47) <= input(45);
output(4, 48) <= input(24);
output(4, 49) <= input(25);
output(4, 50) <= input(26);
output(4, 51) <= input(27);
output(4, 52) <= input(28);
output(4, 53) <= input(29);
output(4, 54) <= input(30);
output(4, 55) <= input(31);
output(4, 56) <= input(33);
output(4, 57) <= input(35);
output(4, 58) <= input(38);
output(4, 59) <= input(39);
output(4, 60) <= input(41);
output(4, 61) <= input(43);
output(4, 62) <= input(45);
output(4, 63) <= input(46);
output(4, 64) <= input(25);
output(4, 65) <= input(26);
output(4, 66) <= input(27);
output(4, 67) <= input(28);
output(4, 68) <= input(29);
output(4, 69) <= input(30);
output(4, 70) <= input(31);
output(4, 71) <= input(33);
output(4, 72) <= input(35);
output(4, 73) <= input(38);
output(4, 74) <= input(39);
output(4, 75) <= input(41);
output(4, 76) <= input(43);
output(4, 77) <= input(45);
output(4, 78) <= input(46);
output(4, 79) <= input(49);
output(4, 80) <= input(10);
output(4, 81) <= input(11);
output(4, 82) <= input(12);
output(4, 83) <= input(13);
output(4, 84) <= input(14);
output(4, 85) <= input(15);
output(4, 86) <= input(32);
output(4, 87) <= input(34);
output(4, 88) <= input(36);
output(4, 89) <= input(37);
output(4, 90) <= input(40);
output(4, 91) <= input(42);
output(4, 92) <= input(44);
output(4, 93) <= input(47);
output(4, 94) <= input(48);
output(4, 95) <= input(51);
output(4, 96) <= input(11);
output(4, 97) <= input(12);
output(4, 98) <= input(13);
output(4, 99) <= input(14);
output(4, 100) <= input(15);
output(4, 101) <= input(32);
output(4, 102) <= input(34);
output(4, 103) <= input(36);
output(4, 104) <= input(37);
output(4, 105) <= input(40);
output(4, 106) <= input(42);
output(4, 107) <= input(44);
output(4, 108) <= input(47);
output(4, 109) <= input(48);
output(4, 110) <= input(51);
output(4, 111) <= input(52);
output(4, 112) <= input(12);
output(4, 113) <= input(13);
output(4, 114) <= input(14);
output(4, 115) <= input(15);
output(4, 116) <= input(32);
output(4, 117) <= input(34);
output(4, 118) <= input(36);
output(4, 119) <= input(37);
output(4, 120) <= input(40);
output(4, 121) <= input(42);
output(4, 122) <= input(44);
output(4, 123) <= input(47);
output(4, 124) <= input(48);
output(4, 125) <= input(51);
output(4, 126) <= input(52);
output(4, 127) <= input(53);
output(4, 128) <= input(13);
output(4, 129) <= input(14);
output(4, 130) <= input(15);
output(4, 131) <= input(32);
output(4, 132) <= input(34);
output(4, 133) <= input(36);
output(4, 134) <= input(37);
output(4, 135) <= input(40);
output(4, 136) <= input(42);
output(4, 137) <= input(44);
output(4, 138) <= input(47);
output(4, 139) <= input(48);
output(4, 140) <= input(51);
output(4, 141) <= input(52);
output(4, 142) <= input(53);
output(4, 143) <= input(57);
output(4, 144) <= input(14);
output(4, 145) <= input(15);
output(4, 146) <= input(32);
output(4, 147) <= input(34);
output(4, 148) <= input(36);
output(4, 149) <= input(37);
output(4, 150) <= input(40);
output(4, 151) <= input(42);
output(4, 152) <= input(44);
output(4, 153) <= input(47);
output(4, 154) <= input(48);
output(4, 155) <= input(51);
output(4, 156) <= input(52);
output(4, 157) <= input(53);
output(4, 158) <= input(57);
output(4, 159) <= input(58);
output(4, 160) <= input(30);
output(4, 161) <= input(31);
output(4, 162) <= input(33);
output(4, 163) <= input(35);
output(4, 164) <= input(38);
output(4, 165) <= input(39);
output(4, 166) <= input(41);
output(4, 167) <= input(43);
output(4, 168) <= input(45);
output(4, 169) <= input(46);
output(4, 170) <= input(49);
output(4, 171) <= input(50);
output(4, 172) <= input(54);
output(4, 173) <= input(55);
output(4, 174) <= input(56);
output(4, 175) <= input(59);
output(4, 176) <= input(31);
output(4, 177) <= input(33);
output(4, 178) <= input(35);
output(4, 179) <= input(38);
output(4, 180) <= input(39);
output(4, 181) <= input(41);
output(4, 182) <= input(43);
output(4, 183) <= input(45);
output(4, 184) <= input(46);
output(4, 185) <= input(49);
output(4, 186) <= input(50);
output(4, 187) <= input(54);
output(4, 188) <= input(55);
output(4, 189) <= input(56);
output(4, 190) <= input(59);
output(4, 191) <= input(60);
output(4, 192) <= input(33);
output(4, 193) <= input(35);
output(4, 194) <= input(38);
output(4, 195) <= input(39);
output(4, 196) <= input(41);
output(4, 197) <= input(43);
output(4, 198) <= input(45);
output(4, 199) <= input(46);
output(4, 200) <= input(49);
output(4, 201) <= input(50);
output(4, 202) <= input(54);
output(4, 203) <= input(55);
output(4, 204) <= input(56);
output(4, 205) <= input(59);
output(4, 206) <= input(60);
output(4, 207) <= input(61);
output(4, 208) <= input(35);
output(4, 209) <= input(38);
output(4, 210) <= input(39);
output(4, 211) <= input(41);
output(4, 212) <= input(43);
output(4, 213) <= input(45);
output(4, 214) <= input(46);
output(4, 215) <= input(49);
output(4, 216) <= input(50);
output(4, 217) <= input(54);
output(4, 218) <= input(55);
output(4, 219) <= input(56);
output(4, 220) <= input(59);
output(4, 221) <= input(60);
output(4, 222) <= input(61);
output(4, 223) <= input(62);
output(4, 224) <= input(38);
output(4, 225) <= input(39);
output(4, 226) <= input(41);
output(4, 227) <= input(43);
output(4, 228) <= input(45);
output(4, 229) <= input(46);
output(4, 230) <= input(49);
output(4, 231) <= input(50);
output(4, 232) <= input(54);
output(4, 233) <= input(55);
output(4, 234) <= input(56);
output(4, 235) <= input(59);
output(4, 236) <= input(60);
output(4, 237) <= input(61);
output(4, 238) <= input(62);
output(4, 239) <= input(63);
output(4, 240) <= input(39);
output(4, 241) <= input(41);
output(4, 242) <= input(43);
output(4, 243) <= input(45);
output(4, 244) <= input(46);
output(4, 245) <= input(49);
output(4, 246) <= input(50);
output(4, 247) <= input(54);
output(4, 248) <= input(55);
output(4, 249) <= input(56);
output(4, 250) <= input(59);
output(4, 251) <= input(60);
output(4, 252) <= input(61);
output(4, 253) <= input(62);
output(4, 254) <= input(63);
output(4, 255) <= input(64);
output(5, 0) <= input(23);
output(5, 1) <= input(24);
output(5, 2) <= input(25);
output(5, 3) <= input(26);
output(5, 4) <= input(27);
output(5, 5) <= input(28);
output(5, 6) <= input(29);
output(5, 7) <= input(30);
output(5, 8) <= input(31);
output(5, 9) <= input(33);
output(5, 10) <= input(35);
output(5, 11) <= input(38);
output(5, 12) <= input(39);
output(5, 13) <= input(41);
output(5, 14) <= input(43);
output(5, 15) <= input(45);
output(5, 16) <= input(24);
output(5, 17) <= input(25);
output(5, 18) <= input(26);
output(5, 19) <= input(27);
output(5, 20) <= input(28);
output(5, 21) <= input(29);
output(5, 22) <= input(30);
output(5, 23) <= input(31);
output(5, 24) <= input(33);
output(5, 25) <= input(35);
output(5, 26) <= input(38);
output(5, 27) <= input(39);
output(5, 28) <= input(41);
output(5, 29) <= input(43);
output(5, 30) <= input(45);
output(5, 31) <= input(46);
output(5, 32) <= input(25);
output(5, 33) <= input(26);
output(5, 34) <= input(27);
output(5, 35) <= input(28);
output(5, 36) <= input(29);
output(5, 37) <= input(30);
output(5, 38) <= input(31);
output(5, 39) <= input(33);
output(5, 40) <= input(35);
output(5, 41) <= input(38);
output(5, 42) <= input(39);
output(5, 43) <= input(41);
output(5, 44) <= input(43);
output(5, 45) <= input(45);
output(5, 46) <= input(46);
output(5, 47) <= input(49);
output(5, 48) <= input(26);
output(5, 49) <= input(27);
output(5, 50) <= input(28);
output(5, 51) <= input(29);
output(5, 52) <= input(30);
output(5, 53) <= input(31);
output(5, 54) <= input(33);
output(5, 55) <= input(35);
output(5, 56) <= input(38);
output(5, 57) <= input(39);
output(5, 58) <= input(41);
output(5, 59) <= input(43);
output(5, 60) <= input(45);
output(5, 61) <= input(46);
output(5, 62) <= input(49);
output(5, 63) <= input(50);
output(5, 64) <= input(27);
output(5, 65) <= input(28);
output(5, 66) <= input(29);
output(5, 67) <= input(30);
output(5, 68) <= input(31);
output(5, 69) <= input(33);
output(5, 70) <= input(35);
output(5, 71) <= input(38);
output(5, 72) <= input(39);
output(5, 73) <= input(41);
output(5, 74) <= input(43);
output(5, 75) <= input(45);
output(5, 76) <= input(46);
output(5, 77) <= input(49);
output(5, 78) <= input(50);
output(5, 79) <= input(54);
output(5, 80) <= input(28);
output(5, 81) <= input(29);
output(5, 82) <= input(30);
output(5, 83) <= input(31);
output(5, 84) <= input(33);
output(5, 85) <= input(35);
output(5, 86) <= input(38);
output(5, 87) <= input(39);
output(5, 88) <= input(41);
output(5, 89) <= input(43);
output(5, 90) <= input(45);
output(5, 91) <= input(46);
output(5, 92) <= input(49);
output(5, 93) <= input(50);
output(5, 94) <= input(54);
output(5, 95) <= input(55);
output(5, 96) <= input(29);
output(5, 97) <= input(30);
output(5, 98) <= input(31);
output(5, 99) <= input(33);
output(5, 100) <= input(35);
output(5, 101) <= input(38);
output(5, 102) <= input(39);
output(5, 103) <= input(41);
output(5, 104) <= input(43);
output(5, 105) <= input(45);
output(5, 106) <= input(46);
output(5, 107) <= input(49);
output(5, 108) <= input(50);
output(5, 109) <= input(54);
output(5, 110) <= input(55);
output(5, 111) <= input(56);
output(5, 112) <= input(30);
output(5, 113) <= input(31);
output(5, 114) <= input(33);
output(5, 115) <= input(35);
output(5, 116) <= input(38);
output(5, 117) <= input(39);
output(5, 118) <= input(41);
output(5, 119) <= input(43);
output(5, 120) <= input(45);
output(5, 121) <= input(46);
output(5, 122) <= input(49);
output(5, 123) <= input(50);
output(5, 124) <= input(54);
output(5, 125) <= input(55);
output(5, 126) <= input(56);
output(5, 127) <= input(59);
output(5, 128) <= input(31);
output(5, 129) <= input(33);
output(5, 130) <= input(35);
output(5, 131) <= input(38);
output(5, 132) <= input(39);
output(5, 133) <= input(41);
output(5, 134) <= input(43);
output(5, 135) <= input(45);
output(5, 136) <= input(46);
output(5, 137) <= input(49);
output(5, 138) <= input(50);
output(5, 139) <= input(54);
output(5, 140) <= input(55);
output(5, 141) <= input(56);
output(5, 142) <= input(59);
output(5, 143) <= input(60);
output(5, 144) <= input(33);
output(5, 145) <= input(35);
output(5, 146) <= input(38);
output(5, 147) <= input(39);
output(5, 148) <= input(41);
output(5, 149) <= input(43);
output(5, 150) <= input(45);
output(5, 151) <= input(46);
output(5, 152) <= input(49);
output(5, 153) <= input(50);
output(5, 154) <= input(54);
output(5, 155) <= input(55);
output(5, 156) <= input(56);
output(5, 157) <= input(59);
output(5, 158) <= input(60);
output(5, 159) <= input(61);
output(5, 160) <= input(35);
output(5, 161) <= input(38);
output(5, 162) <= input(39);
output(5, 163) <= input(41);
output(5, 164) <= input(43);
output(5, 165) <= input(45);
output(5, 166) <= input(46);
output(5, 167) <= input(49);
output(5, 168) <= input(50);
output(5, 169) <= input(54);
output(5, 170) <= input(55);
output(5, 171) <= input(56);
output(5, 172) <= input(59);
output(5, 173) <= input(60);
output(5, 174) <= input(61);
output(5, 175) <= input(62);
output(5, 176) <= input(38);
output(5, 177) <= input(39);
output(5, 178) <= input(41);
output(5, 179) <= input(43);
output(5, 180) <= input(45);
output(5, 181) <= input(46);
output(5, 182) <= input(49);
output(5, 183) <= input(50);
output(5, 184) <= input(54);
output(5, 185) <= input(55);
output(5, 186) <= input(56);
output(5, 187) <= input(59);
output(5, 188) <= input(60);
output(5, 189) <= input(61);
output(5, 190) <= input(62);
output(5, 191) <= input(63);
output(5, 192) <= input(39);
output(5, 193) <= input(41);
output(5, 194) <= input(43);
output(5, 195) <= input(45);
output(5, 196) <= input(46);
output(5, 197) <= input(49);
output(5, 198) <= input(50);
output(5, 199) <= input(54);
output(5, 200) <= input(55);
output(5, 201) <= input(56);
output(5, 202) <= input(59);
output(5, 203) <= input(60);
output(5, 204) <= input(61);
output(5, 205) <= input(62);
output(5, 206) <= input(63);
output(5, 207) <= input(64);
output(5, 208) <= input(41);
output(5, 209) <= input(43);
output(5, 210) <= input(45);
output(5, 211) <= input(46);
output(5, 212) <= input(49);
output(5, 213) <= input(50);
output(5, 214) <= input(54);
output(5, 215) <= input(55);
output(5, 216) <= input(56);
output(5, 217) <= input(59);
output(5, 218) <= input(60);
output(5, 219) <= input(61);
output(5, 220) <= input(62);
output(5, 221) <= input(63);
output(5, 222) <= input(64);
output(5, 223) <= input(65);
output(5, 224) <= input(43);
output(5, 225) <= input(45);
output(5, 226) <= input(46);
output(5, 227) <= input(49);
output(5, 228) <= input(50);
output(5, 229) <= input(54);
output(5, 230) <= input(55);
output(5, 231) <= input(56);
output(5, 232) <= input(59);
output(5, 233) <= input(60);
output(5, 234) <= input(61);
output(5, 235) <= input(62);
output(5, 236) <= input(63);
output(5, 237) <= input(64);
output(5, 238) <= input(65);
output(5, 239) <= input(66);
output(5, 240) <= input(45);
output(5, 241) <= input(46);
output(5, 242) <= input(49);
output(5, 243) <= input(50);
output(5, 244) <= input(54);
output(5, 245) <= input(55);
output(5, 246) <= input(56);
output(5, 247) <= input(59);
output(5, 248) <= input(60);
output(5, 249) <= input(61);
output(5, 250) <= input(62);
output(5, 251) <= input(63);
output(5, 252) <= input(64);
output(5, 253) <= input(65);
output(5, 254) <= input(66);
output(5, 255) <= input(67);
when others => for i in 0 to 7 loop for j in 0 to 255 loop output(i,j) <= "00000000"; end loop; end loop;
end case;
elsif control = "101" then 
case iteration_control is
when "0000" =>
output(0, 0) <= input(0);
output(0, 1) <= input(1);
output(0, 2) <= input(2);
output(0, 3) <= input(3);
output(0, 4) <= input(4);
output(0, 5) <= input(5);
output(0, 6) <= input(6);
output(0, 7) <= input(7);
output(0, 8) <= input(8);
output(0, 9) <= input(9);
output(0, 10) <= input(10);
output(0, 11) <= input(11);
output(0, 12) <= input(12);
output(0, 13) <= input(13);
output(0, 14) <= input(14);
output(0, 15) <= input(15);
output(0, 16) <= input(1);
output(0, 17) <= input(2);
output(0, 18) <= input(3);
output(0, 19) <= input(4);
output(0, 20) <= input(5);
output(0, 21) <= input(6);
output(0, 22) <= input(7);
output(0, 23) <= input(8);
output(0, 24) <= input(9);
output(0, 25) <= input(10);
output(0, 26) <= input(11);
output(0, 27) <= input(12);
output(0, 28) <= input(13);
output(0, 29) <= input(14);
output(0, 30) <= input(15);
output(0, 31) <= input(16);
output(0, 32) <= input(2);
output(0, 33) <= input(3);
output(0, 34) <= input(4);
output(0, 35) <= input(5);
output(0, 36) <= input(6);
output(0, 37) <= input(7);
output(0, 38) <= input(8);
output(0, 39) <= input(9);
output(0, 40) <= input(10);
output(0, 41) <= input(11);
output(0, 42) <= input(12);
output(0, 43) <= input(13);
output(0, 44) <= input(14);
output(0, 45) <= input(15);
output(0, 46) <= input(16);
output(0, 47) <= input(17);
output(0, 48) <= input(3);
output(0, 49) <= input(4);
output(0, 50) <= input(5);
output(0, 51) <= input(6);
output(0, 52) <= input(7);
output(0, 53) <= input(8);
output(0, 54) <= input(9);
output(0, 55) <= input(10);
output(0, 56) <= input(11);
output(0, 57) <= input(12);
output(0, 58) <= input(13);
output(0, 59) <= input(14);
output(0, 60) <= input(15);
output(0, 61) <= input(16);
output(0, 62) <= input(17);
output(0, 63) <= input(18);
output(0, 64) <= input(4);
output(0, 65) <= input(5);
output(0, 66) <= input(6);
output(0, 67) <= input(7);
output(0, 68) <= input(8);
output(0, 69) <= input(9);
output(0, 70) <= input(10);
output(0, 71) <= input(11);
output(0, 72) <= input(12);
output(0, 73) <= input(13);
output(0, 74) <= input(14);
output(0, 75) <= input(15);
output(0, 76) <= input(16);
output(0, 77) <= input(17);
output(0, 78) <= input(18);
output(0, 79) <= input(19);
output(0, 80) <= input(5);
output(0, 81) <= input(6);
output(0, 82) <= input(7);
output(0, 83) <= input(8);
output(0, 84) <= input(9);
output(0, 85) <= input(10);
output(0, 86) <= input(11);
output(0, 87) <= input(12);
output(0, 88) <= input(13);
output(0, 89) <= input(14);
output(0, 90) <= input(15);
output(0, 91) <= input(16);
output(0, 92) <= input(17);
output(0, 93) <= input(18);
output(0, 94) <= input(19);
output(0, 95) <= input(20);
output(0, 96) <= input(6);
output(0, 97) <= input(7);
output(0, 98) <= input(8);
output(0, 99) <= input(9);
output(0, 100) <= input(10);
output(0, 101) <= input(11);
output(0, 102) <= input(12);
output(0, 103) <= input(13);
output(0, 104) <= input(14);
output(0, 105) <= input(15);
output(0, 106) <= input(16);
output(0, 107) <= input(17);
output(0, 108) <= input(18);
output(0, 109) <= input(19);
output(0, 110) <= input(20);
output(0, 111) <= input(21);
output(0, 112) <= input(7);
output(0, 113) <= input(8);
output(0, 114) <= input(9);
output(0, 115) <= input(10);
output(0, 116) <= input(11);
output(0, 117) <= input(12);
output(0, 118) <= input(13);
output(0, 119) <= input(14);
output(0, 120) <= input(15);
output(0, 121) <= input(16);
output(0, 122) <= input(17);
output(0, 123) <= input(18);
output(0, 124) <= input(19);
output(0, 125) <= input(20);
output(0, 126) <= input(21);
output(0, 127) <= input(22);
output(0, 128) <= input(8);
output(0, 129) <= input(9);
output(0, 130) <= input(10);
output(0, 131) <= input(11);
output(0, 132) <= input(12);
output(0, 133) <= input(13);
output(0, 134) <= input(14);
output(0, 135) <= input(15);
output(0, 136) <= input(16);
output(0, 137) <= input(17);
output(0, 138) <= input(18);
output(0, 139) <= input(19);
output(0, 140) <= input(20);
output(0, 141) <= input(21);
output(0, 142) <= input(22);
output(0, 143) <= input(23);
output(0, 144) <= input(9);
output(0, 145) <= input(10);
output(0, 146) <= input(11);
output(0, 147) <= input(12);
output(0, 148) <= input(13);
output(0, 149) <= input(14);
output(0, 150) <= input(15);
output(0, 151) <= input(16);
output(0, 152) <= input(17);
output(0, 153) <= input(18);
output(0, 154) <= input(19);
output(0, 155) <= input(20);
output(0, 156) <= input(21);
output(0, 157) <= input(22);
output(0, 158) <= input(23);
output(0, 159) <= input(24);
output(0, 160) <= input(10);
output(0, 161) <= input(11);
output(0, 162) <= input(12);
output(0, 163) <= input(13);
output(0, 164) <= input(14);
output(0, 165) <= input(15);
output(0, 166) <= input(16);
output(0, 167) <= input(17);
output(0, 168) <= input(18);
output(0, 169) <= input(19);
output(0, 170) <= input(20);
output(0, 171) <= input(21);
output(0, 172) <= input(22);
output(0, 173) <= input(23);
output(0, 174) <= input(24);
output(0, 175) <= input(25);
output(0, 176) <= input(11);
output(0, 177) <= input(12);
output(0, 178) <= input(13);
output(0, 179) <= input(14);
output(0, 180) <= input(15);
output(0, 181) <= input(16);
output(0, 182) <= input(17);
output(0, 183) <= input(18);
output(0, 184) <= input(19);
output(0, 185) <= input(20);
output(0, 186) <= input(21);
output(0, 187) <= input(22);
output(0, 188) <= input(23);
output(0, 189) <= input(24);
output(0, 190) <= input(25);
output(0, 191) <= input(26);
output(0, 192) <= input(12);
output(0, 193) <= input(13);
output(0, 194) <= input(14);
output(0, 195) <= input(15);
output(0, 196) <= input(16);
output(0, 197) <= input(17);
output(0, 198) <= input(18);
output(0, 199) <= input(19);
output(0, 200) <= input(20);
output(0, 201) <= input(21);
output(0, 202) <= input(22);
output(0, 203) <= input(23);
output(0, 204) <= input(24);
output(0, 205) <= input(25);
output(0, 206) <= input(26);
output(0, 207) <= input(27);
output(0, 208) <= input(13);
output(0, 209) <= input(14);
output(0, 210) <= input(15);
output(0, 211) <= input(16);
output(0, 212) <= input(17);
output(0, 213) <= input(18);
output(0, 214) <= input(19);
output(0, 215) <= input(20);
output(0, 216) <= input(21);
output(0, 217) <= input(22);
output(0, 218) <= input(23);
output(0, 219) <= input(24);
output(0, 220) <= input(25);
output(0, 221) <= input(26);
output(0, 222) <= input(27);
output(0, 223) <= input(28);
output(0, 224) <= input(14);
output(0, 225) <= input(15);
output(0, 226) <= input(16);
output(0, 227) <= input(17);
output(0, 228) <= input(18);
output(0, 229) <= input(19);
output(0, 230) <= input(20);
output(0, 231) <= input(21);
output(0, 232) <= input(22);
output(0, 233) <= input(23);
output(0, 234) <= input(24);
output(0, 235) <= input(25);
output(0, 236) <= input(26);
output(0, 237) <= input(27);
output(0, 238) <= input(28);
output(0, 239) <= input(29);
output(0, 240) <= input(15);
output(0, 241) <= input(16);
output(0, 242) <= input(17);
output(0, 243) <= input(18);
output(0, 244) <= input(19);
output(0, 245) <= input(20);
output(0, 246) <= input(21);
output(0, 247) <= input(22);
output(0, 248) <= input(23);
output(0, 249) <= input(24);
output(0, 250) <= input(25);
output(0, 251) <= input(26);
output(0, 252) <= input(27);
output(0, 253) <= input(28);
output(0, 254) <= input(29);
output(0, 255) <= input(30);
output(1, 0) <= input(31);
output(1, 1) <= input(32);
output(1, 2) <= input(0);
output(1, 3) <= input(1);
output(1, 4) <= input(2);
output(1, 5) <= input(3);
output(1, 6) <= input(4);
output(1, 7) <= input(5);
output(1, 8) <= input(6);
output(1, 9) <= input(7);
output(1, 10) <= input(8);
output(1, 11) <= input(9);
output(1, 12) <= input(10);
output(1, 13) <= input(11);
output(1, 14) <= input(12);
output(1, 15) <= input(13);
output(1, 16) <= input(32);
output(1, 17) <= input(0);
output(1, 18) <= input(1);
output(1, 19) <= input(2);
output(1, 20) <= input(3);
output(1, 21) <= input(4);
output(1, 22) <= input(5);
output(1, 23) <= input(6);
output(1, 24) <= input(7);
output(1, 25) <= input(8);
output(1, 26) <= input(9);
output(1, 27) <= input(10);
output(1, 28) <= input(11);
output(1, 29) <= input(12);
output(1, 30) <= input(13);
output(1, 31) <= input(14);
output(1, 32) <= input(0);
output(1, 33) <= input(1);
output(1, 34) <= input(2);
output(1, 35) <= input(3);
output(1, 36) <= input(4);
output(1, 37) <= input(5);
output(1, 38) <= input(6);
output(1, 39) <= input(7);
output(1, 40) <= input(8);
output(1, 41) <= input(9);
output(1, 42) <= input(10);
output(1, 43) <= input(11);
output(1, 44) <= input(12);
output(1, 45) <= input(13);
output(1, 46) <= input(14);
output(1, 47) <= input(15);
output(1, 48) <= input(1);
output(1, 49) <= input(2);
output(1, 50) <= input(3);
output(1, 51) <= input(4);
output(1, 52) <= input(5);
output(1, 53) <= input(6);
output(1, 54) <= input(7);
output(1, 55) <= input(8);
output(1, 56) <= input(9);
output(1, 57) <= input(10);
output(1, 58) <= input(11);
output(1, 59) <= input(12);
output(1, 60) <= input(13);
output(1, 61) <= input(14);
output(1, 62) <= input(15);
output(1, 63) <= input(16);
output(1, 64) <= input(2);
output(1, 65) <= input(3);
output(1, 66) <= input(4);
output(1, 67) <= input(5);
output(1, 68) <= input(6);
output(1, 69) <= input(7);
output(1, 70) <= input(8);
output(1, 71) <= input(9);
output(1, 72) <= input(10);
output(1, 73) <= input(11);
output(1, 74) <= input(12);
output(1, 75) <= input(13);
output(1, 76) <= input(14);
output(1, 77) <= input(15);
output(1, 78) <= input(16);
output(1, 79) <= input(17);
output(1, 80) <= input(33);
output(1, 81) <= input(34);
output(1, 82) <= input(35);
output(1, 83) <= input(36);
output(1, 84) <= input(37);
output(1, 85) <= input(38);
output(1, 86) <= input(39);
output(1, 87) <= input(40);
output(1, 88) <= input(41);
output(1, 89) <= input(42);
output(1, 90) <= input(43);
output(1, 91) <= input(44);
output(1, 92) <= input(45);
output(1, 93) <= input(46);
output(1, 94) <= input(47);
output(1, 95) <= input(48);
output(1, 96) <= input(34);
output(1, 97) <= input(35);
output(1, 98) <= input(36);
output(1, 99) <= input(37);
output(1, 100) <= input(38);
output(1, 101) <= input(39);
output(1, 102) <= input(40);
output(1, 103) <= input(41);
output(1, 104) <= input(42);
output(1, 105) <= input(43);
output(1, 106) <= input(44);
output(1, 107) <= input(45);
output(1, 108) <= input(46);
output(1, 109) <= input(47);
output(1, 110) <= input(48);
output(1, 111) <= input(49);
output(1, 112) <= input(35);
output(1, 113) <= input(36);
output(1, 114) <= input(37);
output(1, 115) <= input(38);
output(1, 116) <= input(39);
output(1, 117) <= input(40);
output(1, 118) <= input(41);
output(1, 119) <= input(42);
output(1, 120) <= input(43);
output(1, 121) <= input(44);
output(1, 122) <= input(45);
output(1, 123) <= input(46);
output(1, 124) <= input(47);
output(1, 125) <= input(48);
output(1, 126) <= input(49);
output(1, 127) <= input(50);
output(1, 128) <= input(36);
output(1, 129) <= input(37);
output(1, 130) <= input(38);
output(1, 131) <= input(39);
output(1, 132) <= input(40);
output(1, 133) <= input(41);
output(1, 134) <= input(42);
output(1, 135) <= input(43);
output(1, 136) <= input(44);
output(1, 137) <= input(45);
output(1, 138) <= input(46);
output(1, 139) <= input(47);
output(1, 140) <= input(48);
output(1, 141) <= input(49);
output(1, 142) <= input(50);
output(1, 143) <= input(51);
output(1, 144) <= input(37);
output(1, 145) <= input(38);
output(1, 146) <= input(39);
output(1, 147) <= input(40);
output(1, 148) <= input(41);
output(1, 149) <= input(42);
output(1, 150) <= input(43);
output(1, 151) <= input(44);
output(1, 152) <= input(45);
output(1, 153) <= input(46);
output(1, 154) <= input(47);
output(1, 155) <= input(48);
output(1, 156) <= input(49);
output(1, 157) <= input(50);
output(1, 158) <= input(51);
output(1, 159) <= input(52);
output(1, 160) <= input(7);
output(1, 161) <= input(8);
output(1, 162) <= input(9);
output(1, 163) <= input(10);
output(1, 164) <= input(11);
output(1, 165) <= input(12);
output(1, 166) <= input(13);
output(1, 167) <= input(14);
output(1, 168) <= input(15);
output(1, 169) <= input(16);
output(1, 170) <= input(17);
output(1, 171) <= input(18);
output(1, 172) <= input(19);
output(1, 173) <= input(20);
output(1, 174) <= input(21);
output(1, 175) <= input(22);
output(1, 176) <= input(8);
output(1, 177) <= input(9);
output(1, 178) <= input(10);
output(1, 179) <= input(11);
output(1, 180) <= input(12);
output(1, 181) <= input(13);
output(1, 182) <= input(14);
output(1, 183) <= input(15);
output(1, 184) <= input(16);
output(1, 185) <= input(17);
output(1, 186) <= input(18);
output(1, 187) <= input(19);
output(1, 188) <= input(20);
output(1, 189) <= input(21);
output(1, 190) <= input(22);
output(1, 191) <= input(23);
output(1, 192) <= input(9);
output(1, 193) <= input(10);
output(1, 194) <= input(11);
output(1, 195) <= input(12);
output(1, 196) <= input(13);
output(1, 197) <= input(14);
output(1, 198) <= input(15);
output(1, 199) <= input(16);
output(1, 200) <= input(17);
output(1, 201) <= input(18);
output(1, 202) <= input(19);
output(1, 203) <= input(20);
output(1, 204) <= input(21);
output(1, 205) <= input(22);
output(1, 206) <= input(23);
output(1, 207) <= input(24);
output(1, 208) <= input(10);
output(1, 209) <= input(11);
output(1, 210) <= input(12);
output(1, 211) <= input(13);
output(1, 212) <= input(14);
output(1, 213) <= input(15);
output(1, 214) <= input(16);
output(1, 215) <= input(17);
output(1, 216) <= input(18);
output(1, 217) <= input(19);
output(1, 218) <= input(20);
output(1, 219) <= input(21);
output(1, 220) <= input(22);
output(1, 221) <= input(23);
output(1, 222) <= input(24);
output(1, 223) <= input(25);
output(1, 224) <= input(11);
output(1, 225) <= input(12);
output(1, 226) <= input(13);
output(1, 227) <= input(14);
output(1, 228) <= input(15);
output(1, 229) <= input(16);
output(1, 230) <= input(17);
output(1, 231) <= input(18);
output(1, 232) <= input(19);
output(1, 233) <= input(20);
output(1, 234) <= input(21);
output(1, 235) <= input(22);
output(1, 236) <= input(23);
output(1, 237) <= input(24);
output(1, 238) <= input(25);
output(1, 239) <= input(26);
output(1, 240) <= input(12);
output(1, 241) <= input(13);
output(1, 242) <= input(14);
output(1, 243) <= input(15);
output(1, 244) <= input(16);
output(1, 245) <= input(17);
output(1, 246) <= input(18);
output(1, 247) <= input(19);
output(1, 248) <= input(20);
output(1, 249) <= input(21);
output(1, 250) <= input(22);
output(1, 251) <= input(23);
output(1, 252) <= input(24);
output(1, 253) <= input(25);
output(1, 254) <= input(26);
output(1, 255) <= input(27);
output(2, 0) <= input(53);
output(2, 1) <= input(54);
output(2, 2) <= input(55);
output(2, 3) <= input(56);
output(2, 4) <= input(57);
output(2, 5) <= input(58);
output(2, 6) <= input(33);
output(2, 7) <= input(34);
output(2, 8) <= input(35);
output(2, 9) <= input(36);
output(2, 10) <= input(37);
output(2, 11) <= input(38);
output(2, 12) <= input(39);
output(2, 13) <= input(40);
output(2, 14) <= input(41);
output(2, 15) <= input(42);
output(2, 16) <= input(54);
output(2, 17) <= input(55);
output(2, 18) <= input(56);
output(2, 19) <= input(57);
output(2, 20) <= input(58);
output(2, 21) <= input(33);
output(2, 22) <= input(34);
output(2, 23) <= input(35);
output(2, 24) <= input(36);
output(2, 25) <= input(37);
output(2, 26) <= input(38);
output(2, 27) <= input(39);
output(2, 28) <= input(40);
output(2, 29) <= input(41);
output(2, 30) <= input(42);
output(2, 31) <= input(43);
output(2, 32) <= input(31);
output(2, 33) <= input(32);
output(2, 34) <= input(0);
output(2, 35) <= input(1);
output(2, 36) <= input(2);
output(2, 37) <= input(3);
output(2, 38) <= input(4);
output(2, 39) <= input(5);
output(2, 40) <= input(6);
output(2, 41) <= input(7);
output(2, 42) <= input(8);
output(2, 43) <= input(9);
output(2, 44) <= input(10);
output(2, 45) <= input(11);
output(2, 46) <= input(12);
output(2, 47) <= input(13);
output(2, 48) <= input(32);
output(2, 49) <= input(0);
output(2, 50) <= input(1);
output(2, 51) <= input(2);
output(2, 52) <= input(3);
output(2, 53) <= input(4);
output(2, 54) <= input(5);
output(2, 55) <= input(6);
output(2, 56) <= input(7);
output(2, 57) <= input(8);
output(2, 58) <= input(9);
output(2, 59) <= input(10);
output(2, 60) <= input(11);
output(2, 61) <= input(12);
output(2, 62) <= input(13);
output(2, 63) <= input(14);
output(2, 64) <= input(0);
output(2, 65) <= input(1);
output(2, 66) <= input(2);
output(2, 67) <= input(3);
output(2, 68) <= input(4);
output(2, 69) <= input(5);
output(2, 70) <= input(6);
output(2, 71) <= input(7);
output(2, 72) <= input(8);
output(2, 73) <= input(9);
output(2, 74) <= input(10);
output(2, 75) <= input(11);
output(2, 76) <= input(12);
output(2, 77) <= input(13);
output(2, 78) <= input(14);
output(2, 79) <= input(15);
output(2, 80) <= input(57);
output(2, 81) <= input(58);
output(2, 82) <= input(33);
output(2, 83) <= input(34);
output(2, 84) <= input(35);
output(2, 85) <= input(36);
output(2, 86) <= input(37);
output(2, 87) <= input(38);
output(2, 88) <= input(39);
output(2, 89) <= input(40);
output(2, 90) <= input(41);
output(2, 91) <= input(42);
output(2, 92) <= input(43);
output(2, 93) <= input(44);
output(2, 94) <= input(45);
output(2, 95) <= input(46);
output(2, 96) <= input(58);
output(2, 97) <= input(33);
output(2, 98) <= input(34);
output(2, 99) <= input(35);
output(2, 100) <= input(36);
output(2, 101) <= input(37);
output(2, 102) <= input(38);
output(2, 103) <= input(39);
output(2, 104) <= input(40);
output(2, 105) <= input(41);
output(2, 106) <= input(42);
output(2, 107) <= input(43);
output(2, 108) <= input(44);
output(2, 109) <= input(45);
output(2, 110) <= input(46);
output(2, 111) <= input(47);
output(2, 112) <= input(33);
output(2, 113) <= input(34);
output(2, 114) <= input(35);
output(2, 115) <= input(36);
output(2, 116) <= input(37);
output(2, 117) <= input(38);
output(2, 118) <= input(39);
output(2, 119) <= input(40);
output(2, 120) <= input(41);
output(2, 121) <= input(42);
output(2, 122) <= input(43);
output(2, 123) <= input(44);
output(2, 124) <= input(45);
output(2, 125) <= input(46);
output(2, 126) <= input(47);
output(2, 127) <= input(48);
output(2, 128) <= input(3);
output(2, 129) <= input(4);
output(2, 130) <= input(5);
output(2, 131) <= input(6);
output(2, 132) <= input(7);
output(2, 133) <= input(8);
output(2, 134) <= input(9);
output(2, 135) <= input(10);
output(2, 136) <= input(11);
output(2, 137) <= input(12);
output(2, 138) <= input(13);
output(2, 139) <= input(14);
output(2, 140) <= input(15);
output(2, 141) <= input(16);
output(2, 142) <= input(17);
output(2, 143) <= input(18);
output(2, 144) <= input(4);
output(2, 145) <= input(5);
output(2, 146) <= input(6);
output(2, 147) <= input(7);
output(2, 148) <= input(8);
output(2, 149) <= input(9);
output(2, 150) <= input(10);
output(2, 151) <= input(11);
output(2, 152) <= input(12);
output(2, 153) <= input(13);
output(2, 154) <= input(14);
output(2, 155) <= input(15);
output(2, 156) <= input(16);
output(2, 157) <= input(17);
output(2, 158) <= input(18);
output(2, 159) <= input(19);
output(2, 160) <= input(35);
output(2, 161) <= input(36);
output(2, 162) <= input(37);
output(2, 163) <= input(38);
output(2, 164) <= input(39);
output(2, 165) <= input(40);
output(2, 166) <= input(41);
output(2, 167) <= input(42);
output(2, 168) <= input(43);
output(2, 169) <= input(44);
output(2, 170) <= input(45);
output(2, 171) <= input(46);
output(2, 172) <= input(47);
output(2, 173) <= input(48);
output(2, 174) <= input(49);
output(2, 175) <= input(50);
output(2, 176) <= input(36);
output(2, 177) <= input(37);
output(2, 178) <= input(38);
output(2, 179) <= input(39);
output(2, 180) <= input(40);
output(2, 181) <= input(41);
output(2, 182) <= input(42);
output(2, 183) <= input(43);
output(2, 184) <= input(44);
output(2, 185) <= input(45);
output(2, 186) <= input(46);
output(2, 187) <= input(47);
output(2, 188) <= input(48);
output(2, 189) <= input(49);
output(2, 190) <= input(50);
output(2, 191) <= input(51);
output(2, 192) <= input(37);
output(2, 193) <= input(38);
output(2, 194) <= input(39);
output(2, 195) <= input(40);
output(2, 196) <= input(41);
output(2, 197) <= input(42);
output(2, 198) <= input(43);
output(2, 199) <= input(44);
output(2, 200) <= input(45);
output(2, 201) <= input(46);
output(2, 202) <= input(47);
output(2, 203) <= input(48);
output(2, 204) <= input(49);
output(2, 205) <= input(50);
output(2, 206) <= input(51);
output(2, 207) <= input(52);
output(2, 208) <= input(7);
output(2, 209) <= input(8);
output(2, 210) <= input(9);
output(2, 211) <= input(10);
output(2, 212) <= input(11);
output(2, 213) <= input(12);
output(2, 214) <= input(13);
output(2, 215) <= input(14);
output(2, 216) <= input(15);
output(2, 217) <= input(16);
output(2, 218) <= input(17);
output(2, 219) <= input(18);
output(2, 220) <= input(19);
output(2, 221) <= input(20);
output(2, 222) <= input(21);
output(2, 223) <= input(22);
output(2, 224) <= input(8);
output(2, 225) <= input(9);
output(2, 226) <= input(10);
output(2, 227) <= input(11);
output(2, 228) <= input(12);
output(2, 229) <= input(13);
output(2, 230) <= input(14);
output(2, 231) <= input(15);
output(2, 232) <= input(16);
output(2, 233) <= input(17);
output(2, 234) <= input(18);
output(2, 235) <= input(19);
output(2, 236) <= input(20);
output(2, 237) <= input(21);
output(2, 238) <= input(22);
output(2, 239) <= input(23);
output(2, 240) <= input(9);
output(2, 241) <= input(10);
output(2, 242) <= input(11);
output(2, 243) <= input(12);
output(2, 244) <= input(13);
output(2, 245) <= input(14);
output(2, 246) <= input(15);
output(2, 247) <= input(16);
output(2, 248) <= input(17);
output(2, 249) <= input(18);
output(2, 250) <= input(19);
output(2, 251) <= input(20);
output(2, 252) <= input(21);
output(2, 253) <= input(22);
output(2, 254) <= input(23);
output(2, 255) <= input(24);
output(3, 0) <= input(59);
output(3, 1) <= input(60);
output(3, 2) <= input(61);
output(3, 3) <= input(31);
output(3, 4) <= input(32);
output(3, 5) <= input(0);
output(3, 6) <= input(1);
output(3, 7) <= input(2);
output(3, 8) <= input(3);
output(3, 9) <= input(4);
output(3, 10) <= input(5);
output(3, 11) <= input(6);
output(3, 12) <= input(7);
output(3, 13) <= input(8);
output(3, 14) <= input(9);
output(3, 15) <= input(10);
output(3, 16) <= input(62);
output(3, 17) <= input(53);
output(3, 18) <= input(54);
output(3, 19) <= input(55);
output(3, 20) <= input(56);
output(3, 21) <= input(57);
output(3, 22) <= input(58);
output(3, 23) <= input(33);
output(3, 24) <= input(34);
output(3, 25) <= input(35);
output(3, 26) <= input(36);
output(3, 27) <= input(37);
output(3, 28) <= input(38);
output(3, 29) <= input(39);
output(3, 30) <= input(40);
output(3, 31) <= input(41);
output(3, 32) <= input(53);
output(3, 33) <= input(54);
output(3, 34) <= input(55);
output(3, 35) <= input(56);
output(3, 36) <= input(57);
output(3, 37) <= input(58);
output(3, 38) <= input(33);
output(3, 39) <= input(34);
output(3, 40) <= input(35);
output(3, 41) <= input(36);
output(3, 42) <= input(37);
output(3, 43) <= input(38);
output(3, 44) <= input(39);
output(3, 45) <= input(40);
output(3, 46) <= input(41);
output(3, 47) <= input(42);
output(3, 48) <= input(61);
output(3, 49) <= input(31);
output(3, 50) <= input(32);
output(3, 51) <= input(0);
output(3, 52) <= input(1);
output(3, 53) <= input(2);
output(3, 54) <= input(3);
output(3, 55) <= input(4);
output(3, 56) <= input(5);
output(3, 57) <= input(6);
output(3, 58) <= input(7);
output(3, 59) <= input(8);
output(3, 60) <= input(9);
output(3, 61) <= input(10);
output(3, 62) <= input(11);
output(3, 63) <= input(12);
output(3, 64) <= input(31);
output(3, 65) <= input(32);
output(3, 66) <= input(0);
output(3, 67) <= input(1);
output(3, 68) <= input(2);
output(3, 69) <= input(3);
output(3, 70) <= input(4);
output(3, 71) <= input(5);
output(3, 72) <= input(6);
output(3, 73) <= input(7);
output(3, 74) <= input(8);
output(3, 75) <= input(9);
output(3, 76) <= input(10);
output(3, 77) <= input(11);
output(3, 78) <= input(12);
output(3, 79) <= input(13);
output(3, 80) <= input(55);
output(3, 81) <= input(56);
output(3, 82) <= input(57);
output(3, 83) <= input(58);
output(3, 84) <= input(33);
output(3, 85) <= input(34);
output(3, 86) <= input(35);
output(3, 87) <= input(36);
output(3, 88) <= input(37);
output(3, 89) <= input(38);
output(3, 90) <= input(39);
output(3, 91) <= input(40);
output(3, 92) <= input(41);
output(3, 93) <= input(42);
output(3, 94) <= input(43);
output(3, 95) <= input(44);
output(3, 96) <= input(56);
output(3, 97) <= input(57);
output(3, 98) <= input(58);
output(3, 99) <= input(33);
output(3, 100) <= input(34);
output(3, 101) <= input(35);
output(3, 102) <= input(36);
output(3, 103) <= input(37);
output(3, 104) <= input(38);
output(3, 105) <= input(39);
output(3, 106) <= input(40);
output(3, 107) <= input(41);
output(3, 108) <= input(42);
output(3, 109) <= input(43);
output(3, 110) <= input(44);
output(3, 111) <= input(45);
output(3, 112) <= input(0);
output(3, 113) <= input(1);
output(3, 114) <= input(2);
output(3, 115) <= input(3);
output(3, 116) <= input(4);
output(3, 117) <= input(5);
output(3, 118) <= input(6);
output(3, 119) <= input(7);
output(3, 120) <= input(8);
output(3, 121) <= input(9);
output(3, 122) <= input(10);
output(3, 123) <= input(11);
output(3, 124) <= input(12);
output(3, 125) <= input(13);
output(3, 126) <= input(14);
output(3, 127) <= input(15);
output(3, 128) <= input(57);
output(3, 129) <= input(58);
output(3, 130) <= input(33);
output(3, 131) <= input(34);
output(3, 132) <= input(35);
output(3, 133) <= input(36);
output(3, 134) <= input(37);
output(3, 135) <= input(38);
output(3, 136) <= input(39);
output(3, 137) <= input(40);
output(3, 138) <= input(41);
output(3, 139) <= input(42);
output(3, 140) <= input(43);
output(3, 141) <= input(44);
output(3, 142) <= input(45);
output(3, 143) <= input(46);
output(3, 144) <= input(58);
output(3, 145) <= input(33);
output(3, 146) <= input(34);
output(3, 147) <= input(35);
output(3, 148) <= input(36);
output(3, 149) <= input(37);
output(3, 150) <= input(38);
output(3, 151) <= input(39);
output(3, 152) <= input(40);
output(3, 153) <= input(41);
output(3, 154) <= input(42);
output(3, 155) <= input(43);
output(3, 156) <= input(44);
output(3, 157) <= input(45);
output(3, 158) <= input(46);
output(3, 159) <= input(47);
output(3, 160) <= input(2);
output(3, 161) <= input(3);
output(3, 162) <= input(4);
output(3, 163) <= input(5);
output(3, 164) <= input(6);
output(3, 165) <= input(7);
output(3, 166) <= input(8);
output(3, 167) <= input(9);
output(3, 168) <= input(10);
output(3, 169) <= input(11);
output(3, 170) <= input(12);
output(3, 171) <= input(13);
output(3, 172) <= input(14);
output(3, 173) <= input(15);
output(3, 174) <= input(16);
output(3, 175) <= input(17);
output(3, 176) <= input(3);
output(3, 177) <= input(4);
output(3, 178) <= input(5);
output(3, 179) <= input(6);
output(3, 180) <= input(7);
output(3, 181) <= input(8);
output(3, 182) <= input(9);
output(3, 183) <= input(10);
output(3, 184) <= input(11);
output(3, 185) <= input(12);
output(3, 186) <= input(13);
output(3, 187) <= input(14);
output(3, 188) <= input(15);
output(3, 189) <= input(16);
output(3, 190) <= input(17);
output(3, 191) <= input(18);
output(3, 192) <= input(34);
output(3, 193) <= input(35);
output(3, 194) <= input(36);
output(3, 195) <= input(37);
output(3, 196) <= input(38);
output(3, 197) <= input(39);
output(3, 198) <= input(40);
output(3, 199) <= input(41);
output(3, 200) <= input(42);
output(3, 201) <= input(43);
output(3, 202) <= input(44);
output(3, 203) <= input(45);
output(3, 204) <= input(46);
output(3, 205) <= input(47);
output(3, 206) <= input(48);
output(3, 207) <= input(49);
output(3, 208) <= input(35);
output(3, 209) <= input(36);
output(3, 210) <= input(37);
output(3, 211) <= input(38);
output(3, 212) <= input(39);
output(3, 213) <= input(40);
output(3, 214) <= input(41);
output(3, 215) <= input(42);
output(3, 216) <= input(43);
output(3, 217) <= input(44);
output(3, 218) <= input(45);
output(3, 219) <= input(46);
output(3, 220) <= input(47);
output(3, 221) <= input(48);
output(3, 222) <= input(49);
output(3, 223) <= input(50);
output(3, 224) <= input(5);
output(3, 225) <= input(6);
output(3, 226) <= input(7);
output(3, 227) <= input(8);
output(3, 228) <= input(9);
output(3, 229) <= input(10);
output(3, 230) <= input(11);
output(3, 231) <= input(12);
output(3, 232) <= input(13);
output(3, 233) <= input(14);
output(3, 234) <= input(15);
output(3, 235) <= input(16);
output(3, 236) <= input(17);
output(3, 237) <= input(18);
output(3, 238) <= input(19);
output(3, 239) <= input(20);
output(3, 240) <= input(6);
output(3, 241) <= input(7);
output(3, 242) <= input(8);
output(3, 243) <= input(9);
output(3, 244) <= input(10);
output(3, 245) <= input(11);
output(3, 246) <= input(12);
output(3, 247) <= input(13);
output(3, 248) <= input(14);
output(3, 249) <= input(15);
output(3, 250) <= input(16);
output(3, 251) <= input(17);
output(3, 252) <= input(18);
output(3, 253) <= input(19);
output(3, 254) <= input(20);
output(3, 255) <= input(21);
output(4, 0) <= input(63);
output(4, 1) <= input(64);
output(4, 2) <= input(62);
output(4, 3) <= input(53);
output(4, 4) <= input(54);
output(4, 5) <= input(55);
output(4, 6) <= input(56);
output(4, 7) <= input(57);
output(4, 8) <= input(58);
output(4, 9) <= input(33);
output(4, 10) <= input(34);
output(4, 11) <= input(35);
output(4, 12) <= input(36);
output(4, 13) <= input(37);
output(4, 14) <= input(38);
output(4, 15) <= input(39);
output(4, 16) <= input(65);
output(4, 17) <= input(59);
output(4, 18) <= input(60);
output(4, 19) <= input(61);
output(4, 20) <= input(31);
output(4, 21) <= input(32);
output(4, 22) <= input(0);
output(4, 23) <= input(1);
output(4, 24) <= input(2);
output(4, 25) <= input(3);
output(4, 26) <= input(4);
output(4, 27) <= input(5);
output(4, 28) <= input(6);
output(4, 29) <= input(7);
output(4, 30) <= input(8);
output(4, 31) <= input(9);
output(4, 32) <= input(64);
output(4, 33) <= input(62);
output(4, 34) <= input(53);
output(4, 35) <= input(54);
output(4, 36) <= input(55);
output(4, 37) <= input(56);
output(4, 38) <= input(57);
output(4, 39) <= input(58);
output(4, 40) <= input(33);
output(4, 41) <= input(34);
output(4, 42) <= input(35);
output(4, 43) <= input(36);
output(4, 44) <= input(37);
output(4, 45) <= input(38);
output(4, 46) <= input(39);
output(4, 47) <= input(40);
output(4, 48) <= input(62);
output(4, 49) <= input(53);
output(4, 50) <= input(54);
output(4, 51) <= input(55);
output(4, 52) <= input(56);
output(4, 53) <= input(57);
output(4, 54) <= input(58);
output(4, 55) <= input(33);
output(4, 56) <= input(34);
output(4, 57) <= input(35);
output(4, 58) <= input(36);
output(4, 59) <= input(37);
output(4, 60) <= input(38);
output(4, 61) <= input(39);
output(4, 62) <= input(40);
output(4, 63) <= input(41);
output(4, 64) <= input(60);
output(4, 65) <= input(61);
output(4, 66) <= input(31);
output(4, 67) <= input(32);
output(4, 68) <= input(0);
output(4, 69) <= input(1);
output(4, 70) <= input(2);
output(4, 71) <= input(3);
output(4, 72) <= input(4);
output(4, 73) <= input(5);
output(4, 74) <= input(6);
output(4, 75) <= input(7);
output(4, 76) <= input(8);
output(4, 77) <= input(9);
output(4, 78) <= input(10);
output(4, 79) <= input(11);
output(4, 80) <= input(53);
output(4, 81) <= input(54);
output(4, 82) <= input(55);
output(4, 83) <= input(56);
output(4, 84) <= input(57);
output(4, 85) <= input(58);
output(4, 86) <= input(33);
output(4, 87) <= input(34);
output(4, 88) <= input(35);
output(4, 89) <= input(36);
output(4, 90) <= input(37);
output(4, 91) <= input(38);
output(4, 92) <= input(39);
output(4, 93) <= input(40);
output(4, 94) <= input(41);
output(4, 95) <= input(42);
output(4, 96) <= input(61);
output(4, 97) <= input(31);
output(4, 98) <= input(32);
output(4, 99) <= input(0);
output(4, 100) <= input(1);
output(4, 101) <= input(2);
output(4, 102) <= input(3);
output(4, 103) <= input(4);
output(4, 104) <= input(5);
output(4, 105) <= input(6);
output(4, 106) <= input(7);
output(4, 107) <= input(8);
output(4, 108) <= input(9);
output(4, 109) <= input(10);
output(4, 110) <= input(11);
output(4, 111) <= input(12);
output(4, 112) <= input(31);
output(4, 113) <= input(32);
output(4, 114) <= input(0);
output(4, 115) <= input(1);
output(4, 116) <= input(2);
output(4, 117) <= input(3);
output(4, 118) <= input(4);
output(4, 119) <= input(5);
output(4, 120) <= input(6);
output(4, 121) <= input(7);
output(4, 122) <= input(8);
output(4, 123) <= input(9);
output(4, 124) <= input(10);
output(4, 125) <= input(11);
output(4, 126) <= input(12);
output(4, 127) <= input(13);
output(4, 128) <= input(55);
output(4, 129) <= input(56);
output(4, 130) <= input(57);
output(4, 131) <= input(58);
output(4, 132) <= input(33);
output(4, 133) <= input(34);
output(4, 134) <= input(35);
output(4, 135) <= input(36);
output(4, 136) <= input(37);
output(4, 137) <= input(38);
output(4, 138) <= input(39);
output(4, 139) <= input(40);
output(4, 140) <= input(41);
output(4, 141) <= input(42);
output(4, 142) <= input(43);
output(4, 143) <= input(44);
output(4, 144) <= input(32);
output(4, 145) <= input(0);
output(4, 146) <= input(1);
output(4, 147) <= input(2);
output(4, 148) <= input(3);
output(4, 149) <= input(4);
output(4, 150) <= input(5);
output(4, 151) <= input(6);
output(4, 152) <= input(7);
output(4, 153) <= input(8);
output(4, 154) <= input(9);
output(4, 155) <= input(10);
output(4, 156) <= input(11);
output(4, 157) <= input(12);
output(4, 158) <= input(13);
output(4, 159) <= input(14);
output(4, 160) <= input(56);
output(4, 161) <= input(57);
output(4, 162) <= input(58);
output(4, 163) <= input(33);
output(4, 164) <= input(34);
output(4, 165) <= input(35);
output(4, 166) <= input(36);
output(4, 167) <= input(37);
output(4, 168) <= input(38);
output(4, 169) <= input(39);
output(4, 170) <= input(40);
output(4, 171) <= input(41);
output(4, 172) <= input(42);
output(4, 173) <= input(43);
output(4, 174) <= input(44);
output(4, 175) <= input(45);
output(4, 176) <= input(57);
output(4, 177) <= input(58);
output(4, 178) <= input(33);
output(4, 179) <= input(34);
output(4, 180) <= input(35);
output(4, 181) <= input(36);
output(4, 182) <= input(37);
output(4, 183) <= input(38);
output(4, 184) <= input(39);
output(4, 185) <= input(40);
output(4, 186) <= input(41);
output(4, 187) <= input(42);
output(4, 188) <= input(43);
output(4, 189) <= input(44);
output(4, 190) <= input(45);
output(4, 191) <= input(46);
output(4, 192) <= input(1);
output(4, 193) <= input(2);
output(4, 194) <= input(3);
output(4, 195) <= input(4);
output(4, 196) <= input(5);
output(4, 197) <= input(6);
output(4, 198) <= input(7);
output(4, 199) <= input(8);
output(4, 200) <= input(9);
output(4, 201) <= input(10);
output(4, 202) <= input(11);
output(4, 203) <= input(12);
output(4, 204) <= input(13);
output(4, 205) <= input(14);
output(4, 206) <= input(15);
output(4, 207) <= input(16);
output(4, 208) <= input(58);
output(4, 209) <= input(33);
output(4, 210) <= input(34);
output(4, 211) <= input(35);
output(4, 212) <= input(36);
output(4, 213) <= input(37);
output(4, 214) <= input(38);
output(4, 215) <= input(39);
output(4, 216) <= input(40);
output(4, 217) <= input(41);
output(4, 218) <= input(42);
output(4, 219) <= input(43);
output(4, 220) <= input(44);
output(4, 221) <= input(45);
output(4, 222) <= input(46);
output(4, 223) <= input(47);
output(4, 224) <= input(2);
output(4, 225) <= input(3);
output(4, 226) <= input(4);
output(4, 227) <= input(5);
output(4, 228) <= input(6);
output(4, 229) <= input(7);
output(4, 230) <= input(8);
output(4, 231) <= input(9);
output(4, 232) <= input(10);
output(4, 233) <= input(11);
output(4, 234) <= input(12);
output(4, 235) <= input(13);
output(4, 236) <= input(14);
output(4, 237) <= input(15);
output(4, 238) <= input(16);
output(4, 239) <= input(17);
output(4, 240) <= input(3);
output(4, 241) <= input(4);
output(4, 242) <= input(5);
output(4, 243) <= input(6);
output(4, 244) <= input(7);
output(4, 245) <= input(8);
output(4, 246) <= input(9);
output(4, 247) <= input(10);
output(4, 248) <= input(11);
output(4, 249) <= input(12);
output(4, 250) <= input(13);
output(4, 251) <= input(14);
output(4, 252) <= input(15);
output(4, 253) <= input(16);
output(4, 254) <= input(17);
output(4, 255) <= input(18);
output(5, 0) <= input(66);
output(5, 1) <= input(63);
output(5, 2) <= input(64);
output(5, 3) <= input(62);
output(5, 4) <= input(53);
output(5, 5) <= input(54);
output(5, 6) <= input(55);
output(5, 7) <= input(56);
output(5, 8) <= input(57);
output(5, 9) <= input(58);
output(5, 10) <= input(33);
output(5, 11) <= input(34);
output(5, 12) <= input(35);
output(5, 13) <= input(36);
output(5, 14) <= input(37);
output(5, 15) <= input(38);
output(5, 16) <= input(67);
output(5, 17) <= input(65);
output(5, 18) <= input(59);
output(5, 19) <= input(60);
output(5, 20) <= input(61);
output(5, 21) <= input(31);
output(5, 22) <= input(32);
output(5, 23) <= input(0);
output(5, 24) <= input(1);
output(5, 25) <= input(2);
output(5, 26) <= input(3);
output(5, 27) <= input(4);
output(5, 28) <= input(5);
output(5, 29) <= input(6);
output(5, 30) <= input(7);
output(5, 31) <= input(8);
output(5, 32) <= input(63);
output(5, 33) <= input(64);
output(5, 34) <= input(62);
output(5, 35) <= input(53);
output(5, 36) <= input(54);
output(5, 37) <= input(55);
output(5, 38) <= input(56);
output(5, 39) <= input(57);
output(5, 40) <= input(58);
output(5, 41) <= input(33);
output(5, 42) <= input(34);
output(5, 43) <= input(35);
output(5, 44) <= input(36);
output(5, 45) <= input(37);
output(5, 46) <= input(38);
output(5, 47) <= input(39);
output(5, 48) <= input(65);
output(5, 49) <= input(59);
output(5, 50) <= input(60);
output(5, 51) <= input(61);
output(5, 52) <= input(31);
output(5, 53) <= input(32);
output(5, 54) <= input(0);
output(5, 55) <= input(1);
output(5, 56) <= input(2);
output(5, 57) <= input(3);
output(5, 58) <= input(4);
output(5, 59) <= input(5);
output(5, 60) <= input(6);
output(5, 61) <= input(7);
output(5, 62) <= input(8);
output(5, 63) <= input(9);
output(5, 64) <= input(64);
output(5, 65) <= input(62);
output(5, 66) <= input(53);
output(5, 67) <= input(54);
output(5, 68) <= input(55);
output(5, 69) <= input(56);
output(5, 70) <= input(57);
output(5, 71) <= input(58);
output(5, 72) <= input(33);
output(5, 73) <= input(34);
output(5, 74) <= input(35);
output(5, 75) <= input(36);
output(5, 76) <= input(37);
output(5, 77) <= input(38);
output(5, 78) <= input(39);
output(5, 79) <= input(40);
output(5, 80) <= input(59);
output(5, 81) <= input(60);
output(5, 82) <= input(61);
output(5, 83) <= input(31);
output(5, 84) <= input(32);
output(5, 85) <= input(0);
output(5, 86) <= input(1);
output(5, 87) <= input(2);
output(5, 88) <= input(3);
output(5, 89) <= input(4);
output(5, 90) <= input(5);
output(5, 91) <= input(6);
output(5, 92) <= input(7);
output(5, 93) <= input(8);
output(5, 94) <= input(9);
output(5, 95) <= input(10);
output(5, 96) <= input(62);
output(5, 97) <= input(53);
output(5, 98) <= input(54);
output(5, 99) <= input(55);
output(5, 100) <= input(56);
output(5, 101) <= input(57);
output(5, 102) <= input(58);
output(5, 103) <= input(33);
output(5, 104) <= input(34);
output(5, 105) <= input(35);
output(5, 106) <= input(36);
output(5, 107) <= input(37);
output(5, 108) <= input(38);
output(5, 109) <= input(39);
output(5, 110) <= input(40);
output(5, 111) <= input(41);
output(5, 112) <= input(53);
output(5, 113) <= input(54);
output(5, 114) <= input(55);
output(5, 115) <= input(56);
output(5, 116) <= input(57);
output(5, 117) <= input(58);
output(5, 118) <= input(33);
output(5, 119) <= input(34);
output(5, 120) <= input(35);
output(5, 121) <= input(36);
output(5, 122) <= input(37);
output(5, 123) <= input(38);
output(5, 124) <= input(39);
output(5, 125) <= input(40);
output(5, 126) <= input(41);
output(5, 127) <= input(42);
output(5, 128) <= input(61);
output(5, 129) <= input(31);
output(5, 130) <= input(32);
output(5, 131) <= input(0);
output(5, 132) <= input(1);
output(5, 133) <= input(2);
output(5, 134) <= input(3);
output(5, 135) <= input(4);
output(5, 136) <= input(5);
output(5, 137) <= input(6);
output(5, 138) <= input(7);
output(5, 139) <= input(8);
output(5, 140) <= input(9);
output(5, 141) <= input(10);
output(5, 142) <= input(11);
output(5, 143) <= input(12);
output(5, 144) <= input(54);
output(5, 145) <= input(55);
output(5, 146) <= input(56);
output(5, 147) <= input(57);
output(5, 148) <= input(58);
output(5, 149) <= input(33);
output(5, 150) <= input(34);
output(5, 151) <= input(35);
output(5, 152) <= input(36);
output(5, 153) <= input(37);
output(5, 154) <= input(38);
output(5, 155) <= input(39);
output(5, 156) <= input(40);
output(5, 157) <= input(41);
output(5, 158) <= input(42);
output(5, 159) <= input(43);
output(5, 160) <= input(31);
output(5, 161) <= input(32);
output(5, 162) <= input(0);
output(5, 163) <= input(1);
output(5, 164) <= input(2);
output(5, 165) <= input(3);
output(5, 166) <= input(4);
output(5, 167) <= input(5);
output(5, 168) <= input(6);
output(5, 169) <= input(7);
output(5, 170) <= input(8);
output(5, 171) <= input(9);
output(5, 172) <= input(10);
output(5, 173) <= input(11);
output(5, 174) <= input(12);
output(5, 175) <= input(13);
output(5, 176) <= input(55);
output(5, 177) <= input(56);
output(5, 178) <= input(57);
output(5, 179) <= input(58);
output(5, 180) <= input(33);
output(5, 181) <= input(34);
output(5, 182) <= input(35);
output(5, 183) <= input(36);
output(5, 184) <= input(37);
output(5, 185) <= input(38);
output(5, 186) <= input(39);
output(5, 187) <= input(40);
output(5, 188) <= input(41);
output(5, 189) <= input(42);
output(5, 190) <= input(43);
output(5, 191) <= input(44);
output(5, 192) <= input(32);
output(5, 193) <= input(0);
output(5, 194) <= input(1);
output(5, 195) <= input(2);
output(5, 196) <= input(3);
output(5, 197) <= input(4);
output(5, 198) <= input(5);
output(5, 199) <= input(6);
output(5, 200) <= input(7);
output(5, 201) <= input(8);
output(5, 202) <= input(9);
output(5, 203) <= input(10);
output(5, 204) <= input(11);
output(5, 205) <= input(12);
output(5, 206) <= input(13);
output(5, 207) <= input(14);
output(5, 208) <= input(56);
output(5, 209) <= input(57);
output(5, 210) <= input(58);
output(5, 211) <= input(33);
output(5, 212) <= input(34);
output(5, 213) <= input(35);
output(5, 214) <= input(36);
output(5, 215) <= input(37);
output(5, 216) <= input(38);
output(5, 217) <= input(39);
output(5, 218) <= input(40);
output(5, 219) <= input(41);
output(5, 220) <= input(42);
output(5, 221) <= input(43);
output(5, 222) <= input(44);
output(5, 223) <= input(45);
output(5, 224) <= input(0);
output(5, 225) <= input(1);
output(5, 226) <= input(2);
output(5, 227) <= input(3);
output(5, 228) <= input(4);
output(5, 229) <= input(5);
output(5, 230) <= input(6);
output(5, 231) <= input(7);
output(5, 232) <= input(8);
output(5, 233) <= input(9);
output(5, 234) <= input(10);
output(5, 235) <= input(11);
output(5, 236) <= input(12);
output(5, 237) <= input(13);
output(5, 238) <= input(14);
output(5, 239) <= input(15);
output(5, 240) <= input(1);
output(5, 241) <= input(2);
output(5, 242) <= input(3);
output(5, 243) <= input(4);
output(5, 244) <= input(5);
output(5, 245) <= input(6);
output(5, 246) <= input(7);
output(5, 247) <= input(8);
output(5, 248) <= input(9);
output(5, 249) <= input(10);
output(5, 250) <= input(11);
output(5, 251) <= input(12);
output(5, 252) <= input(13);
output(5, 253) <= input(14);
output(5, 254) <= input(15);
output(5, 255) <= input(16);
when "0001" =>
output(0, 0) <= input(0);
output(0, 1) <= input(1);
output(0, 2) <= input(2);
output(0, 3) <= input(3);
output(0, 4) <= input(4);
output(0, 5) <= input(5);
output(0, 6) <= input(6);
output(0, 7) <= input(7);
output(0, 8) <= input(8);
output(0, 9) <= input(9);
output(0, 10) <= input(10);
output(0, 11) <= input(11);
output(0, 12) <= input(12);
output(0, 13) <= input(13);
output(0, 14) <= input(14);
output(0, 15) <= input(15);
output(0, 16) <= input(16);
output(0, 17) <= input(17);
output(0, 18) <= input(18);
output(0, 19) <= input(19);
output(0, 20) <= input(20);
output(0, 21) <= input(21);
output(0, 22) <= input(22);
output(0, 23) <= input(23);
output(0, 24) <= input(24);
output(0, 25) <= input(25);
output(0, 26) <= input(26);
output(0, 27) <= input(27);
output(0, 28) <= input(28);
output(0, 29) <= input(29);
output(0, 30) <= input(30);
output(0, 31) <= input(31);
output(0, 32) <= input(1);
output(0, 33) <= input(2);
output(0, 34) <= input(3);
output(0, 35) <= input(4);
output(0, 36) <= input(5);
output(0, 37) <= input(6);
output(0, 38) <= input(7);
output(0, 39) <= input(8);
output(0, 40) <= input(9);
output(0, 41) <= input(10);
output(0, 42) <= input(11);
output(0, 43) <= input(12);
output(0, 44) <= input(13);
output(0, 45) <= input(14);
output(0, 46) <= input(15);
output(0, 47) <= input(32);
output(0, 48) <= input(17);
output(0, 49) <= input(18);
output(0, 50) <= input(19);
output(0, 51) <= input(20);
output(0, 52) <= input(21);
output(0, 53) <= input(22);
output(0, 54) <= input(23);
output(0, 55) <= input(24);
output(0, 56) <= input(25);
output(0, 57) <= input(26);
output(0, 58) <= input(27);
output(0, 59) <= input(28);
output(0, 60) <= input(29);
output(0, 61) <= input(30);
output(0, 62) <= input(31);
output(0, 63) <= input(33);
output(0, 64) <= input(2);
output(0, 65) <= input(3);
output(0, 66) <= input(4);
output(0, 67) <= input(5);
output(0, 68) <= input(6);
output(0, 69) <= input(7);
output(0, 70) <= input(8);
output(0, 71) <= input(9);
output(0, 72) <= input(10);
output(0, 73) <= input(11);
output(0, 74) <= input(12);
output(0, 75) <= input(13);
output(0, 76) <= input(14);
output(0, 77) <= input(15);
output(0, 78) <= input(32);
output(0, 79) <= input(34);
output(0, 80) <= input(18);
output(0, 81) <= input(19);
output(0, 82) <= input(20);
output(0, 83) <= input(21);
output(0, 84) <= input(22);
output(0, 85) <= input(23);
output(0, 86) <= input(24);
output(0, 87) <= input(25);
output(0, 88) <= input(26);
output(0, 89) <= input(27);
output(0, 90) <= input(28);
output(0, 91) <= input(29);
output(0, 92) <= input(30);
output(0, 93) <= input(31);
output(0, 94) <= input(33);
output(0, 95) <= input(35);
output(0, 96) <= input(3);
output(0, 97) <= input(4);
output(0, 98) <= input(5);
output(0, 99) <= input(6);
output(0, 100) <= input(7);
output(0, 101) <= input(8);
output(0, 102) <= input(9);
output(0, 103) <= input(10);
output(0, 104) <= input(11);
output(0, 105) <= input(12);
output(0, 106) <= input(13);
output(0, 107) <= input(14);
output(0, 108) <= input(15);
output(0, 109) <= input(32);
output(0, 110) <= input(34);
output(0, 111) <= input(36);
output(0, 112) <= input(19);
output(0, 113) <= input(20);
output(0, 114) <= input(21);
output(0, 115) <= input(22);
output(0, 116) <= input(23);
output(0, 117) <= input(24);
output(0, 118) <= input(25);
output(0, 119) <= input(26);
output(0, 120) <= input(27);
output(0, 121) <= input(28);
output(0, 122) <= input(29);
output(0, 123) <= input(30);
output(0, 124) <= input(31);
output(0, 125) <= input(33);
output(0, 126) <= input(35);
output(0, 127) <= input(37);
output(0, 128) <= input(4);
output(0, 129) <= input(5);
output(0, 130) <= input(6);
output(0, 131) <= input(7);
output(0, 132) <= input(8);
output(0, 133) <= input(9);
output(0, 134) <= input(10);
output(0, 135) <= input(11);
output(0, 136) <= input(12);
output(0, 137) <= input(13);
output(0, 138) <= input(14);
output(0, 139) <= input(15);
output(0, 140) <= input(32);
output(0, 141) <= input(34);
output(0, 142) <= input(36);
output(0, 143) <= input(38);
output(0, 144) <= input(20);
output(0, 145) <= input(21);
output(0, 146) <= input(22);
output(0, 147) <= input(23);
output(0, 148) <= input(24);
output(0, 149) <= input(25);
output(0, 150) <= input(26);
output(0, 151) <= input(27);
output(0, 152) <= input(28);
output(0, 153) <= input(29);
output(0, 154) <= input(30);
output(0, 155) <= input(31);
output(0, 156) <= input(33);
output(0, 157) <= input(35);
output(0, 158) <= input(37);
output(0, 159) <= input(39);
output(0, 160) <= input(5);
output(0, 161) <= input(6);
output(0, 162) <= input(7);
output(0, 163) <= input(8);
output(0, 164) <= input(9);
output(0, 165) <= input(10);
output(0, 166) <= input(11);
output(0, 167) <= input(12);
output(0, 168) <= input(13);
output(0, 169) <= input(14);
output(0, 170) <= input(15);
output(0, 171) <= input(32);
output(0, 172) <= input(34);
output(0, 173) <= input(36);
output(0, 174) <= input(38);
output(0, 175) <= input(40);
output(0, 176) <= input(21);
output(0, 177) <= input(22);
output(0, 178) <= input(23);
output(0, 179) <= input(24);
output(0, 180) <= input(25);
output(0, 181) <= input(26);
output(0, 182) <= input(27);
output(0, 183) <= input(28);
output(0, 184) <= input(29);
output(0, 185) <= input(30);
output(0, 186) <= input(31);
output(0, 187) <= input(33);
output(0, 188) <= input(35);
output(0, 189) <= input(37);
output(0, 190) <= input(39);
output(0, 191) <= input(41);
output(0, 192) <= input(6);
output(0, 193) <= input(7);
output(0, 194) <= input(8);
output(0, 195) <= input(9);
output(0, 196) <= input(10);
output(0, 197) <= input(11);
output(0, 198) <= input(12);
output(0, 199) <= input(13);
output(0, 200) <= input(14);
output(0, 201) <= input(15);
output(0, 202) <= input(32);
output(0, 203) <= input(34);
output(0, 204) <= input(36);
output(0, 205) <= input(38);
output(0, 206) <= input(40);
output(0, 207) <= input(42);
output(0, 208) <= input(22);
output(0, 209) <= input(23);
output(0, 210) <= input(24);
output(0, 211) <= input(25);
output(0, 212) <= input(26);
output(0, 213) <= input(27);
output(0, 214) <= input(28);
output(0, 215) <= input(29);
output(0, 216) <= input(30);
output(0, 217) <= input(31);
output(0, 218) <= input(33);
output(0, 219) <= input(35);
output(0, 220) <= input(37);
output(0, 221) <= input(39);
output(0, 222) <= input(41);
output(0, 223) <= input(43);
output(0, 224) <= input(7);
output(0, 225) <= input(8);
output(0, 226) <= input(9);
output(0, 227) <= input(10);
output(0, 228) <= input(11);
output(0, 229) <= input(12);
output(0, 230) <= input(13);
output(0, 231) <= input(14);
output(0, 232) <= input(15);
output(0, 233) <= input(32);
output(0, 234) <= input(34);
output(0, 235) <= input(36);
output(0, 236) <= input(38);
output(0, 237) <= input(40);
output(0, 238) <= input(42);
output(0, 239) <= input(44);
output(0, 240) <= input(23);
output(0, 241) <= input(24);
output(0, 242) <= input(25);
output(0, 243) <= input(26);
output(0, 244) <= input(27);
output(0, 245) <= input(28);
output(0, 246) <= input(29);
output(0, 247) <= input(30);
output(0, 248) <= input(31);
output(0, 249) <= input(33);
output(0, 250) <= input(35);
output(0, 251) <= input(37);
output(0, 252) <= input(39);
output(0, 253) <= input(41);
output(0, 254) <= input(43);
output(0, 255) <= input(45);
output(1, 0) <= input(46);
output(1, 1) <= input(47);
output(1, 2) <= input(16);
output(1, 3) <= input(17);
output(1, 4) <= input(18);
output(1, 5) <= input(19);
output(1, 6) <= input(20);
output(1, 7) <= input(21);
output(1, 8) <= input(22);
output(1, 9) <= input(23);
output(1, 10) <= input(24);
output(1, 11) <= input(25);
output(1, 12) <= input(26);
output(1, 13) <= input(27);
output(1, 14) <= input(28);
output(1, 15) <= input(29);
output(1, 16) <= input(48);
output(1, 17) <= input(0);
output(1, 18) <= input(1);
output(1, 19) <= input(2);
output(1, 20) <= input(3);
output(1, 21) <= input(4);
output(1, 22) <= input(5);
output(1, 23) <= input(6);
output(1, 24) <= input(7);
output(1, 25) <= input(8);
output(1, 26) <= input(9);
output(1, 27) <= input(10);
output(1, 28) <= input(11);
output(1, 29) <= input(12);
output(1, 30) <= input(13);
output(1, 31) <= input(14);
output(1, 32) <= input(47);
output(1, 33) <= input(16);
output(1, 34) <= input(17);
output(1, 35) <= input(18);
output(1, 36) <= input(19);
output(1, 37) <= input(20);
output(1, 38) <= input(21);
output(1, 39) <= input(22);
output(1, 40) <= input(23);
output(1, 41) <= input(24);
output(1, 42) <= input(25);
output(1, 43) <= input(26);
output(1, 44) <= input(27);
output(1, 45) <= input(28);
output(1, 46) <= input(29);
output(1, 47) <= input(30);
output(1, 48) <= input(0);
output(1, 49) <= input(1);
output(1, 50) <= input(2);
output(1, 51) <= input(3);
output(1, 52) <= input(4);
output(1, 53) <= input(5);
output(1, 54) <= input(6);
output(1, 55) <= input(7);
output(1, 56) <= input(8);
output(1, 57) <= input(9);
output(1, 58) <= input(10);
output(1, 59) <= input(11);
output(1, 60) <= input(12);
output(1, 61) <= input(13);
output(1, 62) <= input(14);
output(1, 63) <= input(15);
output(1, 64) <= input(16);
output(1, 65) <= input(17);
output(1, 66) <= input(18);
output(1, 67) <= input(19);
output(1, 68) <= input(20);
output(1, 69) <= input(21);
output(1, 70) <= input(22);
output(1, 71) <= input(23);
output(1, 72) <= input(24);
output(1, 73) <= input(25);
output(1, 74) <= input(26);
output(1, 75) <= input(27);
output(1, 76) <= input(28);
output(1, 77) <= input(29);
output(1, 78) <= input(30);
output(1, 79) <= input(31);
output(1, 80) <= input(1);
output(1, 81) <= input(2);
output(1, 82) <= input(3);
output(1, 83) <= input(4);
output(1, 84) <= input(5);
output(1, 85) <= input(6);
output(1, 86) <= input(7);
output(1, 87) <= input(8);
output(1, 88) <= input(9);
output(1, 89) <= input(10);
output(1, 90) <= input(11);
output(1, 91) <= input(12);
output(1, 92) <= input(13);
output(1, 93) <= input(14);
output(1, 94) <= input(15);
output(1, 95) <= input(32);
output(1, 96) <= input(17);
output(1, 97) <= input(18);
output(1, 98) <= input(19);
output(1, 99) <= input(20);
output(1, 100) <= input(21);
output(1, 101) <= input(22);
output(1, 102) <= input(23);
output(1, 103) <= input(24);
output(1, 104) <= input(25);
output(1, 105) <= input(26);
output(1, 106) <= input(27);
output(1, 107) <= input(28);
output(1, 108) <= input(29);
output(1, 109) <= input(30);
output(1, 110) <= input(31);
output(1, 111) <= input(33);
output(1, 112) <= input(2);
output(1, 113) <= input(3);
output(1, 114) <= input(4);
output(1, 115) <= input(5);
output(1, 116) <= input(6);
output(1, 117) <= input(7);
output(1, 118) <= input(8);
output(1, 119) <= input(9);
output(1, 120) <= input(10);
output(1, 121) <= input(11);
output(1, 122) <= input(12);
output(1, 123) <= input(13);
output(1, 124) <= input(14);
output(1, 125) <= input(15);
output(1, 126) <= input(32);
output(1, 127) <= input(34);
output(1, 128) <= input(2);
output(1, 129) <= input(3);
output(1, 130) <= input(4);
output(1, 131) <= input(5);
output(1, 132) <= input(6);
output(1, 133) <= input(7);
output(1, 134) <= input(8);
output(1, 135) <= input(9);
output(1, 136) <= input(10);
output(1, 137) <= input(11);
output(1, 138) <= input(12);
output(1, 139) <= input(13);
output(1, 140) <= input(14);
output(1, 141) <= input(15);
output(1, 142) <= input(32);
output(1, 143) <= input(34);
output(1, 144) <= input(18);
output(1, 145) <= input(19);
output(1, 146) <= input(20);
output(1, 147) <= input(21);
output(1, 148) <= input(22);
output(1, 149) <= input(23);
output(1, 150) <= input(24);
output(1, 151) <= input(25);
output(1, 152) <= input(26);
output(1, 153) <= input(27);
output(1, 154) <= input(28);
output(1, 155) <= input(29);
output(1, 156) <= input(30);
output(1, 157) <= input(31);
output(1, 158) <= input(33);
output(1, 159) <= input(35);
output(1, 160) <= input(3);
output(1, 161) <= input(4);
output(1, 162) <= input(5);
output(1, 163) <= input(6);
output(1, 164) <= input(7);
output(1, 165) <= input(8);
output(1, 166) <= input(9);
output(1, 167) <= input(10);
output(1, 168) <= input(11);
output(1, 169) <= input(12);
output(1, 170) <= input(13);
output(1, 171) <= input(14);
output(1, 172) <= input(15);
output(1, 173) <= input(32);
output(1, 174) <= input(34);
output(1, 175) <= input(36);
output(1, 176) <= input(19);
output(1, 177) <= input(20);
output(1, 178) <= input(21);
output(1, 179) <= input(22);
output(1, 180) <= input(23);
output(1, 181) <= input(24);
output(1, 182) <= input(25);
output(1, 183) <= input(26);
output(1, 184) <= input(27);
output(1, 185) <= input(28);
output(1, 186) <= input(29);
output(1, 187) <= input(30);
output(1, 188) <= input(31);
output(1, 189) <= input(33);
output(1, 190) <= input(35);
output(1, 191) <= input(37);
output(1, 192) <= input(4);
output(1, 193) <= input(5);
output(1, 194) <= input(6);
output(1, 195) <= input(7);
output(1, 196) <= input(8);
output(1, 197) <= input(9);
output(1, 198) <= input(10);
output(1, 199) <= input(11);
output(1, 200) <= input(12);
output(1, 201) <= input(13);
output(1, 202) <= input(14);
output(1, 203) <= input(15);
output(1, 204) <= input(32);
output(1, 205) <= input(34);
output(1, 206) <= input(36);
output(1, 207) <= input(38);
output(1, 208) <= input(20);
output(1, 209) <= input(21);
output(1, 210) <= input(22);
output(1, 211) <= input(23);
output(1, 212) <= input(24);
output(1, 213) <= input(25);
output(1, 214) <= input(26);
output(1, 215) <= input(27);
output(1, 216) <= input(28);
output(1, 217) <= input(29);
output(1, 218) <= input(30);
output(1, 219) <= input(31);
output(1, 220) <= input(33);
output(1, 221) <= input(35);
output(1, 222) <= input(37);
output(1, 223) <= input(39);
output(1, 224) <= input(5);
output(1, 225) <= input(6);
output(1, 226) <= input(7);
output(1, 227) <= input(8);
output(1, 228) <= input(9);
output(1, 229) <= input(10);
output(1, 230) <= input(11);
output(1, 231) <= input(12);
output(1, 232) <= input(13);
output(1, 233) <= input(14);
output(1, 234) <= input(15);
output(1, 235) <= input(32);
output(1, 236) <= input(34);
output(1, 237) <= input(36);
output(1, 238) <= input(38);
output(1, 239) <= input(40);
output(1, 240) <= input(21);
output(1, 241) <= input(22);
output(1, 242) <= input(23);
output(1, 243) <= input(24);
output(1, 244) <= input(25);
output(1, 245) <= input(26);
output(1, 246) <= input(27);
output(1, 247) <= input(28);
output(1, 248) <= input(29);
output(1, 249) <= input(30);
output(1, 250) <= input(31);
output(1, 251) <= input(33);
output(1, 252) <= input(35);
output(1, 253) <= input(37);
output(1, 254) <= input(39);
output(1, 255) <= input(41);
output(2, 0) <= input(49);
output(2, 1) <= input(46);
output(2, 2) <= input(47);
output(2, 3) <= input(16);
output(2, 4) <= input(17);
output(2, 5) <= input(18);
output(2, 6) <= input(19);
output(2, 7) <= input(20);
output(2, 8) <= input(21);
output(2, 9) <= input(22);
output(2, 10) <= input(23);
output(2, 11) <= input(24);
output(2, 12) <= input(25);
output(2, 13) <= input(26);
output(2, 14) <= input(27);
output(2, 15) <= input(28);
output(2, 16) <= input(50);
output(2, 17) <= input(48);
output(2, 18) <= input(0);
output(2, 19) <= input(1);
output(2, 20) <= input(2);
output(2, 21) <= input(3);
output(2, 22) <= input(4);
output(2, 23) <= input(5);
output(2, 24) <= input(6);
output(2, 25) <= input(7);
output(2, 26) <= input(8);
output(2, 27) <= input(9);
output(2, 28) <= input(10);
output(2, 29) <= input(11);
output(2, 30) <= input(12);
output(2, 31) <= input(13);
output(2, 32) <= input(46);
output(2, 33) <= input(47);
output(2, 34) <= input(16);
output(2, 35) <= input(17);
output(2, 36) <= input(18);
output(2, 37) <= input(19);
output(2, 38) <= input(20);
output(2, 39) <= input(21);
output(2, 40) <= input(22);
output(2, 41) <= input(23);
output(2, 42) <= input(24);
output(2, 43) <= input(25);
output(2, 44) <= input(26);
output(2, 45) <= input(27);
output(2, 46) <= input(28);
output(2, 47) <= input(29);
output(2, 48) <= input(48);
output(2, 49) <= input(0);
output(2, 50) <= input(1);
output(2, 51) <= input(2);
output(2, 52) <= input(3);
output(2, 53) <= input(4);
output(2, 54) <= input(5);
output(2, 55) <= input(6);
output(2, 56) <= input(7);
output(2, 57) <= input(8);
output(2, 58) <= input(9);
output(2, 59) <= input(10);
output(2, 60) <= input(11);
output(2, 61) <= input(12);
output(2, 62) <= input(13);
output(2, 63) <= input(14);
output(2, 64) <= input(48);
output(2, 65) <= input(0);
output(2, 66) <= input(1);
output(2, 67) <= input(2);
output(2, 68) <= input(3);
output(2, 69) <= input(4);
output(2, 70) <= input(5);
output(2, 71) <= input(6);
output(2, 72) <= input(7);
output(2, 73) <= input(8);
output(2, 74) <= input(9);
output(2, 75) <= input(10);
output(2, 76) <= input(11);
output(2, 77) <= input(12);
output(2, 78) <= input(13);
output(2, 79) <= input(14);
output(2, 80) <= input(47);
output(2, 81) <= input(16);
output(2, 82) <= input(17);
output(2, 83) <= input(18);
output(2, 84) <= input(19);
output(2, 85) <= input(20);
output(2, 86) <= input(21);
output(2, 87) <= input(22);
output(2, 88) <= input(23);
output(2, 89) <= input(24);
output(2, 90) <= input(25);
output(2, 91) <= input(26);
output(2, 92) <= input(27);
output(2, 93) <= input(28);
output(2, 94) <= input(29);
output(2, 95) <= input(30);
output(2, 96) <= input(0);
output(2, 97) <= input(1);
output(2, 98) <= input(2);
output(2, 99) <= input(3);
output(2, 100) <= input(4);
output(2, 101) <= input(5);
output(2, 102) <= input(6);
output(2, 103) <= input(7);
output(2, 104) <= input(8);
output(2, 105) <= input(9);
output(2, 106) <= input(10);
output(2, 107) <= input(11);
output(2, 108) <= input(12);
output(2, 109) <= input(13);
output(2, 110) <= input(14);
output(2, 111) <= input(15);
output(2, 112) <= input(16);
output(2, 113) <= input(17);
output(2, 114) <= input(18);
output(2, 115) <= input(19);
output(2, 116) <= input(20);
output(2, 117) <= input(21);
output(2, 118) <= input(22);
output(2, 119) <= input(23);
output(2, 120) <= input(24);
output(2, 121) <= input(25);
output(2, 122) <= input(26);
output(2, 123) <= input(27);
output(2, 124) <= input(28);
output(2, 125) <= input(29);
output(2, 126) <= input(30);
output(2, 127) <= input(31);
output(2, 128) <= input(16);
output(2, 129) <= input(17);
output(2, 130) <= input(18);
output(2, 131) <= input(19);
output(2, 132) <= input(20);
output(2, 133) <= input(21);
output(2, 134) <= input(22);
output(2, 135) <= input(23);
output(2, 136) <= input(24);
output(2, 137) <= input(25);
output(2, 138) <= input(26);
output(2, 139) <= input(27);
output(2, 140) <= input(28);
output(2, 141) <= input(29);
output(2, 142) <= input(30);
output(2, 143) <= input(31);
output(2, 144) <= input(1);
output(2, 145) <= input(2);
output(2, 146) <= input(3);
output(2, 147) <= input(4);
output(2, 148) <= input(5);
output(2, 149) <= input(6);
output(2, 150) <= input(7);
output(2, 151) <= input(8);
output(2, 152) <= input(9);
output(2, 153) <= input(10);
output(2, 154) <= input(11);
output(2, 155) <= input(12);
output(2, 156) <= input(13);
output(2, 157) <= input(14);
output(2, 158) <= input(15);
output(2, 159) <= input(32);
output(2, 160) <= input(17);
output(2, 161) <= input(18);
output(2, 162) <= input(19);
output(2, 163) <= input(20);
output(2, 164) <= input(21);
output(2, 165) <= input(22);
output(2, 166) <= input(23);
output(2, 167) <= input(24);
output(2, 168) <= input(25);
output(2, 169) <= input(26);
output(2, 170) <= input(27);
output(2, 171) <= input(28);
output(2, 172) <= input(29);
output(2, 173) <= input(30);
output(2, 174) <= input(31);
output(2, 175) <= input(33);
output(2, 176) <= input(2);
output(2, 177) <= input(3);
output(2, 178) <= input(4);
output(2, 179) <= input(5);
output(2, 180) <= input(6);
output(2, 181) <= input(7);
output(2, 182) <= input(8);
output(2, 183) <= input(9);
output(2, 184) <= input(10);
output(2, 185) <= input(11);
output(2, 186) <= input(12);
output(2, 187) <= input(13);
output(2, 188) <= input(14);
output(2, 189) <= input(15);
output(2, 190) <= input(32);
output(2, 191) <= input(34);
output(2, 192) <= input(2);
output(2, 193) <= input(3);
output(2, 194) <= input(4);
output(2, 195) <= input(5);
output(2, 196) <= input(6);
output(2, 197) <= input(7);
output(2, 198) <= input(8);
output(2, 199) <= input(9);
output(2, 200) <= input(10);
output(2, 201) <= input(11);
output(2, 202) <= input(12);
output(2, 203) <= input(13);
output(2, 204) <= input(14);
output(2, 205) <= input(15);
output(2, 206) <= input(32);
output(2, 207) <= input(34);
output(2, 208) <= input(18);
output(2, 209) <= input(19);
output(2, 210) <= input(20);
output(2, 211) <= input(21);
output(2, 212) <= input(22);
output(2, 213) <= input(23);
output(2, 214) <= input(24);
output(2, 215) <= input(25);
output(2, 216) <= input(26);
output(2, 217) <= input(27);
output(2, 218) <= input(28);
output(2, 219) <= input(29);
output(2, 220) <= input(30);
output(2, 221) <= input(31);
output(2, 222) <= input(33);
output(2, 223) <= input(35);
output(2, 224) <= input(3);
output(2, 225) <= input(4);
output(2, 226) <= input(5);
output(2, 227) <= input(6);
output(2, 228) <= input(7);
output(2, 229) <= input(8);
output(2, 230) <= input(9);
output(2, 231) <= input(10);
output(2, 232) <= input(11);
output(2, 233) <= input(12);
output(2, 234) <= input(13);
output(2, 235) <= input(14);
output(2, 236) <= input(15);
output(2, 237) <= input(32);
output(2, 238) <= input(34);
output(2, 239) <= input(36);
output(2, 240) <= input(19);
output(2, 241) <= input(20);
output(2, 242) <= input(21);
output(2, 243) <= input(22);
output(2, 244) <= input(23);
output(2, 245) <= input(24);
output(2, 246) <= input(25);
output(2, 247) <= input(26);
output(2, 248) <= input(27);
output(2, 249) <= input(28);
output(2, 250) <= input(29);
output(2, 251) <= input(30);
output(2, 252) <= input(31);
output(2, 253) <= input(33);
output(2, 254) <= input(35);
output(2, 255) <= input(37);
output(3, 0) <= input(51);
output(3, 1) <= input(49);
output(3, 2) <= input(46);
output(3, 3) <= input(47);
output(3, 4) <= input(16);
output(3, 5) <= input(17);
output(3, 6) <= input(18);
output(3, 7) <= input(19);
output(3, 8) <= input(20);
output(3, 9) <= input(21);
output(3, 10) <= input(22);
output(3, 11) <= input(23);
output(3, 12) <= input(24);
output(3, 13) <= input(25);
output(3, 14) <= input(26);
output(3, 15) <= input(27);
output(3, 16) <= input(52);
output(3, 17) <= input(50);
output(3, 18) <= input(48);
output(3, 19) <= input(0);
output(3, 20) <= input(1);
output(3, 21) <= input(2);
output(3, 22) <= input(3);
output(3, 23) <= input(4);
output(3, 24) <= input(5);
output(3, 25) <= input(6);
output(3, 26) <= input(7);
output(3, 27) <= input(8);
output(3, 28) <= input(9);
output(3, 29) <= input(10);
output(3, 30) <= input(11);
output(3, 31) <= input(12);
output(3, 32) <= input(52);
output(3, 33) <= input(50);
output(3, 34) <= input(48);
output(3, 35) <= input(0);
output(3, 36) <= input(1);
output(3, 37) <= input(2);
output(3, 38) <= input(3);
output(3, 39) <= input(4);
output(3, 40) <= input(5);
output(3, 41) <= input(6);
output(3, 42) <= input(7);
output(3, 43) <= input(8);
output(3, 44) <= input(9);
output(3, 45) <= input(10);
output(3, 46) <= input(11);
output(3, 47) <= input(12);
output(3, 48) <= input(49);
output(3, 49) <= input(46);
output(3, 50) <= input(47);
output(3, 51) <= input(16);
output(3, 52) <= input(17);
output(3, 53) <= input(18);
output(3, 54) <= input(19);
output(3, 55) <= input(20);
output(3, 56) <= input(21);
output(3, 57) <= input(22);
output(3, 58) <= input(23);
output(3, 59) <= input(24);
output(3, 60) <= input(25);
output(3, 61) <= input(26);
output(3, 62) <= input(27);
output(3, 63) <= input(28);
output(3, 64) <= input(50);
output(3, 65) <= input(48);
output(3, 66) <= input(0);
output(3, 67) <= input(1);
output(3, 68) <= input(2);
output(3, 69) <= input(3);
output(3, 70) <= input(4);
output(3, 71) <= input(5);
output(3, 72) <= input(6);
output(3, 73) <= input(7);
output(3, 74) <= input(8);
output(3, 75) <= input(9);
output(3, 76) <= input(10);
output(3, 77) <= input(11);
output(3, 78) <= input(12);
output(3, 79) <= input(13);
output(3, 80) <= input(50);
output(3, 81) <= input(48);
output(3, 82) <= input(0);
output(3, 83) <= input(1);
output(3, 84) <= input(2);
output(3, 85) <= input(3);
output(3, 86) <= input(4);
output(3, 87) <= input(5);
output(3, 88) <= input(6);
output(3, 89) <= input(7);
output(3, 90) <= input(8);
output(3, 91) <= input(9);
output(3, 92) <= input(10);
output(3, 93) <= input(11);
output(3, 94) <= input(12);
output(3, 95) <= input(13);
output(3, 96) <= input(46);
output(3, 97) <= input(47);
output(3, 98) <= input(16);
output(3, 99) <= input(17);
output(3, 100) <= input(18);
output(3, 101) <= input(19);
output(3, 102) <= input(20);
output(3, 103) <= input(21);
output(3, 104) <= input(22);
output(3, 105) <= input(23);
output(3, 106) <= input(24);
output(3, 107) <= input(25);
output(3, 108) <= input(26);
output(3, 109) <= input(27);
output(3, 110) <= input(28);
output(3, 111) <= input(29);
output(3, 112) <= input(48);
output(3, 113) <= input(0);
output(3, 114) <= input(1);
output(3, 115) <= input(2);
output(3, 116) <= input(3);
output(3, 117) <= input(4);
output(3, 118) <= input(5);
output(3, 119) <= input(6);
output(3, 120) <= input(7);
output(3, 121) <= input(8);
output(3, 122) <= input(9);
output(3, 123) <= input(10);
output(3, 124) <= input(11);
output(3, 125) <= input(12);
output(3, 126) <= input(13);
output(3, 127) <= input(14);
output(3, 128) <= input(48);
output(3, 129) <= input(0);
output(3, 130) <= input(1);
output(3, 131) <= input(2);
output(3, 132) <= input(3);
output(3, 133) <= input(4);
output(3, 134) <= input(5);
output(3, 135) <= input(6);
output(3, 136) <= input(7);
output(3, 137) <= input(8);
output(3, 138) <= input(9);
output(3, 139) <= input(10);
output(3, 140) <= input(11);
output(3, 141) <= input(12);
output(3, 142) <= input(13);
output(3, 143) <= input(14);
output(3, 144) <= input(47);
output(3, 145) <= input(16);
output(3, 146) <= input(17);
output(3, 147) <= input(18);
output(3, 148) <= input(19);
output(3, 149) <= input(20);
output(3, 150) <= input(21);
output(3, 151) <= input(22);
output(3, 152) <= input(23);
output(3, 153) <= input(24);
output(3, 154) <= input(25);
output(3, 155) <= input(26);
output(3, 156) <= input(27);
output(3, 157) <= input(28);
output(3, 158) <= input(29);
output(3, 159) <= input(30);
output(3, 160) <= input(47);
output(3, 161) <= input(16);
output(3, 162) <= input(17);
output(3, 163) <= input(18);
output(3, 164) <= input(19);
output(3, 165) <= input(20);
output(3, 166) <= input(21);
output(3, 167) <= input(22);
output(3, 168) <= input(23);
output(3, 169) <= input(24);
output(3, 170) <= input(25);
output(3, 171) <= input(26);
output(3, 172) <= input(27);
output(3, 173) <= input(28);
output(3, 174) <= input(29);
output(3, 175) <= input(30);
output(3, 176) <= input(0);
output(3, 177) <= input(1);
output(3, 178) <= input(2);
output(3, 179) <= input(3);
output(3, 180) <= input(4);
output(3, 181) <= input(5);
output(3, 182) <= input(6);
output(3, 183) <= input(7);
output(3, 184) <= input(8);
output(3, 185) <= input(9);
output(3, 186) <= input(10);
output(3, 187) <= input(11);
output(3, 188) <= input(12);
output(3, 189) <= input(13);
output(3, 190) <= input(14);
output(3, 191) <= input(15);
output(3, 192) <= input(16);
output(3, 193) <= input(17);
output(3, 194) <= input(18);
output(3, 195) <= input(19);
output(3, 196) <= input(20);
output(3, 197) <= input(21);
output(3, 198) <= input(22);
output(3, 199) <= input(23);
output(3, 200) <= input(24);
output(3, 201) <= input(25);
output(3, 202) <= input(26);
output(3, 203) <= input(27);
output(3, 204) <= input(28);
output(3, 205) <= input(29);
output(3, 206) <= input(30);
output(3, 207) <= input(31);
output(3, 208) <= input(16);
output(3, 209) <= input(17);
output(3, 210) <= input(18);
output(3, 211) <= input(19);
output(3, 212) <= input(20);
output(3, 213) <= input(21);
output(3, 214) <= input(22);
output(3, 215) <= input(23);
output(3, 216) <= input(24);
output(3, 217) <= input(25);
output(3, 218) <= input(26);
output(3, 219) <= input(27);
output(3, 220) <= input(28);
output(3, 221) <= input(29);
output(3, 222) <= input(30);
output(3, 223) <= input(31);
output(3, 224) <= input(1);
output(3, 225) <= input(2);
output(3, 226) <= input(3);
output(3, 227) <= input(4);
output(3, 228) <= input(5);
output(3, 229) <= input(6);
output(3, 230) <= input(7);
output(3, 231) <= input(8);
output(3, 232) <= input(9);
output(3, 233) <= input(10);
output(3, 234) <= input(11);
output(3, 235) <= input(12);
output(3, 236) <= input(13);
output(3, 237) <= input(14);
output(3, 238) <= input(15);
output(3, 239) <= input(32);
output(3, 240) <= input(17);
output(3, 241) <= input(18);
output(3, 242) <= input(19);
output(3, 243) <= input(20);
output(3, 244) <= input(21);
output(3, 245) <= input(22);
output(3, 246) <= input(23);
output(3, 247) <= input(24);
output(3, 248) <= input(25);
output(3, 249) <= input(26);
output(3, 250) <= input(27);
output(3, 251) <= input(28);
output(3, 252) <= input(29);
output(3, 253) <= input(30);
output(3, 254) <= input(31);
output(3, 255) <= input(33);
output(4, 0) <= input(53);
output(4, 1) <= input(51);
output(4, 2) <= input(49);
output(4, 3) <= input(46);
output(4, 4) <= input(47);
output(4, 5) <= input(16);
output(4, 6) <= input(17);
output(4, 7) <= input(18);
output(4, 8) <= input(19);
output(4, 9) <= input(20);
output(4, 10) <= input(21);
output(4, 11) <= input(22);
output(4, 12) <= input(23);
output(4, 13) <= input(24);
output(4, 14) <= input(25);
output(4, 15) <= input(26);
output(4, 16) <= input(54);
output(4, 17) <= input(52);
output(4, 18) <= input(50);
output(4, 19) <= input(48);
output(4, 20) <= input(0);
output(4, 21) <= input(1);
output(4, 22) <= input(2);
output(4, 23) <= input(3);
output(4, 24) <= input(4);
output(4, 25) <= input(5);
output(4, 26) <= input(6);
output(4, 27) <= input(7);
output(4, 28) <= input(8);
output(4, 29) <= input(9);
output(4, 30) <= input(10);
output(4, 31) <= input(11);
output(4, 32) <= input(54);
output(4, 33) <= input(52);
output(4, 34) <= input(50);
output(4, 35) <= input(48);
output(4, 36) <= input(0);
output(4, 37) <= input(1);
output(4, 38) <= input(2);
output(4, 39) <= input(3);
output(4, 40) <= input(4);
output(4, 41) <= input(5);
output(4, 42) <= input(6);
output(4, 43) <= input(7);
output(4, 44) <= input(8);
output(4, 45) <= input(9);
output(4, 46) <= input(10);
output(4, 47) <= input(11);
output(4, 48) <= input(51);
output(4, 49) <= input(49);
output(4, 50) <= input(46);
output(4, 51) <= input(47);
output(4, 52) <= input(16);
output(4, 53) <= input(17);
output(4, 54) <= input(18);
output(4, 55) <= input(19);
output(4, 56) <= input(20);
output(4, 57) <= input(21);
output(4, 58) <= input(22);
output(4, 59) <= input(23);
output(4, 60) <= input(24);
output(4, 61) <= input(25);
output(4, 62) <= input(26);
output(4, 63) <= input(27);
output(4, 64) <= input(51);
output(4, 65) <= input(49);
output(4, 66) <= input(46);
output(4, 67) <= input(47);
output(4, 68) <= input(16);
output(4, 69) <= input(17);
output(4, 70) <= input(18);
output(4, 71) <= input(19);
output(4, 72) <= input(20);
output(4, 73) <= input(21);
output(4, 74) <= input(22);
output(4, 75) <= input(23);
output(4, 76) <= input(24);
output(4, 77) <= input(25);
output(4, 78) <= input(26);
output(4, 79) <= input(27);
output(4, 80) <= input(52);
output(4, 81) <= input(50);
output(4, 82) <= input(48);
output(4, 83) <= input(0);
output(4, 84) <= input(1);
output(4, 85) <= input(2);
output(4, 86) <= input(3);
output(4, 87) <= input(4);
output(4, 88) <= input(5);
output(4, 89) <= input(6);
output(4, 90) <= input(7);
output(4, 91) <= input(8);
output(4, 92) <= input(9);
output(4, 93) <= input(10);
output(4, 94) <= input(11);
output(4, 95) <= input(12);
output(4, 96) <= input(52);
output(4, 97) <= input(50);
output(4, 98) <= input(48);
output(4, 99) <= input(0);
output(4, 100) <= input(1);
output(4, 101) <= input(2);
output(4, 102) <= input(3);
output(4, 103) <= input(4);
output(4, 104) <= input(5);
output(4, 105) <= input(6);
output(4, 106) <= input(7);
output(4, 107) <= input(8);
output(4, 108) <= input(9);
output(4, 109) <= input(10);
output(4, 110) <= input(11);
output(4, 111) <= input(12);
output(4, 112) <= input(49);
output(4, 113) <= input(46);
output(4, 114) <= input(47);
output(4, 115) <= input(16);
output(4, 116) <= input(17);
output(4, 117) <= input(18);
output(4, 118) <= input(19);
output(4, 119) <= input(20);
output(4, 120) <= input(21);
output(4, 121) <= input(22);
output(4, 122) <= input(23);
output(4, 123) <= input(24);
output(4, 124) <= input(25);
output(4, 125) <= input(26);
output(4, 126) <= input(27);
output(4, 127) <= input(28);
output(4, 128) <= input(49);
output(4, 129) <= input(46);
output(4, 130) <= input(47);
output(4, 131) <= input(16);
output(4, 132) <= input(17);
output(4, 133) <= input(18);
output(4, 134) <= input(19);
output(4, 135) <= input(20);
output(4, 136) <= input(21);
output(4, 137) <= input(22);
output(4, 138) <= input(23);
output(4, 139) <= input(24);
output(4, 140) <= input(25);
output(4, 141) <= input(26);
output(4, 142) <= input(27);
output(4, 143) <= input(28);
output(4, 144) <= input(50);
output(4, 145) <= input(48);
output(4, 146) <= input(0);
output(4, 147) <= input(1);
output(4, 148) <= input(2);
output(4, 149) <= input(3);
output(4, 150) <= input(4);
output(4, 151) <= input(5);
output(4, 152) <= input(6);
output(4, 153) <= input(7);
output(4, 154) <= input(8);
output(4, 155) <= input(9);
output(4, 156) <= input(10);
output(4, 157) <= input(11);
output(4, 158) <= input(12);
output(4, 159) <= input(13);
output(4, 160) <= input(50);
output(4, 161) <= input(48);
output(4, 162) <= input(0);
output(4, 163) <= input(1);
output(4, 164) <= input(2);
output(4, 165) <= input(3);
output(4, 166) <= input(4);
output(4, 167) <= input(5);
output(4, 168) <= input(6);
output(4, 169) <= input(7);
output(4, 170) <= input(8);
output(4, 171) <= input(9);
output(4, 172) <= input(10);
output(4, 173) <= input(11);
output(4, 174) <= input(12);
output(4, 175) <= input(13);
output(4, 176) <= input(46);
output(4, 177) <= input(47);
output(4, 178) <= input(16);
output(4, 179) <= input(17);
output(4, 180) <= input(18);
output(4, 181) <= input(19);
output(4, 182) <= input(20);
output(4, 183) <= input(21);
output(4, 184) <= input(22);
output(4, 185) <= input(23);
output(4, 186) <= input(24);
output(4, 187) <= input(25);
output(4, 188) <= input(26);
output(4, 189) <= input(27);
output(4, 190) <= input(28);
output(4, 191) <= input(29);
output(4, 192) <= input(46);
output(4, 193) <= input(47);
output(4, 194) <= input(16);
output(4, 195) <= input(17);
output(4, 196) <= input(18);
output(4, 197) <= input(19);
output(4, 198) <= input(20);
output(4, 199) <= input(21);
output(4, 200) <= input(22);
output(4, 201) <= input(23);
output(4, 202) <= input(24);
output(4, 203) <= input(25);
output(4, 204) <= input(26);
output(4, 205) <= input(27);
output(4, 206) <= input(28);
output(4, 207) <= input(29);
output(4, 208) <= input(48);
output(4, 209) <= input(0);
output(4, 210) <= input(1);
output(4, 211) <= input(2);
output(4, 212) <= input(3);
output(4, 213) <= input(4);
output(4, 214) <= input(5);
output(4, 215) <= input(6);
output(4, 216) <= input(7);
output(4, 217) <= input(8);
output(4, 218) <= input(9);
output(4, 219) <= input(10);
output(4, 220) <= input(11);
output(4, 221) <= input(12);
output(4, 222) <= input(13);
output(4, 223) <= input(14);
output(4, 224) <= input(48);
output(4, 225) <= input(0);
output(4, 226) <= input(1);
output(4, 227) <= input(2);
output(4, 228) <= input(3);
output(4, 229) <= input(4);
output(4, 230) <= input(5);
output(4, 231) <= input(6);
output(4, 232) <= input(7);
output(4, 233) <= input(8);
output(4, 234) <= input(9);
output(4, 235) <= input(10);
output(4, 236) <= input(11);
output(4, 237) <= input(12);
output(4, 238) <= input(13);
output(4, 239) <= input(14);
output(4, 240) <= input(47);
output(4, 241) <= input(16);
output(4, 242) <= input(17);
output(4, 243) <= input(18);
output(4, 244) <= input(19);
output(4, 245) <= input(20);
output(4, 246) <= input(21);
output(4, 247) <= input(22);
output(4, 248) <= input(23);
output(4, 249) <= input(24);
output(4, 250) <= input(25);
output(4, 251) <= input(26);
output(4, 252) <= input(27);
output(4, 253) <= input(28);
output(4, 254) <= input(29);
output(4, 255) <= input(30);
output(5, 0) <= input(55);
output(5, 1) <= input(53);
output(5, 2) <= input(51);
output(5, 3) <= input(49);
output(5, 4) <= input(46);
output(5, 5) <= input(47);
output(5, 6) <= input(16);
output(5, 7) <= input(17);
output(5, 8) <= input(18);
output(5, 9) <= input(19);
output(5, 10) <= input(20);
output(5, 11) <= input(21);
output(5, 12) <= input(22);
output(5, 13) <= input(23);
output(5, 14) <= input(24);
output(5, 15) <= input(25);
output(5, 16) <= input(55);
output(5, 17) <= input(53);
output(5, 18) <= input(51);
output(5, 19) <= input(49);
output(5, 20) <= input(46);
output(5, 21) <= input(47);
output(5, 22) <= input(16);
output(5, 23) <= input(17);
output(5, 24) <= input(18);
output(5, 25) <= input(19);
output(5, 26) <= input(20);
output(5, 27) <= input(21);
output(5, 28) <= input(22);
output(5, 29) <= input(23);
output(5, 30) <= input(24);
output(5, 31) <= input(25);
output(5, 32) <= input(56);
output(5, 33) <= input(54);
output(5, 34) <= input(52);
output(5, 35) <= input(50);
output(5, 36) <= input(48);
output(5, 37) <= input(0);
output(5, 38) <= input(1);
output(5, 39) <= input(2);
output(5, 40) <= input(3);
output(5, 41) <= input(4);
output(5, 42) <= input(5);
output(5, 43) <= input(6);
output(5, 44) <= input(7);
output(5, 45) <= input(8);
output(5, 46) <= input(9);
output(5, 47) <= input(10);
output(5, 48) <= input(56);
output(5, 49) <= input(54);
output(5, 50) <= input(52);
output(5, 51) <= input(50);
output(5, 52) <= input(48);
output(5, 53) <= input(0);
output(5, 54) <= input(1);
output(5, 55) <= input(2);
output(5, 56) <= input(3);
output(5, 57) <= input(4);
output(5, 58) <= input(5);
output(5, 59) <= input(6);
output(5, 60) <= input(7);
output(5, 61) <= input(8);
output(5, 62) <= input(9);
output(5, 63) <= input(10);
output(5, 64) <= input(56);
output(5, 65) <= input(54);
output(5, 66) <= input(52);
output(5, 67) <= input(50);
output(5, 68) <= input(48);
output(5, 69) <= input(0);
output(5, 70) <= input(1);
output(5, 71) <= input(2);
output(5, 72) <= input(3);
output(5, 73) <= input(4);
output(5, 74) <= input(5);
output(5, 75) <= input(6);
output(5, 76) <= input(7);
output(5, 77) <= input(8);
output(5, 78) <= input(9);
output(5, 79) <= input(10);
output(5, 80) <= input(53);
output(5, 81) <= input(51);
output(5, 82) <= input(49);
output(5, 83) <= input(46);
output(5, 84) <= input(47);
output(5, 85) <= input(16);
output(5, 86) <= input(17);
output(5, 87) <= input(18);
output(5, 88) <= input(19);
output(5, 89) <= input(20);
output(5, 90) <= input(21);
output(5, 91) <= input(22);
output(5, 92) <= input(23);
output(5, 93) <= input(24);
output(5, 94) <= input(25);
output(5, 95) <= input(26);
output(5, 96) <= input(53);
output(5, 97) <= input(51);
output(5, 98) <= input(49);
output(5, 99) <= input(46);
output(5, 100) <= input(47);
output(5, 101) <= input(16);
output(5, 102) <= input(17);
output(5, 103) <= input(18);
output(5, 104) <= input(19);
output(5, 105) <= input(20);
output(5, 106) <= input(21);
output(5, 107) <= input(22);
output(5, 108) <= input(23);
output(5, 109) <= input(24);
output(5, 110) <= input(25);
output(5, 111) <= input(26);
output(5, 112) <= input(54);
output(5, 113) <= input(52);
output(5, 114) <= input(50);
output(5, 115) <= input(48);
output(5, 116) <= input(0);
output(5, 117) <= input(1);
output(5, 118) <= input(2);
output(5, 119) <= input(3);
output(5, 120) <= input(4);
output(5, 121) <= input(5);
output(5, 122) <= input(6);
output(5, 123) <= input(7);
output(5, 124) <= input(8);
output(5, 125) <= input(9);
output(5, 126) <= input(10);
output(5, 127) <= input(11);
output(5, 128) <= input(54);
output(5, 129) <= input(52);
output(5, 130) <= input(50);
output(5, 131) <= input(48);
output(5, 132) <= input(0);
output(5, 133) <= input(1);
output(5, 134) <= input(2);
output(5, 135) <= input(3);
output(5, 136) <= input(4);
output(5, 137) <= input(5);
output(5, 138) <= input(6);
output(5, 139) <= input(7);
output(5, 140) <= input(8);
output(5, 141) <= input(9);
output(5, 142) <= input(10);
output(5, 143) <= input(11);
output(5, 144) <= input(54);
output(5, 145) <= input(52);
output(5, 146) <= input(50);
output(5, 147) <= input(48);
output(5, 148) <= input(0);
output(5, 149) <= input(1);
output(5, 150) <= input(2);
output(5, 151) <= input(3);
output(5, 152) <= input(4);
output(5, 153) <= input(5);
output(5, 154) <= input(6);
output(5, 155) <= input(7);
output(5, 156) <= input(8);
output(5, 157) <= input(9);
output(5, 158) <= input(10);
output(5, 159) <= input(11);
output(5, 160) <= input(51);
output(5, 161) <= input(49);
output(5, 162) <= input(46);
output(5, 163) <= input(47);
output(5, 164) <= input(16);
output(5, 165) <= input(17);
output(5, 166) <= input(18);
output(5, 167) <= input(19);
output(5, 168) <= input(20);
output(5, 169) <= input(21);
output(5, 170) <= input(22);
output(5, 171) <= input(23);
output(5, 172) <= input(24);
output(5, 173) <= input(25);
output(5, 174) <= input(26);
output(5, 175) <= input(27);
output(5, 176) <= input(51);
output(5, 177) <= input(49);
output(5, 178) <= input(46);
output(5, 179) <= input(47);
output(5, 180) <= input(16);
output(5, 181) <= input(17);
output(5, 182) <= input(18);
output(5, 183) <= input(19);
output(5, 184) <= input(20);
output(5, 185) <= input(21);
output(5, 186) <= input(22);
output(5, 187) <= input(23);
output(5, 188) <= input(24);
output(5, 189) <= input(25);
output(5, 190) <= input(26);
output(5, 191) <= input(27);
output(5, 192) <= input(51);
output(5, 193) <= input(49);
output(5, 194) <= input(46);
output(5, 195) <= input(47);
output(5, 196) <= input(16);
output(5, 197) <= input(17);
output(5, 198) <= input(18);
output(5, 199) <= input(19);
output(5, 200) <= input(20);
output(5, 201) <= input(21);
output(5, 202) <= input(22);
output(5, 203) <= input(23);
output(5, 204) <= input(24);
output(5, 205) <= input(25);
output(5, 206) <= input(26);
output(5, 207) <= input(27);
output(5, 208) <= input(52);
output(5, 209) <= input(50);
output(5, 210) <= input(48);
output(5, 211) <= input(0);
output(5, 212) <= input(1);
output(5, 213) <= input(2);
output(5, 214) <= input(3);
output(5, 215) <= input(4);
output(5, 216) <= input(5);
output(5, 217) <= input(6);
output(5, 218) <= input(7);
output(5, 219) <= input(8);
output(5, 220) <= input(9);
output(5, 221) <= input(10);
output(5, 222) <= input(11);
output(5, 223) <= input(12);
output(5, 224) <= input(52);
output(5, 225) <= input(50);
output(5, 226) <= input(48);
output(5, 227) <= input(0);
output(5, 228) <= input(1);
output(5, 229) <= input(2);
output(5, 230) <= input(3);
output(5, 231) <= input(4);
output(5, 232) <= input(5);
output(5, 233) <= input(6);
output(5, 234) <= input(7);
output(5, 235) <= input(8);
output(5, 236) <= input(9);
output(5, 237) <= input(10);
output(5, 238) <= input(11);
output(5, 239) <= input(12);
output(5, 240) <= input(49);
output(5, 241) <= input(46);
output(5, 242) <= input(47);
output(5, 243) <= input(16);
output(5, 244) <= input(17);
output(5, 245) <= input(18);
output(5, 246) <= input(19);
output(5, 247) <= input(20);
output(5, 248) <= input(21);
output(5, 249) <= input(22);
output(5, 250) <= input(23);
output(5, 251) <= input(24);
output(5, 252) <= input(25);
output(5, 253) <= input(26);
output(5, 254) <= input(27);
output(5, 255) <= input(28);
when "0010" =>
output(0, 0) <= input(0);
output(0, 1) <= input(1);
output(0, 2) <= input(2);
output(0, 3) <= input(3);
output(0, 4) <= input(4);
output(0, 5) <= input(5);
output(0, 6) <= input(6);
output(0, 7) <= input(7);
output(0, 8) <= input(8);
output(0, 9) <= input(9);
output(0, 10) <= input(10);
output(0, 11) <= input(11);
output(0, 12) <= input(12);
output(0, 13) <= input(13);
output(0, 14) <= input(14);
output(0, 15) <= input(15);
output(0, 16) <= input(0);
output(0, 17) <= input(1);
output(0, 18) <= input(2);
output(0, 19) <= input(3);
output(0, 20) <= input(4);
output(0, 21) <= input(5);
output(0, 22) <= input(6);
output(0, 23) <= input(7);
output(0, 24) <= input(8);
output(0, 25) <= input(9);
output(0, 26) <= input(10);
output(0, 27) <= input(11);
output(0, 28) <= input(12);
output(0, 29) <= input(13);
output(0, 30) <= input(14);
output(0, 31) <= input(15);
output(0, 32) <= input(0);
output(0, 33) <= input(1);
output(0, 34) <= input(2);
output(0, 35) <= input(3);
output(0, 36) <= input(4);
output(0, 37) <= input(5);
output(0, 38) <= input(6);
output(0, 39) <= input(7);
output(0, 40) <= input(8);
output(0, 41) <= input(9);
output(0, 42) <= input(10);
output(0, 43) <= input(11);
output(0, 44) <= input(12);
output(0, 45) <= input(13);
output(0, 46) <= input(14);
output(0, 47) <= input(15);
output(0, 48) <= input(16);
output(0, 49) <= input(17);
output(0, 50) <= input(18);
output(0, 51) <= input(19);
output(0, 52) <= input(20);
output(0, 53) <= input(21);
output(0, 54) <= input(22);
output(0, 55) <= input(23);
output(0, 56) <= input(24);
output(0, 57) <= input(25);
output(0, 58) <= input(26);
output(0, 59) <= input(27);
output(0, 60) <= input(28);
output(0, 61) <= input(29);
output(0, 62) <= input(30);
output(0, 63) <= input(31);
output(0, 64) <= input(16);
output(0, 65) <= input(17);
output(0, 66) <= input(18);
output(0, 67) <= input(19);
output(0, 68) <= input(20);
output(0, 69) <= input(21);
output(0, 70) <= input(22);
output(0, 71) <= input(23);
output(0, 72) <= input(24);
output(0, 73) <= input(25);
output(0, 74) <= input(26);
output(0, 75) <= input(27);
output(0, 76) <= input(28);
output(0, 77) <= input(29);
output(0, 78) <= input(30);
output(0, 79) <= input(31);
output(0, 80) <= input(16);
output(0, 81) <= input(17);
output(0, 82) <= input(18);
output(0, 83) <= input(19);
output(0, 84) <= input(20);
output(0, 85) <= input(21);
output(0, 86) <= input(22);
output(0, 87) <= input(23);
output(0, 88) <= input(24);
output(0, 89) <= input(25);
output(0, 90) <= input(26);
output(0, 91) <= input(27);
output(0, 92) <= input(28);
output(0, 93) <= input(29);
output(0, 94) <= input(30);
output(0, 95) <= input(31);
output(0, 96) <= input(16);
output(0, 97) <= input(17);
output(0, 98) <= input(18);
output(0, 99) <= input(19);
output(0, 100) <= input(20);
output(0, 101) <= input(21);
output(0, 102) <= input(22);
output(0, 103) <= input(23);
output(0, 104) <= input(24);
output(0, 105) <= input(25);
output(0, 106) <= input(26);
output(0, 107) <= input(27);
output(0, 108) <= input(28);
output(0, 109) <= input(29);
output(0, 110) <= input(30);
output(0, 111) <= input(31);
output(0, 112) <= input(1);
output(0, 113) <= input(2);
output(0, 114) <= input(3);
output(0, 115) <= input(4);
output(0, 116) <= input(5);
output(0, 117) <= input(6);
output(0, 118) <= input(7);
output(0, 119) <= input(8);
output(0, 120) <= input(9);
output(0, 121) <= input(10);
output(0, 122) <= input(11);
output(0, 123) <= input(12);
output(0, 124) <= input(13);
output(0, 125) <= input(14);
output(0, 126) <= input(15);
output(0, 127) <= input(32);
output(0, 128) <= input(1);
output(0, 129) <= input(2);
output(0, 130) <= input(3);
output(0, 131) <= input(4);
output(0, 132) <= input(5);
output(0, 133) <= input(6);
output(0, 134) <= input(7);
output(0, 135) <= input(8);
output(0, 136) <= input(9);
output(0, 137) <= input(10);
output(0, 138) <= input(11);
output(0, 139) <= input(12);
output(0, 140) <= input(13);
output(0, 141) <= input(14);
output(0, 142) <= input(15);
output(0, 143) <= input(32);
output(0, 144) <= input(1);
output(0, 145) <= input(2);
output(0, 146) <= input(3);
output(0, 147) <= input(4);
output(0, 148) <= input(5);
output(0, 149) <= input(6);
output(0, 150) <= input(7);
output(0, 151) <= input(8);
output(0, 152) <= input(9);
output(0, 153) <= input(10);
output(0, 154) <= input(11);
output(0, 155) <= input(12);
output(0, 156) <= input(13);
output(0, 157) <= input(14);
output(0, 158) <= input(15);
output(0, 159) <= input(32);
output(0, 160) <= input(1);
output(0, 161) <= input(2);
output(0, 162) <= input(3);
output(0, 163) <= input(4);
output(0, 164) <= input(5);
output(0, 165) <= input(6);
output(0, 166) <= input(7);
output(0, 167) <= input(8);
output(0, 168) <= input(9);
output(0, 169) <= input(10);
output(0, 170) <= input(11);
output(0, 171) <= input(12);
output(0, 172) <= input(13);
output(0, 173) <= input(14);
output(0, 174) <= input(15);
output(0, 175) <= input(32);
output(0, 176) <= input(17);
output(0, 177) <= input(18);
output(0, 178) <= input(19);
output(0, 179) <= input(20);
output(0, 180) <= input(21);
output(0, 181) <= input(22);
output(0, 182) <= input(23);
output(0, 183) <= input(24);
output(0, 184) <= input(25);
output(0, 185) <= input(26);
output(0, 186) <= input(27);
output(0, 187) <= input(28);
output(0, 188) <= input(29);
output(0, 189) <= input(30);
output(0, 190) <= input(31);
output(0, 191) <= input(33);
output(0, 192) <= input(17);
output(0, 193) <= input(18);
output(0, 194) <= input(19);
output(0, 195) <= input(20);
output(0, 196) <= input(21);
output(0, 197) <= input(22);
output(0, 198) <= input(23);
output(0, 199) <= input(24);
output(0, 200) <= input(25);
output(0, 201) <= input(26);
output(0, 202) <= input(27);
output(0, 203) <= input(28);
output(0, 204) <= input(29);
output(0, 205) <= input(30);
output(0, 206) <= input(31);
output(0, 207) <= input(33);
output(0, 208) <= input(17);
output(0, 209) <= input(18);
output(0, 210) <= input(19);
output(0, 211) <= input(20);
output(0, 212) <= input(21);
output(0, 213) <= input(22);
output(0, 214) <= input(23);
output(0, 215) <= input(24);
output(0, 216) <= input(25);
output(0, 217) <= input(26);
output(0, 218) <= input(27);
output(0, 219) <= input(28);
output(0, 220) <= input(29);
output(0, 221) <= input(30);
output(0, 222) <= input(31);
output(0, 223) <= input(33);
output(0, 224) <= input(17);
output(0, 225) <= input(18);
output(0, 226) <= input(19);
output(0, 227) <= input(20);
output(0, 228) <= input(21);
output(0, 229) <= input(22);
output(0, 230) <= input(23);
output(0, 231) <= input(24);
output(0, 232) <= input(25);
output(0, 233) <= input(26);
output(0, 234) <= input(27);
output(0, 235) <= input(28);
output(0, 236) <= input(29);
output(0, 237) <= input(30);
output(0, 238) <= input(31);
output(0, 239) <= input(33);
output(0, 240) <= input(2);
output(0, 241) <= input(3);
output(0, 242) <= input(4);
output(0, 243) <= input(5);
output(0, 244) <= input(6);
output(0, 245) <= input(7);
output(0, 246) <= input(8);
output(0, 247) <= input(9);
output(0, 248) <= input(10);
output(0, 249) <= input(11);
output(0, 250) <= input(12);
output(0, 251) <= input(13);
output(0, 252) <= input(14);
output(0, 253) <= input(15);
output(0, 254) <= input(32);
output(0, 255) <= input(34);
output(1, 0) <= input(35);
output(1, 1) <= input(16);
output(1, 2) <= input(17);
output(1, 3) <= input(18);
output(1, 4) <= input(19);
output(1, 5) <= input(20);
output(1, 6) <= input(21);
output(1, 7) <= input(22);
output(1, 8) <= input(23);
output(1, 9) <= input(24);
output(1, 10) <= input(25);
output(1, 11) <= input(26);
output(1, 12) <= input(27);
output(1, 13) <= input(28);
output(1, 14) <= input(29);
output(1, 15) <= input(30);
output(1, 16) <= input(35);
output(1, 17) <= input(16);
output(1, 18) <= input(17);
output(1, 19) <= input(18);
output(1, 20) <= input(19);
output(1, 21) <= input(20);
output(1, 22) <= input(21);
output(1, 23) <= input(22);
output(1, 24) <= input(23);
output(1, 25) <= input(24);
output(1, 26) <= input(25);
output(1, 27) <= input(26);
output(1, 28) <= input(27);
output(1, 29) <= input(28);
output(1, 30) <= input(29);
output(1, 31) <= input(30);
output(1, 32) <= input(35);
output(1, 33) <= input(16);
output(1, 34) <= input(17);
output(1, 35) <= input(18);
output(1, 36) <= input(19);
output(1, 37) <= input(20);
output(1, 38) <= input(21);
output(1, 39) <= input(22);
output(1, 40) <= input(23);
output(1, 41) <= input(24);
output(1, 42) <= input(25);
output(1, 43) <= input(26);
output(1, 44) <= input(27);
output(1, 45) <= input(28);
output(1, 46) <= input(29);
output(1, 47) <= input(30);
output(1, 48) <= input(35);
output(1, 49) <= input(16);
output(1, 50) <= input(17);
output(1, 51) <= input(18);
output(1, 52) <= input(19);
output(1, 53) <= input(20);
output(1, 54) <= input(21);
output(1, 55) <= input(22);
output(1, 56) <= input(23);
output(1, 57) <= input(24);
output(1, 58) <= input(25);
output(1, 59) <= input(26);
output(1, 60) <= input(27);
output(1, 61) <= input(28);
output(1, 62) <= input(29);
output(1, 63) <= input(30);
output(1, 64) <= input(35);
output(1, 65) <= input(16);
output(1, 66) <= input(17);
output(1, 67) <= input(18);
output(1, 68) <= input(19);
output(1, 69) <= input(20);
output(1, 70) <= input(21);
output(1, 71) <= input(22);
output(1, 72) <= input(23);
output(1, 73) <= input(24);
output(1, 74) <= input(25);
output(1, 75) <= input(26);
output(1, 76) <= input(27);
output(1, 77) <= input(28);
output(1, 78) <= input(29);
output(1, 79) <= input(30);
output(1, 80) <= input(0);
output(1, 81) <= input(1);
output(1, 82) <= input(2);
output(1, 83) <= input(3);
output(1, 84) <= input(4);
output(1, 85) <= input(5);
output(1, 86) <= input(6);
output(1, 87) <= input(7);
output(1, 88) <= input(8);
output(1, 89) <= input(9);
output(1, 90) <= input(10);
output(1, 91) <= input(11);
output(1, 92) <= input(12);
output(1, 93) <= input(13);
output(1, 94) <= input(14);
output(1, 95) <= input(15);
output(1, 96) <= input(0);
output(1, 97) <= input(1);
output(1, 98) <= input(2);
output(1, 99) <= input(3);
output(1, 100) <= input(4);
output(1, 101) <= input(5);
output(1, 102) <= input(6);
output(1, 103) <= input(7);
output(1, 104) <= input(8);
output(1, 105) <= input(9);
output(1, 106) <= input(10);
output(1, 107) <= input(11);
output(1, 108) <= input(12);
output(1, 109) <= input(13);
output(1, 110) <= input(14);
output(1, 111) <= input(15);
output(1, 112) <= input(0);
output(1, 113) <= input(1);
output(1, 114) <= input(2);
output(1, 115) <= input(3);
output(1, 116) <= input(4);
output(1, 117) <= input(5);
output(1, 118) <= input(6);
output(1, 119) <= input(7);
output(1, 120) <= input(8);
output(1, 121) <= input(9);
output(1, 122) <= input(10);
output(1, 123) <= input(11);
output(1, 124) <= input(12);
output(1, 125) <= input(13);
output(1, 126) <= input(14);
output(1, 127) <= input(15);
output(1, 128) <= input(0);
output(1, 129) <= input(1);
output(1, 130) <= input(2);
output(1, 131) <= input(3);
output(1, 132) <= input(4);
output(1, 133) <= input(5);
output(1, 134) <= input(6);
output(1, 135) <= input(7);
output(1, 136) <= input(8);
output(1, 137) <= input(9);
output(1, 138) <= input(10);
output(1, 139) <= input(11);
output(1, 140) <= input(12);
output(1, 141) <= input(13);
output(1, 142) <= input(14);
output(1, 143) <= input(15);
output(1, 144) <= input(0);
output(1, 145) <= input(1);
output(1, 146) <= input(2);
output(1, 147) <= input(3);
output(1, 148) <= input(4);
output(1, 149) <= input(5);
output(1, 150) <= input(6);
output(1, 151) <= input(7);
output(1, 152) <= input(8);
output(1, 153) <= input(9);
output(1, 154) <= input(10);
output(1, 155) <= input(11);
output(1, 156) <= input(12);
output(1, 157) <= input(13);
output(1, 158) <= input(14);
output(1, 159) <= input(15);
output(1, 160) <= input(16);
output(1, 161) <= input(17);
output(1, 162) <= input(18);
output(1, 163) <= input(19);
output(1, 164) <= input(20);
output(1, 165) <= input(21);
output(1, 166) <= input(22);
output(1, 167) <= input(23);
output(1, 168) <= input(24);
output(1, 169) <= input(25);
output(1, 170) <= input(26);
output(1, 171) <= input(27);
output(1, 172) <= input(28);
output(1, 173) <= input(29);
output(1, 174) <= input(30);
output(1, 175) <= input(31);
output(1, 176) <= input(16);
output(1, 177) <= input(17);
output(1, 178) <= input(18);
output(1, 179) <= input(19);
output(1, 180) <= input(20);
output(1, 181) <= input(21);
output(1, 182) <= input(22);
output(1, 183) <= input(23);
output(1, 184) <= input(24);
output(1, 185) <= input(25);
output(1, 186) <= input(26);
output(1, 187) <= input(27);
output(1, 188) <= input(28);
output(1, 189) <= input(29);
output(1, 190) <= input(30);
output(1, 191) <= input(31);
output(1, 192) <= input(16);
output(1, 193) <= input(17);
output(1, 194) <= input(18);
output(1, 195) <= input(19);
output(1, 196) <= input(20);
output(1, 197) <= input(21);
output(1, 198) <= input(22);
output(1, 199) <= input(23);
output(1, 200) <= input(24);
output(1, 201) <= input(25);
output(1, 202) <= input(26);
output(1, 203) <= input(27);
output(1, 204) <= input(28);
output(1, 205) <= input(29);
output(1, 206) <= input(30);
output(1, 207) <= input(31);
output(1, 208) <= input(16);
output(1, 209) <= input(17);
output(1, 210) <= input(18);
output(1, 211) <= input(19);
output(1, 212) <= input(20);
output(1, 213) <= input(21);
output(1, 214) <= input(22);
output(1, 215) <= input(23);
output(1, 216) <= input(24);
output(1, 217) <= input(25);
output(1, 218) <= input(26);
output(1, 219) <= input(27);
output(1, 220) <= input(28);
output(1, 221) <= input(29);
output(1, 222) <= input(30);
output(1, 223) <= input(31);
output(1, 224) <= input(16);
output(1, 225) <= input(17);
output(1, 226) <= input(18);
output(1, 227) <= input(19);
output(1, 228) <= input(20);
output(1, 229) <= input(21);
output(1, 230) <= input(22);
output(1, 231) <= input(23);
output(1, 232) <= input(24);
output(1, 233) <= input(25);
output(1, 234) <= input(26);
output(1, 235) <= input(27);
output(1, 236) <= input(28);
output(1, 237) <= input(29);
output(1, 238) <= input(30);
output(1, 239) <= input(31);
output(1, 240) <= input(1);
output(1, 241) <= input(2);
output(1, 242) <= input(3);
output(1, 243) <= input(4);
output(1, 244) <= input(5);
output(1, 245) <= input(6);
output(1, 246) <= input(7);
output(1, 247) <= input(8);
output(1, 248) <= input(9);
output(1, 249) <= input(10);
output(1, 250) <= input(11);
output(1, 251) <= input(12);
output(1, 252) <= input(13);
output(1, 253) <= input(14);
output(1, 254) <= input(15);
output(1, 255) <= input(32);
output(2, 0) <= input(36);
output(2, 1) <= input(0);
output(2, 2) <= input(1);
output(2, 3) <= input(2);
output(2, 4) <= input(3);
output(2, 5) <= input(4);
output(2, 6) <= input(5);
output(2, 7) <= input(6);
output(2, 8) <= input(7);
output(2, 9) <= input(8);
output(2, 10) <= input(9);
output(2, 11) <= input(10);
output(2, 12) <= input(11);
output(2, 13) <= input(12);
output(2, 14) <= input(13);
output(2, 15) <= input(14);
output(2, 16) <= input(36);
output(2, 17) <= input(0);
output(2, 18) <= input(1);
output(2, 19) <= input(2);
output(2, 20) <= input(3);
output(2, 21) <= input(4);
output(2, 22) <= input(5);
output(2, 23) <= input(6);
output(2, 24) <= input(7);
output(2, 25) <= input(8);
output(2, 26) <= input(9);
output(2, 27) <= input(10);
output(2, 28) <= input(11);
output(2, 29) <= input(12);
output(2, 30) <= input(13);
output(2, 31) <= input(14);
output(2, 32) <= input(36);
output(2, 33) <= input(0);
output(2, 34) <= input(1);
output(2, 35) <= input(2);
output(2, 36) <= input(3);
output(2, 37) <= input(4);
output(2, 38) <= input(5);
output(2, 39) <= input(6);
output(2, 40) <= input(7);
output(2, 41) <= input(8);
output(2, 42) <= input(9);
output(2, 43) <= input(10);
output(2, 44) <= input(11);
output(2, 45) <= input(12);
output(2, 46) <= input(13);
output(2, 47) <= input(14);
output(2, 48) <= input(36);
output(2, 49) <= input(0);
output(2, 50) <= input(1);
output(2, 51) <= input(2);
output(2, 52) <= input(3);
output(2, 53) <= input(4);
output(2, 54) <= input(5);
output(2, 55) <= input(6);
output(2, 56) <= input(7);
output(2, 57) <= input(8);
output(2, 58) <= input(9);
output(2, 59) <= input(10);
output(2, 60) <= input(11);
output(2, 61) <= input(12);
output(2, 62) <= input(13);
output(2, 63) <= input(14);
output(2, 64) <= input(36);
output(2, 65) <= input(0);
output(2, 66) <= input(1);
output(2, 67) <= input(2);
output(2, 68) <= input(3);
output(2, 69) <= input(4);
output(2, 70) <= input(5);
output(2, 71) <= input(6);
output(2, 72) <= input(7);
output(2, 73) <= input(8);
output(2, 74) <= input(9);
output(2, 75) <= input(10);
output(2, 76) <= input(11);
output(2, 77) <= input(12);
output(2, 78) <= input(13);
output(2, 79) <= input(14);
output(2, 80) <= input(36);
output(2, 81) <= input(0);
output(2, 82) <= input(1);
output(2, 83) <= input(2);
output(2, 84) <= input(3);
output(2, 85) <= input(4);
output(2, 86) <= input(5);
output(2, 87) <= input(6);
output(2, 88) <= input(7);
output(2, 89) <= input(8);
output(2, 90) <= input(9);
output(2, 91) <= input(10);
output(2, 92) <= input(11);
output(2, 93) <= input(12);
output(2, 94) <= input(13);
output(2, 95) <= input(14);
output(2, 96) <= input(36);
output(2, 97) <= input(0);
output(2, 98) <= input(1);
output(2, 99) <= input(2);
output(2, 100) <= input(3);
output(2, 101) <= input(4);
output(2, 102) <= input(5);
output(2, 103) <= input(6);
output(2, 104) <= input(7);
output(2, 105) <= input(8);
output(2, 106) <= input(9);
output(2, 107) <= input(10);
output(2, 108) <= input(11);
output(2, 109) <= input(12);
output(2, 110) <= input(13);
output(2, 111) <= input(14);
output(2, 112) <= input(35);
output(2, 113) <= input(16);
output(2, 114) <= input(17);
output(2, 115) <= input(18);
output(2, 116) <= input(19);
output(2, 117) <= input(20);
output(2, 118) <= input(21);
output(2, 119) <= input(22);
output(2, 120) <= input(23);
output(2, 121) <= input(24);
output(2, 122) <= input(25);
output(2, 123) <= input(26);
output(2, 124) <= input(27);
output(2, 125) <= input(28);
output(2, 126) <= input(29);
output(2, 127) <= input(30);
output(2, 128) <= input(35);
output(2, 129) <= input(16);
output(2, 130) <= input(17);
output(2, 131) <= input(18);
output(2, 132) <= input(19);
output(2, 133) <= input(20);
output(2, 134) <= input(21);
output(2, 135) <= input(22);
output(2, 136) <= input(23);
output(2, 137) <= input(24);
output(2, 138) <= input(25);
output(2, 139) <= input(26);
output(2, 140) <= input(27);
output(2, 141) <= input(28);
output(2, 142) <= input(29);
output(2, 143) <= input(30);
output(2, 144) <= input(35);
output(2, 145) <= input(16);
output(2, 146) <= input(17);
output(2, 147) <= input(18);
output(2, 148) <= input(19);
output(2, 149) <= input(20);
output(2, 150) <= input(21);
output(2, 151) <= input(22);
output(2, 152) <= input(23);
output(2, 153) <= input(24);
output(2, 154) <= input(25);
output(2, 155) <= input(26);
output(2, 156) <= input(27);
output(2, 157) <= input(28);
output(2, 158) <= input(29);
output(2, 159) <= input(30);
output(2, 160) <= input(35);
output(2, 161) <= input(16);
output(2, 162) <= input(17);
output(2, 163) <= input(18);
output(2, 164) <= input(19);
output(2, 165) <= input(20);
output(2, 166) <= input(21);
output(2, 167) <= input(22);
output(2, 168) <= input(23);
output(2, 169) <= input(24);
output(2, 170) <= input(25);
output(2, 171) <= input(26);
output(2, 172) <= input(27);
output(2, 173) <= input(28);
output(2, 174) <= input(29);
output(2, 175) <= input(30);
output(2, 176) <= input(35);
output(2, 177) <= input(16);
output(2, 178) <= input(17);
output(2, 179) <= input(18);
output(2, 180) <= input(19);
output(2, 181) <= input(20);
output(2, 182) <= input(21);
output(2, 183) <= input(22);
output(2, 184) <= input(23);
output(2, 185) <= input(24);
output(2, 186) <= input(25);
output(2, 187) <= input(26);
output(2, 188) <= input(27);
output(2, 189) <= input(28);
output(2, 190) <= input(29);
output(2, 191) <= input(30);
output(2, 192) <= input(35);
output(2, 193) <= input(16);
output(2, 194) <= input(17);
output(2, 195) <= input(18);
output(2, 196) <= input(19);
output(2, 197) <= input(20);
output(2, 198) <= input(21);
output(2, 199) <= input(22);
output(2, 200) <= input(23);
output(2, 201) <= input(24);
output(2, 202) <= input(25);
output(2, 203) <= input(26);
output(2, 204) <= input(27);
output(2, 205) <= input(28);
output(2, 206) <= input(29);
output(2, 207) <= input(30);
output(2, 208) <= input(35);
output(2, 209) <= input(16);
output(2, 210) <= input(17);
output(2, 211) <= input(18);
output(2, 212) <= input(19);
output(2, 213) <= input(20);
output(2, 214) <= input(21);
output(2, 215) <= input(22);
output(2, 216) <= input(23);
output(2, 217) <= input(24);
output(2, 218) <= input(25);
output(2, 219) <= input(26);
output(2, 220) <= input(27);
output(2, 221) <= input(28);
output(2, 222) <= input(29);
output(2, 223) <= input(30);
output(2, 224) <= input(35);
output(2, 225) <= input(16);
output(2, 226) <= input(17);
output(2, 227) <= input(18);
output(2, 228) <= input(19);
output(2, 229) <= input(20);
output(2, 230) <= input(21);
output(2, 231) <= input(22);
output(2, 232) <= input(23);
output(2, 233) <= input(24);
output(2, 234) <= input(25);
output(2, 235) <= input(26);
output(2, 236) <= input(27);
output(2, 237) <= input(28);
output(2, 238) <= input(29);
output(2, 239) <= input(30);
output(2, 240) <= input(0);
output(2, 241) <= input(1);
output(2, 242) <= input(2);
output(2, 243) <= input(3);
output(2, 244) <= input(4);
output(2, 245) <= input(5);
output(2, 246) <= input(6);
output(2, 247) <= input(7);
output(2, 248) <= input(8);
output(2, 249) <= input(9);
output(2, 250) <= input(10);
output(2, 251) <= input(11);
output(2, 252) <= input(12);
output(2, 253) <= input(13);
output(2, 254) <= input(14);
output(2, 255) <= input(15);
output(3, 0) <= input(37);
output(3, 1) <= input(35);
output(3, 2) <= input(16);
output(3, 3) <= input(17);
output(3, 4) <= input(18);
output(3, 5) <= input(19);
output(3, 6) <= input(20);
output(3, 7) <= input(21);
output(3, 8) <= input(22);
output(3, 9) <= input(23);
output(3, 10) <= input(24);
output(3, 11) <= input(25);
output(3, 12) <= input(26);
output(3, 13) <= input(27);
output(3, 14) <= input(28);
output(3, 15) <= input(29);
output(3, 16) <= input(37);
output(3, 17) <= input(35);
output(3, 18) <= input(16);
output(3, 19) <= input(17);
output(3, 20) <= input(18);
output(3, 21) <= input(19);
output(3, 22) <= input(20);
output(3, 23) <= input(21);
output(3, 24) <= input(22);
output(3, 25) <= input(23);
output(3, 26) <= input(24);
output(3, 27) <= input(25);
output(3, 28) <= input(26);
output(3, 29) <= input(27);
output(3, 30) <= input(28);
output(3, 31) <= input(29);
output(3, 32) <= input(37);
output(3, 33) <= input(35);
output(3, 34) <= input(16);
output(3, 35) <= input(17);
output(3, 36) <= input(18);
output(3, 37) <= input(19);
output(3, 38) <= input(20);
output(3, 39) <= input(21);
output(3, 40) <= input(22);
output(3, 41) <= input(23);
output(3, 42) <= input(24);
output(3, 43) <= input(25);
output(3, 44) <= input(26);
output(3, 45) <= input(27);
output(3, 46) <= input(28);
output(3, 47) <= input(29);
output(3, 48) <= input(37);
output(3, 49) <= input(35);
output(3, 50) <= input(16);
output(3, 51) <= input(17);
output(3, 52) <= input(18);
output(3, 53) <= input(19);
output(3, 54) <= input(20);
output(3, 55) <= input(21);
output(3, 56) <= input(22);
output(3, 57) <= input(23);
output(3, 58) <= input(24);
output(3, 59) <= input(25);
output(3, 60) <= input(26);
output(3, 61) <= input(27);
output(3, 62) <= input(28);
output(3, 63) <= input(29);
output(3, 64) <= input(37);
output(3, 65) <= input(35);
output(3, 66) <= input(16);
output(3, 67) <= input(17);
output(3, 68) <= input(18);
output(3, 69) <= input(19);
output(3, 70) <= input(20);
output(3, 71) <= input(21);
output(3, 72) <= input(22);
output(3, 73) <= input(23);
output(3, 74) <= input(24);
output(3, 75) <= input(25);
output(3, 76) <= input(26);
output(3, 77) <= input(27);
output(3, 78) <= input(28);
output(3, 79) <= input(29);
output(3, 80) <= input(37);
output(3, 81) <= input(35);
output(3, 82) <= input(16);
output(3, 83) <= input(17);
output(3, 84) <= input(18);
output(3, 85) <= input(19);
output(3, 86) <= input(20);
output(3, 87) <= input(21);
output(3, 88) <= input(22);
output(3, 89) <= input(23);
output(3, 90) <= input(24);
output(3, 91) <= input(25);
output(3, 92) <= input(26);
output(3, 93) <= input(27);
output(3, 94) <= input(28);
output(3, 95) <= input(29);
output(3, 96) <= input(37);
output(3, 97) <= input(35);
output(3, 98) <= input(16);
output(3, 99) <= input(17);
output(3, 100) <= input(18);
output(3, 101) <= input(19);
output(3, 102) <= input(20);
output(3, 103) <= input(21);
output(3, 104) <= input(22);
output(3, 105) <= input(23);
output(3, 106) <= input(24);
output(3, 107) <= input(25);
output(3, 108) <= input(26);
output(3, 109) <= input(27);
output(3, 110) <= input(28);
output(3, 111) <= input(29);
output(3, 112) <= input(37);
output(3, 113) <= input(35);
output(3, 114) <= input(16);
output(3, 115) <= input(17);
output(3, 116) <= input(18);
output(3, 117) <= input(19);
output(3, 118) <= input(20);
output(3, 119) <= input(21);
output(3, 120) <= input(22);
output(3, 121) <= input(23);
output(3, 122) <= input(24);
output(3, 123) <= input(25);
output(3, 124) <= input(26);
output(3, 125) <= input(27);
output(3, 126) <= input(28);
output(3, 127) <= input(29);
output(3, 128) <= input(37);
output(3, 129) <= input(35);
output(3, 130) <= input(16);
output(3, 131) <= input(17);
output(3, 132) <= input(18);
output(3, 133) <= input(19);
output(3, 134) <= input(20);
output(3, 135) <= input(21);
output(3, 136) <= input(22);
output(3, 137) <= input(23);
output(3, 138) <= input(24);
output(3, 139) <= input(25);
output(3, 140) <= input(26);
output(3, 141) <= input(27);
output(3, 142) <= input(28);
output(3, 143) <= input(29);
output(3, 144) <= input(37);
output(3, 145) <= input(35);
output(3, 146) <= input(16);
output(3, 147) <= input(17);
output(3, 148) <= input(18);
output(3, 149) <= input(19);
output(3, 150) <= input(20);
output(3, 151) <= input(21);
output(3, 152) <= input(22);
output(3, 153) <= input(23);
output(3, 154) <= input(24);
output(3, 155) <= input(25);
output(3, 156) <= input(26);
output(3, 157) <= input(27);
output(3, 158) <= input(28);
output(3, 159) <= input(29);
output(3, 160) <= input(37);
output(3, 161) <= input(35);
output(3, 162) <= input(16);
output(3, 163) <= input(17);
output(3, 164) <= input(18);
output(3, 165) <= input(19);
output(3, 166) <= input(20);
output(3, 167) <= input(21);
output(3, 168) <= input(22);
output(3, 169) <= input(23);
output(3, 170) <= input(24);
output(3, 171) <= input(25);
output(3, 172) <= input(26);
output(3, 173) <= input(27);
output(3, 174) <= input(28);
output(3, 175) <= input(29);
output(3, 176) <= input(37);
output(3, 177) <= input(35);
output(3, 178) <= input(16);
output(3, 179) <= input(17);
output(3, 180) <= input(18);
output(3, 181) <= input(19);
output(3, 182) <= input(20);
output(3, 183) <= input(21);
output(3, 184) <= input(22);
output(3, 185) <= input(23);
output(3, 186) <= input(24);
output(3, 187) <= input(25);
output(3, 188) <= input(26);
output(3, 189) <= input(27);
output(3, 190) <= input(28);
output(3, 191) <= input(29);
output(3, 192) <= input(37);
output(3, 193) <= input(35);
output(3, 194) <= input(16);
output(3, 195) <= input(17);
output(3, 196) <= input(18);
output(3, 197) <= input(19);
output(3, 198) <= input(20);
output(3, 199) <= input(21);
output(3, 200) <= input(22);
output(3, 201) <= input(23);
output(3, 202) <= input(24);
output(3, 203) <= input(25);
output(3, 204) <= input(26);
output(3, 205) <= input(27);
output(3, 206) <= input(28);
output(3, 207) <= input(29);
output(3, 208) <= input(37);
output(3, 209) <= input(35);
output(3, 210) <= input(16);
output(3, 211) <= input(17);
output(3, 212) <= input(18);
output(3, 213) <= input(19);
output(3, 214) <= input(20);
output(3, 215) <= input(21);
output(3, 216) <= input(22);
output(3, 217) <= input(23);
output(3, 218) <= input(24);
output(3, 219) <= input(25);
output(3, 220) <= input(26);
output(3, 221) <= input(27);
output(3, 222) <= input(28);
output(3, 223) <= input(29);
output(3, 224) <= input(37);
output(3, 225) <= input(35);
output(3, 226) <= input(16);
output(3, 227) <= input(17);
output(3, 228) <= input(18);
output(3, 229) <= input(19);
output(3, 230) <= input(20);
output(3, 231) <= input(21);
output(3, 232) <= input(22);
output(3, 233) <= input(23);
output(3, 234) <= input(24);
output(3, 235) <= input(25);
output(3, 236) <= input(26);
output(3, 237) <= input(27);
output(3, 238) <= input(28);
output(3, 239) <= input(29);
output(3, 240) <= input(36);
output(3, 241) <= input(0);
output(3, 242) <= input(1);
output(3, 243) <= input(2);
output(3, 244) <= input(3);
output(3, 245) <= input(4);
output(3, 246) <= input(5);
output(3, 247) <= input(6);
output(3, 248) <= input(7);
output(3, 249) <= input(8);
output(3, 250) <= input(9);
output(3, 251) <= input(10);
output(3, 252) <= input(11);
output(3, 253) <= input(12);
output(3, 254) <= input(13);
output(3, 255) <= input(14);
output(4, 0) <= input(38);
output(4, 1) <= input(36);
output(4, 2) <= input(0);
output(4, 3) <= input(1);
output(4, 4) <= input(2);
output(4, 5) <= input(3);
output(4, 6) <= input(4);
output(4, 7) <= input(5);
output(4, 8) <= input(6);
output(4, 9) <= input(7);
output(4, 10) <= input(8);
output(4, 11) <= input(9);
output(4, 12) <= input(10);
output(4, 13) <= input(11);
output(4, 14) <= input(12);
output(4, 15) <= input(13);
output(4, 16) <= input(38);
output(4, 17) <= input(36);
output(4, 18) <= input(0);
output(4, 19) <= input(1);
output(4, 20) <= input(2);
output(4, 21) <= input(3);
output(4, 22) <= input(4);
output(4, 23) <= input(5);
output(4, 24) <= input(6);
output(4, 25) <= input(7);
output(4, 26) <= input(8);
output(4, 27) <= input(9);
output(4, 28) <= input(10);
output(4, 29) <= input(11);
output(4, 30) <= input(12);
output(4, 31) <= input(13);
output(4, 32) <= input(38);
output(4, 33) <= input(36);
output(4, 34) <= input(0);
output(4, 35) <= input(1);
output(4, 36) <= input(2);
output(4, 37) <= input(3);
output(4, 38) <= input(4);
output(4, 39) <= input(5);
output(4, 40) <= input(6);
output(4, 41) <= input(7);
output(4, 42) <= input(8);
output(4, 43) <= input(9);
output(4, 44) <= input(10);
output(4, 45) <= input(11);
output(4, 46) <= input(12);
output(4, 47) <= input(13);
output(4, 48) <= input(38);
output(4, 49) <= input(36);
output(4, 50) <= input(0);
output(4, 51) <= input(1);
output(4, 52) <= input(2);
output(4, 53) <= input(3);
output(4, 54) <= input(4);
output(4, 55) <= input(5);
output(4, 56) <= input(6);
output(4, 57) <= input(7);
output(4, 58) <= input(8);
output(4, 59) <= input(9);
output(4, 60) <= input(10);
output(4, 61) <= input(11);
output(4, 62) <= input(12);
output(4, 63) <= input(13);
output(4, 64) <= input(38);
output(4, 65) <= input(36);
output(4, 66) <= input(0);
output(4, 67) <= input(1);
output(4, 68) <= input(2);
output(4, 69) <= input(3);
output(4, 70) <= input(4);
output(4, 71) <= input(5);
output(4, 72) <= input(6);
output(4, 73) <= input(7);
output(4, 74) <= input(8);
output(4, 75) <= input(9);
output(4, 76) <= input(10);
output(4, 77) <= input(11);
output(4, 78) <= input(12);
output(4, 79) <= input(13);
output(4, 80) <= input(38);
output(4, 81) <= input(36);
output(4, 82) <= input(0);
output(4, 83) <= input(1);
output(4, 84) <= input(2);
output(4, 85) <= input(3);
output(4, 86) <= input(4);
output(4, 87) <= input(5);
output(4, 88) <= input(6);
output(4, 89) <= input(7);
output(4, 90) <= input(8);
output(4, 91) <= input(9);
output(4, 92) <= input(10);
output(4, 93) <= input(11);
output(4, 94) <= input(12);
output(4, 95) <= input(13);
output(4, 96) <= input(38);
output(4, 97) <= input(36);
output(4, 98) <= input(0);
output(4, 99) <= input(1);
output(4, 100) <= input(2);
output(4, 101) <= input(3);
output(4, 102) <= input(4);
output(4, 103) <= input(5);
output(4, 104) <= input(6);
output(4, 105) <= input(7);
output(4, 106) <= input(8);
output(4, 107) <= input(9);
output(4, 108) <= input(10);
output(4, 109) <= input(11);
output(4, 110) <= input(12);
output(4, 111) <= input(13);
output(4, 112) <= input(38);
output(4, 113) <= input(36);
output(4, 114) <= input(0);
output(4, 115) <= input(1);
output(4, 116) <= input(2);
output(4, 117) <= input(3);
output(4, 118) <= input(4);
output(4, 119) <= input(5);
output(4, 120) <= input(6);
output(4, 121) <= input(7);
output(4, 122) <= input(8);
output(4, 123) <= input(9);
output(4, 124) <= input(10);
output(4, 125) <= input(11);
output(4, 126) <= input(12);
output(4, 127) <= input(13);
output(4, 128) <= input(38);
output(4, 129) <= input(36);
output(4, 130) <= input(0);
output(4, 131) <= input(1);
output(4, 132) <= input(2);
output(4, 133) <= input(3);
output(4, 134) <= input(4);
output(4, 135) <= input(5);
output(4, 136) <= input(6);
output(4, 137) <= input(7);
output(4, 138) <= input(8);
output(4, 139) <= input(9);
output(4, 140) <= input(10);
output(4, 141) <= input(11);
output(4, 142) <= input(12);
output(4, 143) <= input(13);
output(4, 144) <= input(38);
output(4, 145) <= input(36);
output(4, 146) <= input(0);
output(4, 147) <= input(1);
output(4, 148) <= input(2);
output(4, 149) <= input(3);
output(4, 150) <= input(4);
output(4, 151) <= input(5);
output(4, 152) <= input(6);
output(4, 153) <= input(7);
output(4, 154) <= input(8);
output(4, 155) <= input(9);
output(4, 156) <= input(10);
output(4, 157) <= input(11);
output(4, 158) <= input(12);
output(4, 159) <= input(13);
output(4, 160) <= input(38);
output(4, 161) <= input(36);
output(4, 162) <= input(0);
output(4, 163) <= input(1);
output(4, 164) <= input(2);
output(4, 165) <= input(3);
output(4, 166) <= input(4);
output(4, 167) <= input(5);
output(4, 168) <= input(6);
output(4, 169) <= input(7);
output(4, 170) <= input(8);
output(4, 171) <= input(9);
output(4, 172) <= input(10);
output(4, 173) <= input(11);
output(4, 174) <= input(12);
output(4, 175) <= input(13);
output(4, 176) <= input(38);
output(4, 177) <= input(36);
output(4, 178) <= input(0);
output(4, 179) <= input(1);
output(4, 180) <= input(2);
output(4, 181) <= input(3);
output(4, 182) <= input(4);
output(4, 183) <= input(5);
output(4, 184) <= input(6);
output(4, 185) <= input(7);
output(4, 186) <= input(8);
output(4, 187) <= input(9);
output(4, 188) <= input(10);
output(4, 189) <= input(11);
output(4, 190) <= input(12);
output(4, 191) <= input(13);
output(4, 192) <= input(38);
output(4, 193) <= input(36);
output(4, 194) <= input(0);
output(4, 195) <= input(1);
output(4, 196) <= input(2);
output(4, 197) <= input(3);
output(4, 198) <= input(4);
output(4, 199) <= input(5);
output(4, 200) <= input(6);
output(4, 201) <= input(7);
output(4, 202) <= input(8);
output(4, 203) <= input(9);
output(4, 204) <= input(10);
output(4, 205) <= input(11);
output(4, 206) <= input(12);
output(4, 207) <= input(13);
output(4, 208) <= input(38);
output(4, 209) <= input(36);
output(4, 210) <= input(0);
output(4, 211) <= input(1);
output(4, 212) <= input(2);
output(4, 213) <= input(3);
output(4, 214) <= input(4);
output(4, 215) <= input(5);
output(4, 216) <= input(6);
output(4, 217) <= input(7);
output(4, 218) <= input(8);
output(4, 219) <= input(9);
output(4, 220) <= input(10);
output(4, 221) <= input(11);
output(4, 222) <= input(12);
output(4, 223) <= input(13);
output(4, 224) <= input(38);
output(4, 225) <= input(36);
output(4, 226) <= input(0);
output(4, 227) <= input(1);
output(4, 228) <= input(2);
output(4, 229) <= input(3);
output(4, 230) <= input(4);
output(4, 231) <= input(5);
output(4, 232) <= input(6);
output(4, 233) <= input(7);
output(4, 234) <= input(8);
output(4, 235) <= input(9);
output(4, 236) <= input(10);
output(4, 237) <= input(11);
output(4, 238) <= input(12);
output(4, 239) <= input(13);
output(4, 240) <= input(38);
output(4, 241) <= input(36);
output(4, 242) <= input(0);
output(4, 243) <= input(1);
output(4, 244) <= input(2);
output(4, 245) <= input(3);
output(4, 246) <= input(4);
output(4, 247) <= input(5);
output(4, 248) <= input(6);
output(4, 249) <= input(7);
output(4, 250) <= input(8);
output(4, 251) <= input(9);
output(4, 252) <= input(10);
output(4, 253) <= input(11);
output(4, 254) <= input(12);
output(4, 255) <= input(13);
output(5, 0) <= input(39);
output(5, 1) <= input(38);
output(5, 2) <= input(36);
output(5, 3) <= input(0);
output(5, 4) <= input(1);
output(5, 5) <= input(2);
output(5, 6) <= input(3);
output(5, 7) <= input(4);
output(5, 8) <= input(5);
output(5, 9) <= input(6);
output(5, 10) <= input(7);
output(5, 11) <= input(8);
output(5, 12) <= input(9);
output(5, 13) <= input(10);
output(5, 14) <= input(11);
output(5, 15) <= input(12);
output(5, 16) <= input(39);
output(5, 17) <= input(38);
output(5, 18) <= input(36);
output(5, 19) <= input(0);
output(5, 20) <= input(1);
output(5, 21) <= input(2);
output(5, 22) <= input(3);
output(5, 23) <= input(4);
output(5, 24) <= input(5);
output(5, 25) <= input(6);
output(5, 26) <= input(7);
output(5, 27) <= input(8);
output(5, 28) <= input(9);
output(5, 29) <= input(10);
output(5, 30) <= input(11);
output(5, 31) <= input(12);
output(5, 32) <= input(39);
output(5, 33) <= input(38);
output(5, 34) <= input(36);
output(5, 35) <= input(0);
output(5, 36) <= input(1);
output(5, 37) <= input(2);
output(5, 38) <= input(3);
output(5, 39) <= input(4);
output(5, 40) <= input(5);
output(5, 41) <= input(6);
output(5, 42) <= input(7);
output(5, 43) <= input(8);
output(5, 44) <= input(9);
output(5, 45) <= input(10);
output(5, 46) <= input(11);
output(5, 47) <= input(12);
output(5, 48) <= input(39);
output(5, 49) <= input(38);
output(5, 50) <= input(36);
output(5, 51) <= input(0);
output(5, 52) <= input(1);
output(5, 53) <= input(2);
output(5, 54) <= input(3);
output(5, 55) <= input(4);
output(5, 56) <= input(5);
output(5, 57) <= input(6);
output(5, 58) <= input(7);
output(5, 59) <= input(8);
output(5, 60) <= input(9);
output(5, 61) <= input(10);
output(5, 62) <= input(11);
output(5, 63) <= input(12);
output(5, 64) <= input(39);
output(5, 65) <= input(38);
output(5, 66) <= input(36);
output(5, 67) <= input(0);
output(5, 68) <= input(1);
output(5, 69) <= input(2);
output(5, 70) <= input(3);
output(5, 71) <= input(4);
output(5, 72) <= input(5);
output(5, 73) <= input(6);
output(5, 74) <= input(7);
output(5, 75) <= input(8);
output(5, 76) <= input(9);
output(5, 77) <= input(10);
output(5, 78) <= input(11);
output(5, 79) <= input(12);
output(5, 80) <= input(39);
output(5, 81) <= input(38);
output(5, 82) <= input(36);
output(5, 83) <= input(0);
output(5, 84) <= input(1);
output(5, 85) <= input(2);
output(5, 86) <= input(3);
output(5, 87) <= input(4);
output(5, 88) <= input(5);
output(5, 89) <= input(6);
output(5, 90) <= input(7);
output(5, 91) <= input(8);
output(5, 92) <= input(9);
output(5, 93) <= input(10);
output(5, 94) <= input(11);
output(5, 95) <= input(12);
output(5, 96) <= input(39);
output(5, 97) <= input(38);
output(5, 98) <= input(36);
output(5, 99) <= input(0);
output(5, 100) <= input(1);
output(5, 101) <= input(2);
output(5, 102) <= input(3);
output(5, 103) <= input(4);
output(5, 104) <= input(5);
output(5, 105) <= input(6);
output(5, 106) <= input(7);
output(5, 107) <= input(8);
output(5, 108) <= input(9);
output(5, 109) <= input(10);
output(5, 110) <= input(11);
output(5, 111) <= input(12);
output(5, 112) <= input(39);
output(5, 113) <= input(38);
output(5, 114) <= input(36);
output(5, 115) <= input(0);
output(5, 116) <= input(1);
output(5, 117) <= input(2);
output(5, 118) <= input(3);
output(5, 119) <= input(4);
output(5, 120) <= input(5);
output(5, 121) <= input(6);
output(5, 122) <= input(7);
output(5, 123) <= input(8);
output(5, 124) <= input(9);
output(5, 125) <= input(10);
output(5, 126) <= input(11);
output(5, 127) <= input(12);
output(5, 128) <= input(39);
output(5, 129) <= input(38);
output(5, 130) <= input(36);
output(5, 131) <= input(0);
output(5, 132) <= input(1);
output(5, 133) <= input(2);
output(5, 134) <= input(3);
output(5, 135) <= input(4);
output(5, 136) <= input(5);
output(5, 137) <= input(6);
output(5, 138) <= input(7);
output(5, 139) <= input(8);
output(5, 140) <= input(9);
output(5, 141) <= input(10);
output(5, 142) <= input(11);
output(5, 143) <= input(12);
output(5, 144) <= input(39);
output(5, 145) <= input(38);
output(5, 146) <= input(36);
output(5, 147) <= input(0);
output(5, 148) <= input(1);
output(5, 149) <= input(2);
output(5, 150) <= input(3);
output(5, 151) <= input(4);
output(5, 152) <= input(5);
output(5, 153) <= input(6);
output(5, 154) <= input(7);
output(5, 155) <= input(8);
output(5, 156) <= input(9);
output(5, 157) <= input(10);
output(5, 158) <= input(11);
output(5, 159) <= input(12);
output(5, 160) <= input(39);
output(5, 161) <= input(38);
output(5, 162) <= input(36);
output(5, 163) <= input(0);
output(5, 164) <= input(1);
output(5, 165) <= input(2);
output(5, 166) <= input(3);
output(5, 167) <= input(4);
output(5, 168) <= input(5);
output(5, 169) <= input(6);
output(5, 170) <= input(7);
output(5, 171) <= input(8);
output(5, 172) <= input(9);
output(5, 173) <= input(10);
output(5, 174) <= input(11);
output(5, 175) <= input(12);
output(5, 176) <= input(39);
output(5, 177) <= input(38);
output(5, 178) <= input(36);
output(5, 179) <= input(0);
output(5, 180) <= input(1);
output(5, 181) <= input(2);
output(5, 182) <= input(3);
output(5, 183) <= input(4);
output(5, 184) <= input(5);
output(5, 185) <= input(6);
output(5, 186) <= input(7);
output(5, 187) <= input(8);
output(5, 188) <= input(9);
output(5, 189) <= input(10);
output(5, 190) <= input(11);
output(5, 191) <= input(12);
output(5, 192) <= input(39);
output(5, 193) <= input(38);
output(5, 194) <= input(36);
output(5, 195) <= input(0);
output(5, 196) <= input(1);
output(5, 197) <= input(2);
output(5, 198) <= input(3);
output(5, 199) <= input(4);
output(5, 200) <= input(5);
output(5, 201) <= input(6);
output(5, 202) <= input(7);
output(5, 203) <= input(8);
output(5, 204) <= input(9);
output(5, 205) <= input(10);
output(5, 206) <= input(11);
output(5, 207) <= input(12);
output(5, 208) <= input(39);
output(5, 209) <= input(38);
output(5, 210) <= input(36);
output(5, 211) <= input(0);
output(5, 212) <= input(1);
output(5, 213) <= input(2);
output(5, 214) <= input(3);
output(5, 215) <= input(4);
output(5, 216) <= input(5);
output(5, 217) <= input(6);
output(5, 218) <= input(7);
output(5, 219) <= input(8);
output(5, 220) <= input(9);
output(5, 221) <= input(10);
output(5, 222) <= input(11);
output(5, 223) <= input(12);
output(5, 224) <= input(39);
output(5, 225) <= input(38);
output(5, 226) <= input(36);
output(5, 227) <= input(0);
output(5, 228) <= input(1);
output(5, 229) <= input(2);
output(5, 230) <= input(3);
output(5, 231) <= input(4);
output(5, 232) <= input(5);
output(5, 233) <= input(6);
output(5, 234) <= input(7);
output(5, 235) <= input(8);
output(5, 236) <= input(9);
output(5, 237) <= input(10);
output(5, 238) <= input(11);
output(5, 239) <= input(12);
output(5, 240) <= input(39);
output(5, 241) <= input(38);
output(5, 242) <= input(36);
output(5, 243) <= input(0);
output(5, 244) <= input(1);
output(5, 245) <= input(2);
output(5, 246) <= input(3);
output(5, 247) <= input(4);
output(5, 248) <= input(5);
output(5, 249) <= input(6);
output(5, 250) <= input(7);
output(5, 251) <= input(8);
output(5, 252) <= input(9);
output(5, 253) <= input(10);
output(5, 254) <= input(11);
output(5, 255) <= input(12);
output(6, 0) <= input(40);
output(6, 1) <= input(41);
output(6, 2) <= input(37);
output(6, 3) <= input(35);
output(6, 4) <= input(16);
output(6, 5) <= input(17);
output(6, 6) <= input(18);
output(6, 7) <= input(19);
output(6, 8) <= input(20);
output(6, 9) <= input(21);
output(6, 10) <= input(22);
output(6, 11) <= input(23);
output(6, 12) <= input(24);
output(6, 13) <= input(25);
output(6, 14) <= input(26);
output(6, 15) <= input(27);
output(6, 16) <= input(40);
output(6, 17) <= input(41);
output(6, 18) <= input(37);
output(6, 19) <= input(35);
output(6, 20) <= input(16);
output(6, 21) <= input(17);
output(6, 22) <= input(18);
output(6, 23) <= input(19);
output(6, 24) <= input(20);
output(6, 25) <= input(21);
output(6, 26) <= input(22);
output(6, 27) <= input(23);
output(6, 28) <= input(24);
output(6, 29) <= input(25);
output(6, 30) <= input(26);
output(6, 31) <= input(27);
output(6, 32) <= input(40);
output(6, 33) <= input(41);
output(6, 34) <= input(37);
output(6, 35) <= input(35);
output(6, 36) <= input(16);
output(6, 37) <= input(17);
output(6, 38) <= input(18);
output(6, 39) <= input(19);
output(6, 40) <= input(20);
output(6, 41) <= input(21);
output(6, 42) <= input(22);
output(6, 43) <= input(23);
output(6, 44) <= input(24);
output(6, 45) <= input(25);
output(6, 46) <= input(26);
output(6, 47) <= input(27);
output(6, 48) <= input(40);
output(6, 49) <= input(41);
output(6, 50) <= input(37);
output(6, 51) <= input(35);
output(6, 52) <= input(16);
output(6, 53) <= input(17);
output(6, 54) <= input(18);
output(6, 55) <= input(19);
output(6, 56) <= input(20);
output(6, 57) <= input(21);
output(6, 58) <= input(22);
output(6, 59) <= input(23);
output(6, 60) <= input(24);
output(6, 61) <= input(25);
output(6, 62) <= input(26);
output(6, 63) <= input(27);
output(6, 64) <= input(40);
output(6, 65) <= input(41);
output(6, 66) <= input(37);
output(6, 67) <= input(35);
output(6, 68) <= input(16);
output(6, 69) <= input(17);
output(6, 70) <= input(18);
output(6, 71) <= input(19);
output(6, 72) <= input(20);
output(6, 73) <= input(21);
output(6, 74) <= input(22);
output(6, 75) <= input(23);
output(6, 76) <= input(24);
output(6, 77) <= input(25);
output(6, 78) <= input(26);
output(6, 79) <= input(27);
output(6, 80) <= input(40);
output(6, 81) <= input(41);
output(6, 82) <= input(37);
output(6, 83) <= input(35);
output(6, 84) <= input(16);
output(6, 85) <= input(17);
output(6, 86) <= input(18);
output(6, 87) <= input(19);
output(6, 88) <= input(20);
output(6, 89) <= input(21);
output(6, 90) <= input(22);
output(6, 91) <= input(23);
output(6, 92) <= input(24);
output(6, 93) <= input(25);
output(6, 94) <= input(26);
output(6, 95) <= input(27);
output(6, 96) <= input(40);
output(6, 97) <= input(41);
output(6, 98) <= input(37);
output(6, 99) <= input(35);
output(6, 100) <= input(16);
output(6, 101) <= input(17);
output(6, 102) <= input(18);
output(6, 103) <= input(19);
output(6, 104) <= input(20);
output(6, 105) <= input(21);
output(6, 106) <= input(22);
output(6, 107) <= input(23);
output(6, 108) <= input(24);
output(6, 109) <= input(25);
output(6, 110) <= input(26);
output(6, 111) <= input(27);
output(6, 112) <= input(40);
output(6, 113) <= input(41);
output(6, 114) <= input(37);
output(6, 115) <= input(35);
output(6, 116) <= input(16);
output(6, 117) <= input(17);
output(6, 118) <= input(18);
output(6, 119) <= input(19);
output(6, 120) <= input(20);
output(6, 121) <= input(21);
output(6, 122) <= input(22);
output(6, 123) <= input(23);
output(6, 124) <= input(24);
output(6, 125) <= input(25);
output(6, 126) <= input(26);
output(6, 127) <= input(27);
output(6, 128) <= input(42);
output(6, 129) <= input(39);
output(6, 130) <= input(38);
output(6, 131) <= input(36);
output(6, 132) <= input(0);
output(6, 133) <= input(1);
output(6, 134) <= input(2);
output(6, 135) <= input(3);
output(6, 136) <= input(4);
output(6, 137) <= input(5);
output(6, 138) <= input(6);
output(6, 139) <= input(7);
output(6, 140) <= input(8);
output(6, 141) <= input(9);
output(6, 142) <= input(10);
output(6, 143) <= input(11);
output(6, 144) <= input(42);
output(6, 145) <= input(39);
output(6, 146) <= input(38);
output(6, 147) <= input(36);
output(6, 148) <= input(0);
output(6, 149) <= input(1);
output(6, 150) <= input(2);
output(6, 151) <= input(3);
output(6, 152) <= input(4);
output(6, 153) <= input(5);
output(6, 154) <= input(6);
output(6, 155) <= input(7);
output(6, 156) <= input(8);
output(6, 157) <= input(9);
output(6, 158) <= input(10);
output(6, 159) <= input(11);
output(6, 160) <= input(42);
output(6, 161) <= input(39);
output(6, 162) <= input(38);
output(6, 163) <= input(36);
output(6, 164) <= input(0);
output(6, 165) <= input(1);
output(6, 166) <= input(2);
output(6, 167) <= input(3);
output(6, 168) <= input(4);
output(6, 169) <= input(5);
output(6, 170) <= input(6);
output(6, 171) <= input(7);
output(6, 172) <= input(8);
output(6, 173) <= input(9);
output(6, 174) <= input(10);
output(6, 175) <= input(11);
output(6, 176) <= input(42);
output(6, 177) <= input(39);
output(6, 178) <= input(38);
output(6, 179) <= input(36);
output(6, 180) <= input(0);
output(6, 181) <= input(1);
output(6, 182) <= input(2);
output(6, 183) <= input(3);
output(6, 184) <= input(4);
output(6, 185) <= input(5);
output(6, 186) <= input(6);
output(6, 187) <= input(7);
output(6, 188) <= input(8);
output(6, 189) <= input(9);
output(6, 190) <= input(10);
output(6, 191) <= input(11);
output(6, 192) <= input(42);
output(6, 193) <= input(39);
output(6, 194) <= input(38);
output(6, 195) <= input(36);
output(6, 196) <= input(0);
output(6, 197) <= input(1);
output(6, 198) <= input(2);
output(6, 199) <= input(3);
output(6, 200) <= input(4);
output(6, 201) <= input(5);
output(6, 202) <= input(6);
output(6, 203) <= input(7);
output(6, 204) <= input(8);
output(6, 205) <= input(9);
output(6, 206) <= input(10);
output(6, 207) <= input(11);
output(6, 208) <= input(42);
output(6, 209) <= input(39);
output(6, 210) <= input(38);
output(6, 211) <= input(36);
output(6, 212) <= input(0);
output(6, 213) <= input(1);
output(6, 214) <= input(2);
output(6, 215) <= input(3);
output(6, 216) <= input(4);
output(6, 217) <= input(5);
output(6, 218) <= input(6);
output(6, 219) <= input(7);
output(6, 220) <= input(8);
output(6, 221) <= input(9);
output(6, 222) <= input(10);
output(6, 223) <= input(11);
output(6, 224) <= input(42);
output(6, 225) <= input(39);
output(6, 226) <= input(38);
output(6, 227) <= input(36);
output(6, 228) <= input(0);
output(6, 229) <= input(1);
output(6, 230) <= input(2);
output(6, 231) <= input(3);
output(6, 232) <= input(4);
output(6, 233) <= input(5);
output(6, 234) <= input(6);
output(6, 235) <= input(7);
output(6, 236) <= input(8);
output(6, 237) <= input(9);
output(6, 238) <= input(10);
output(6, 239) <= input(11);
output(6, 240) <= input(42);
output(6, 241) <= input(39);
output(6, 242) <= input(38);
output(6, 243) <= input(36);
output(6, 244) <= input(0);
output(6, 245) <= input(1);
output(6, 246) <= input(2);
output(6, 247) <= input(3);
output(6, 248) <= input(4);
output(6, 249) <= input(5);
output(6, 250) <= input(6);
output(6, 251) <= input(7);
output(6, 252) <= input(8);
output(6, 253) <= input(9);
output(6, 254) <= input(10);
output(6, 255) <= input(11);
output(7, 0) <= input(42);
output(7, 1) <= input(39);
output(7, 2) <= input(38);
output(7, 3) <= input(36);
output(7, 4) <= input(0);
output(7, 5) <= input(1);
output(7, 6) <= input(2);
output(7, 7) <= input(3);
output(7, 8) <= input(4);
output(7, 9) <= input(5);
output(7, 10) <= input(6);
output(7, 11) <= input(7);
output(7, 12) <= input(8);
output(7, 13) <= input(9);
output(7, 14) <= input(10);
output(7, 15) <= input(11);
output(7, 16) <= input(42);
output(7, 17) <= input(39);
output(7, 18) <= input(38);
output(7, 19) <= input(36);
output(7, 20) <= input(0);
output(7, 21) <= input(1);
output(7, 22) <= input(2);
output(7, 23) <= input(3);
output(7, 24) <= input(4);
output(7, 25) <= input(5);
output(7, 26) <= input(6);
output(7, 27) <= input(7);
output(7, 28) <= input(8);
output(7, 29) <= input(9);
output(7, 30) <= input(10);
output(7, 31) <= input(11);
output(7, 32) <= input(42);
output(7, 33) <= input(39);
output(7, 34) <= input(38);
output(7, 35) <= input(36);
output(7, 36) <= input(0);
output(7, 37) <= input(1);
output(7, 38) <= input(2);
output(7, 39) <= input(3);
output(7, 40) <= input(4);
output(7, 41) <= input(5);
output(7, 42) <= input(6);
output(7, 43) <= input(7);
output(7, 44) <= input(8);
output(7, 45) <= input(9);
output(7, 46) <= input(10);
output(7, 47) <= input(11);
output(7, 48) <= input(42);
output(7, 49) <= input(39);
output(7, 50) <= input(38);
output(7, 51) <= input(36);
output(7, 52) <= input(0);
output(7, 53) <= input(1);
output(7, 54) <= input(2);
output(7, 55) <= input(3);
output(7, 56) <= input(4);
output(7, 57) <= input(5);
output(7, 58) <= input(6);
output(7, 59) <= input(7);
output(7, 60) <= input(8);
output(7, 61) <= input(9);
output(7, 62) <= input(10);
output(7, 63) <= input(11);
output(7, 64) <= input(42);
output(7, 65) <= input(39);
output(7, 66) <= input(38);
output(7, 67) <= input(36);
output(7, 68) <= input(0);
output(7, 69) <= input(1);
output(7, 70) <= input(2);
output(7, 71) <= input(3);
output(7, 72) <= input(4);
output(7, 73) <= input(5);
output(7, 74) <= input(6);
output(7, 75) <= input(7);
output(7, 76) <= input(8);
output(7, 77) <= input(9);
output(7, 78) <= input(10);
output(7, 79) <= input(11);
output(7, 80) <= input(43);
output(7, 81) <= input(40);
output(7, 82) <= input(41);
output(7, 83) <= input(37);
output(7, 84) <= input(35);
output(7, 85) <= input(16);
output(7, 86) <= input(17);
output(7, 87) <= input(18);
output(7, 88) <= input(19);
output(7, 89) <= input(20);
output(7, 90) <= input(21);
output(7, 91) <= input(22);
output(7, 92) <= input(23);
output(7, 93) <= input(24);
output(7, 94) <= input(25);
output(7, 95) <= input(26);
output(7, 96) <= input(43);
output(7, 97) <= input(40);
output(7, 98) <= input(41);
output(7, 99) <= input(37);
output(7, 100) <= input(35);
output(7, 101) <= input(16);
output(7, 102) <= input(17);
output(7, 103) <= input(18);
output(7, 104) <= input(19);
output(7, 105) <= input(20);
output(7, 106) <= input(21);
output(7, 107) <= input(22);
output(7, 108) <= input(23);
output(7, 109) <= input(24);
output(7, 110) <= input(25);
output(7, 111) <= input(26);
output(7, 112) <= input(43);
output(7, 113) <= input(40);
output(7, 114) <= input(41);
output(7, 115) <= input(37);
output(7, 116) <= input(35);
output(7, 117) <= input(16);
output(7, 118) <= input(17);
output(7, 119) <= input(18);
output(7, 120) <= input(19);
output(7, 121) <= input(20);
output(7, 122) <= input(21);
output(7, 123) <= input(22);
output(7, 124) <= input(23);
output(7, 125) <= input(24);
output(7, 126) <= input(25);
output(7, 127) <= input(26);
output(7, 128) <= input(43);
output(7, 129) <= input(40);
output(7, 130) <= input(41);
output(7, 131) <= input(37);
output(7, 132) <= input(35);
output(7, 133) <= input(16);
output(7, 134) <= input(17);
output(7, 135) <= input(18);
output(7, 136) <= input(19);
output(7, 137) <= input(20);
output(7, 138) <= input(21);
output(7, 139) <= input(22);
output(7, 140) <= input(23);
output(7, 141) <= input(24);
output(7, 142) <= input(25);
output(7, 143) <= input(26);
output(7, 144) <= input(43);
output(7, 145) <= input(40);
output(7, 146) <= input(41);
output(7, 147) <= input(37);
output(7, 148) <= input(35);
output(7, 149) <= input(16);
output(7, 150) <= input(17);
output(7, 151) <= input(18);
output(7, 152) <= input(19);
output(7, 153) <= input(20);
output(7, 154) <= input(21);
output(7, 155) <= input(22);
output(7, 156) <= input(23);
output(7, 157) <= input(24);
output(7, 158) <= input(25);
output(7, 159) <= input(26);
output(7, 160) <= input(44);
output(7, 161) <= input(42);
output(7, 162) <= input(39);
output(7, 163) <= input(38);
output(7, 164) <= input(36);
output(7, 165) <= input(0);
output(7, 166) <= input(1);
output(7, 167) <= input(2);
output(7, 168) <= input(3);
output(7, 169) <= input(4);
output(7, 170) <= input(5);
output(7, 171) <= input(6);
output(7, 172) <= input(7);
output(7, 173) <= input(8);
output(7, 174) <= input(9);
output(7, 175) <= input(10);
output(7, 176) <= input(44);
output(7, 177) <= input(42);
output(7, 178) <= input(39);
output(7, 179) <= input(38);
output(7, 180) <= input(36);
output(7, 181) <= input(0);
output(7, 182) <= input(1);
output(7, 183) <= input(2);
output(7, 184) <= input(3);
output(7, 185) <= input(4);
output(7, 186) <= input(5);
output(7, 187) <= input(6);
output(7, 188) <= input(7);
output(7, 189) <= input(8);
output(7, 190) <= input(9);
output(7, 191) <= input(10);
output(7, 192) <= input(44);
output(7, 193) <= input(42);
output(7, 194) <= input(39);
output(7, 195) <= input(38);
output(7, 196) <= input(36);
output(7, 197) <= input(0);
output(7, 198) <= input(1);
output(7, 199) <= input(2);
output(7, 200) <= input(3);
output(7, 201) <= input(4);
output(7, 202) <= input(5);
output(7, 203) <= input(6);
output(7, 204) <= input(7);
output(7, 205) <= input(8);
output(7, 206) <= input(9);
output(7, 207) <= input(10);
output(7, 208) <= input(44);
output(7, 209) <= input(42);
output(7, 210) <= input(39);
output(7, 211) <= input(38);
output(7, 212) <= input(36);
output(7, 213) <= input(0);
output(7, 214) <= input(1);
output(7, 215) <= input(2);
output(7, 216) <= input(3);
output(7, 217) <= input(4);
output(7, 218) <= input(5);
output(7, 219) <= input(6);
output(7, 220) <= input(7);
output(7, 221) <= input(8);
output(7, 222) <= input(9);
output(7, 223) <= input(10);
output(7, 224) <= input(44);
output(7, 225) <= input(42);
output(7, 226) <= input(39);
output(7, 227) <= input(38);
output(7, 228) <= input(36);
output(7, 229) <= input(0);
output(7, 230) <= input(1);
output(7, 231) <= input(2);
output(7, 232) <= input(3);
output(7, 233) <= input(4);
output(7, 234) <= input(5);
output(7, 235) <= input(6);
output(7, 236) <= input(7);
output(7, 237) <= input(8);
output(7, 238) <= input(9);
output(7, 239) <= input(10);
output(7, 240) <= input(44);
output(7, 241) <= input(42);
output(7, 242) <= input(39);
output(7, 243) <= input(38);
output(7, 244) <= input(36);
output(7, 245) <= input(0);
output(7, 246) <= input(1);
output(7, 247) <= input(2);
output(7, 248) <= input(3);
output(7, 249) <= input(4);
output(7, 250) <= input(5);
output(7, 251) <= input(6);
output(7, 252) <= input(7);
output(7, 253) <= input(8);
output(7, 254) <= input(9);
output(7, 255) <= input(10);
when "0011" =>
output(0, 0) <= input(0);
output(0, 1) <= input(1);
output(0, 2) <= input(2);
output(0, 3) <= input(3);
output(0, 4) <= input(4);
output(0, 5) <= input(5);
output(0, 6) <= input(6);
output(0, 7) <= input(7);
output(0, 8) <= input(8);
output(0, 9) <= input(9);
output(0, 10) <= input(10);
output(0, 11) <= input(11);
output(0, 12) <= input(12);
output(0, 13) <= input(13);
output(0, 14) <= input(14);
output(0, 15) <= input(15);
output(0, 16) <= input(0);
output(0, 17) <= input(1);
output(0, 18) <= input(2);
output(0, 19) <= input(3);
output(0, 20) <= input(4);
output(0, 21) <= input(5);
output(0, 22) <= input(6);
output(0, 23) <= input(7);
output(0, 24) <= input(8);
output(0, 25) <= input(9);
output(0, 26) <= input(10);
output(0, 27) <= input(11);
output(0, 28) <= input(12);
output(0, 29) <= input(13);
output(0, 30) <= input(14);
output(0, 31) <= input(15);
output(0, 32) <= input(0);
output(0, 33) <= input(1);
output(0, 34) <= input(2);
output(0, 35) <= input(3);
output(0, 36) <= input(4);
output(0, 37) <= input(5);
output(0, 38) <= input(6);
output(0, 39) <= input(7);
output(0, 40) <= input(8);
output(0, 41) <= input(9);
output(0, 42) <= input(10);
output(0, 43) <= input(11);
output(0, 44) <= input(12);
output(0, 45) <= input(13);
output(0, 46) <= input(14);
output(0, 47) <= input(15);
output(0, 48) <= input(0);
output(0, 49) <= input(1);
output(0, 50) <= input(2);
output(0, 51) <= input(3);
output(0, 52) <= input(4);
output(0, 53) <= input(5);
output(0, 54) <= input(6);
output(0, 55) <= input(7);
output(0, 56) <= input(8);
output(0, 57) <= input(9);
output(0, 58) <= input(10);
output(0, 59) <= input(11);
output(0, 60) <= input(12);
output(0, 61) <= input(13);
output(0, 62) <= input(14);
output(0, 63) <= input(15);
output(0, 64) <= input(16);
output(0, 65) <= input(17);
output(0, 66) <= input(18);
output(0, 67) <= input(19);
output(0, 68) <= input(20);
output(0, 69) <= input(21);
output(0, 70) <= input(22);
output(0, 71) <= input(23);
output(0, 72) <= input(24);
output(0, 73) <= input(25);
output(0, 74) <= input(26);
output(0, 75) <= input(27);
output(0, 76) <= input(28);
output(0, 77) <= input(29);
output(0, 78) <= input(30);
output(0, 79) <= input(31);
output(0, 80) <= input(16);
output(0, 81) <= input(17);
output(0, 82) <= input(18);
output(0, 83) <= input(19);
output(0, 84) <= input(20);
output(0, 85) <= input(21);
output(0, 86) <= input(22);
output(0, 87) <= input(23);
output(0, 88) <= input(24);
output(0, 89) <= input(25);
output(0, 90) <= input(26);
output(0, 91) <= input(27);
output(0, 92) <= input(28);
output(0, 93) <= input(29);
output(0, 94) <= input(30);
output(0, 95) <= input(31);
output(0, 96) <= input(16);
output(0, 97) <= input(17);
output(0, 98) <= input(18);
output(0, 99) <= input(19);
output(0, 100) <= input(20);
output(0, 101) <= input(21);
output(0, 102) <= input(22);
output(0, 103) <= input(23);
output(0, 104) <= input(24);
output(0, 105) <= input(25);
output(0, 106) <= input(26);
output(0, 107) <= input(27);
output(0, 108) <= input(28);
output(0, 109) <= input(29);
output(0, 110) <= input(30);
output(0, 111) <= input(31);
output(0, 112) <= input(16);
output(0, 113) <= input(17);
output(0, 114) <= input(18);
output(0, 115) <= input(19);
output(0, 116) <= input(20);
output(0, 117) <= input(21);
output(0, 118) <= input(22);
output(0, 119) <= input(23);
output(0, 120) <= input(24);
output(0, 121) <= input(25);
output(0, 122) <= input(26);
output(0, 123) <= input(27);
output(0, 124) <= input(28);
output(0, 125) <= input(29);
output(0, 126) <= input(30);
output(0, 127) <= input(31);
output(0, 128) <= input(32);
output(0, 129) <= input(0);
output(0, 130) <= input(1);
output(0, 131) <= input(2);
output(0, 132) <= input(3);
output(0, 133) <= input(4);
output(0, 134) <= input(5);
output(0, 135) <= input(6);
output(0, 136) <= input(7);
output(0, 137) <= input(8);
output(0, 138) <= input(9);
output(0, 139) <= input(10);
output(0, 140) <= input(11);
output(0, 141) <= input(12);
output(0, 142) <= input(13);
output(0, 143) <= input(14);
output(0, 144) <= input(32);
output(0, 145) <= input(0);
output(0, 146) <= input(1);
output(0, 147) <= input(2);
output(0, 148) <= input(3);
output(0, 149) <= input(4);
output(0, 150) <= input(5);
output(0, 151) <= input(6);
output(0, 152) <= input(7);
output(0, 153) <= input(8);
output(0, 154) <= input(9);
output(0, 155) <= input(10);
output(0, 156) <= input(11);
output(0, 157) <= input(12);
output(0, 158) <= input(13);
output(0, 159) <= input(14);
output(0, 160) <= input(32);
output(0, 161) <= input(0);
output(0, 162) <= input(1);
output(0, 163) <= input(2);
output(0, 164) <= input(3);
output(0, 165) <= input(4);
output(0, 166) <= input(5);
output(0, 167) <= input(6);
output(0, 168) <= input(7);
output(0, 169) <= input(8);
output(0, 170) <= input(9);
output(0, 171) <= input(10);
output(0, 172) <= input(11);
output(0, 173) <= input(12);
output(0, 174) <= input(13);
output(0, 175) <= input(14);
output(0, 176) <= input(32);
output(0, 177) <= input(0);
output(0, 178) <= input(1);
output(0, 179) <= input(2);
output(0, 180) <= input(3);
output(0, 181) <= input(4);
output(0, 182) <= input(5);
output(0, 183) <= input(6);
output(0, 184) <= input(7);
output(0, 185) <= input(8);
output(0, 186) <= input(9);
output(0, 187) <= input(10);
output(0, 188) <= input(11);
output(0, 189) <= input(12);
output(0, 190) <= input(13);
output(0, 191) <= input(14);
output(0, 192) <= input(33);
output(0, 193) <= input(16);
output(0, 194) <= input(17);
output(0, 195) <= input(18);
output(0, 196) <= input(19);
output(0, 197) <= input(20);
output(0, 198) <= input(21);
output(0, 199) <= input(22);
output(0, 200) <= input(23);
output(0, 201) <= input(24);
output(0, 202) <= input(25);
output(0, 203) <= input(26);
output(0, 204) <= input(27);
output(0, 205) <= input(28);
output(0, 206) <= input(29);
output(0, 207) <= input(30);
output(0, 208) <= input(33);
output(0, 209) <= input(16);
output(0, 210) <= input(17);
output(0, 211) <= input(18);
output(0, 212) <= input(19);
output(0, 213) <= input(20);
output(0, 214) <= input(21);
output(0, 215) <= input(22);
output(0, 216) <= input(23);
output(0, 217) <= input(24);
output(0, 218) <= input(25);
output(0, 219) <= input(26);
output(0, 220) <= input(27);
output(0, 221) <= input(28);
output(0, 222) <= input(29);
output(0, 223) <= input(30);
output(0, 224) <= input(33);
output(0, 225) <= input(16);
output(0, 226) <= input(17);
output(0, 227) <= input(18);
output(0, 228) <= input(19);
output(0, 229) <= input(20);
output(0, 230) <= input(21);
output(0, 231) <= input(22);
output(0, 232) <= input(23);
output(0, 233) <= input(24);
output(0, 234) <= input(25);
output(0, 235) <= input(26);
output(0, 236) <= input(27);
output(0, 237) <= input(28);
output(0, 238) <= input(29);
output(0, 239) <= input(30);
output(0, 240) <= input(33);
output(0, 241) <= input(16);
output(0, 242) <= input(17);
output(0, 243) <= input(18);
output(0, 244) <= input(19);
output(0, 245) <= input(20);
output(0, 246) <= input(21);
output(0, 247) <= input(22);
output(0, 248) <= input(23);
output(0, 249) <= input(24);
output(0, 250) <= input(25);
output(0, 251) <= input(26);
output(0, 252) <= input(27);
output(0, 253) <= input(28);
output(0, 254) <= input(29);
output(0, 255) <= input(30);
output(1, 0) <= input(32);
output(1, 1) <= input(0);
output(1, 2) <= input(1);
output(1, 3) <= input(2);
output(1, 4) <= input(3);
output(1, 5) <= input(4);
output(1, 6) <= input(5);
output(1, 7) <= input(6);
output(1, 8) <= input(7);
output(1, 9) <= input(8);
output(1, 10) <= input(9);
output(1, 11) <= input(10);
output(1, 12) <= input(11);
output(1, 13) <= input(12);
output(1, 14) <= input(13);
output(1, 15) <= input(14);
output(1, 16) <= input(32);
output(1, 17) <= input(0);
output(1, 18) <= input(1);
output(1, 19) <= input(2);
output(1, 20) <= input(3);
output(1, 21) <= input(4);
output(1, 22) <= input(5);
output(1, 23) <= input(6);
output(1, 24) <= input(7);
output(1, 25) <= input(8);
output(1, 26) <= input(9);
output(1, 27) <= input(10);
output(1, 28) <= input(11);
output(1, 29) <= input(12);
output(1, 30) <= input(13);
output(1, 31) <= input(14);
output(1, 32) <= input(33);
output(1, 33) <= input(16);
output(1, 34) <= input(17);
output(1, 35) <= input(18);
output(1, 36) <= input(19);
output(1, 37) <= input(20);
output(1, 38) <= input(21);
output(1, 39) <= input(22);
output(1, 40) <= input(23);
output(1, 41) <= input(24);
output(1, 42) <= input(25);
output(1, 43) <= input(26);
output(1, 44) <= input(27);
output(1, 45) <= input(28);
output(1, 46) <= input(29);
output(1, 47) <= input(30);
output(1, 48) <= input(33);
output(1, 49) <= input(16);
output(1, 50) <= input(17);
output(1, 51) <= input(18);
output(1, 52) <= input(19);
output(1, 53) <= input(20);
output(1, 54) <= input(21);
output(1, 55) <= input(22);
output(1, 56) <= input(23);
output(1, 57) <= input(24);
output(1, 58) <= input(25);
output(1, 59) <= input(26);
output(1, 60) <= input(27);
output(1, 61) <= input(28);
output(1, 62) <= input(29);
output(1, 63) <= input(30);
output(1, 64) <= input(33);
output(1, 65) <= input(16);
output(1, 66) <= input(17);
output(1, 67) <= input(18);
output(1, 68) <= input(19);
output(1, 69) <= input(20);
output(1, 70) <= input(21);
output(1, 71) <= input(22);
output(1, 72) <= input(23);
output(1, 73) <= input(24);
output(1, 74) <= input(25);
output(1, 75) <= input(26);
output(1, 76) <= input(27);
output(1, 77) <= input(28);
output(1, 78) <= input(29);
output(1, 79) <= input(30);
output(1, 80) <= input(34);
output(1, 81) <= input(32);
output(1, 82) <= input(0);
output(1, 83) <= input(1);
output(1, 84) <= input(2);
output(1, 85) <= input(3);
output(1, 86) <= input(4);
output(1, 87) <= input(5);
output(1, 88) <= input(6);
output(1, 89) <= input(7);
output(1, 90) <= input(8);
output(1, 91) <= input(9);
output(1, 92) <= input(10);
output(1, 93) <= input(11);
output(1, 94) <= input(12);
output(1, 95) <= input(13);
output(1, 96) <= input(34);
output(1, 97) <= input(32);
output(1, 98) <= input(0);
output(1, 99) <= input(1);
output(1, 100) <= input(2);
output(1, 101) <= input(3);
output(1, 102) <= input(4);
output(1, 103) <= input(5);
output(1, 104) <= input(6);
output(1, 105) <= input(7);
output(1, 106) <= input(8);
output(1, 107) <= input(9);
output(1, 108) <= input(10);
output(1, 109) <= input(11);
output(1, 110) <= input(12);
output(1, 111) <= input(13);
output(1, 112) <= input(34);
output(1, 113) <= input(32);
output(1, 114) <= input(0);
output(1, 115) <= input(1);
output(1, 116) <= input(2);
output(1, 117) <= input(3);
output(1, 118) <= input(4);
output(1, 119) <= input(5);
output(1, 120) <= input(6);
output(1, 121) <= input(7);
output(1, 122) <= input(8);
output(1, 123) <= input(9);
output(1, 124) <= input(10);
output(1, 125) <= input(11);
output(1, 126) <= input(12);
output(1, 127) <= input(13);
output(1, 128) <= input(35);
output(1, 129) <= input(33);
output(1, 130) <= input(16);
output(1, 131) <= input(17);
output(1, 132) <= input(18);
output(1, 133) <= input(19);
output(1, 134) <= input(20);
output(1, 135) <= input(21);
output(1, 136) <= input(22);
output(1, 137) <= input(23);
output(1, 138) <= input(24);
output(1, 139) <= input(25);
output(1, 140) <= input(26);
output(1, 141) <= input(27);
output(1, 142) <= input(28);
output(1, 143) <= input(29);
output(1, 144) <= input(35);
output(1, 145) <= input(33);
output(1, 146) <= input(16);
output(1, 147) <= input(17);
output(1, 148) <= input(18);
output(1, 149) <= input(19);
output(1, 150) <= input(20);
output(1, 151) <= input(21);
output(1, 152) <= input(22);
output(1, 153) <= input(23);
output(1, 154) <= input(24);
output(1, 155) <= input(25);
output(1, 156) <= input(26);
output(1, 157) <= input(27);
output(1, 158) <= input(28);
output(1, 159) <= input(29);
output(1, 160) <= input(36);
output(1, 161) <= input(34);
output(1, 162) <= input(32);
output(1, 163) <= input(0);
output(1, 164) <= input(1);
output(1, 165) <= input(2);
output(1, 166) <= input(3);
output(1, 167) <= input(4);
output(1, 168) <= input(5);
output(1, 169) <= input(6);
output(1, 170) <= input(7);
output(1, 171) <= input(8);
output(1, 172) <= input(9);
output(1, 173) <= input(10);
output(1, 174) <= input(11);
output(1, 175) <= input(12);
output(1, 176) <= input(36);
output(1, 177) <= input(34);
output(1, 178) <= input(32);
output(1, 179) <= input(0);
output(1, 180) <= input(1);
output(1, 181) <= input(2);
output(1, 182) <= input(3);
output(1, 183) <= input(4);
output(1, 184) <= input(5);
output(1, 185) <= input(6);
output(1, 186) <= input(7);
output(1, 187) <= input(8);
output(1, 188) <= input(9);
output(1, 189) <= input(10);
output(1, 190) <= input(11);
output(1, 191) <= input(12);
output(1, 192) <= input(36);
output(1, 193) <= input(34);
output(1, 194) <= input(32);
output(1, 195) <= input(0);
output(1, 196) <= input(1);
output(1, 197) <= input(2);
output(1, 198) <= input(3);
output(1, 199) <= input(4);
output(1, 200) <= input(5);
output(1, 201) <= input(6);
output(1, 202) <= input(7);
output(1, 203) <= input(8);
output(1, 204) <= input(9);
output(1, 205) <= input(10);
output(1, 206) <= input(11);
output(1, 207) <= input(12);
output(1, 208) <= input(37);
output(1, 209) <= input(35);
output(1, 210) <= input(33);
output(1, 211) <= input(16);
output(1, 212) <= input(17);
output(1, 213) <= input(18);
output(1, 214) <= input(19);
output(1, 215) <= input(20);
output(1, 216) <= input(21);
output(1, 217) <= input(22);
output(1, 218) <= input(23);
output(1, 219) <= input(24);
output(1, 220) <= input(25);
output(1, 221) <= input(26);
output(1, 222) <= input(27);
output(1, 223) <= input(28);
output(1, 224) <= input(37);
output(1, 225) <= input(35);
output(1, 226) <= input(33);
output(1, 227) <= input(16);
output(1, 228) <= input(17);
output(1, 229) <= input(18);
output(1, 230) <= input(19);
output(1, 231) <= input(20);
output(1, 232) <= input(21);
output(1, 233) <= input(22);
output(1, 234) <= input(23);
output(1, 235) <= input(24);
output(1, 236) <= input(25);
output(1, 237) <= input(26);
output(1, 238) <= input(27);
output(1, 239) <= input(28);
output(1, 240) <= input(37);
output(1, 241) <= input(35);
output(1, 242) <= input(33);
output(1, 243) <= input(16);
output(1, 244) <= input(17);
output(1, 245) <= input(18);
output(1, 246) <= input(19);
output(1, 247) <= input(20);
output(1, 248) <= input(21);
output(1, 249) <= input(22);
output(1, 250) <= input(23);
output(1, 251) <= input(24);
output(1, 252) <= input(25);
output(1, 253) <= input(26);
output(1, 254) <= input(27);
output(1, 255) <= input(28);
output(2, 0) <= input(34);
output(2, 1) <= input(32);
output(2, 2) <= input(0);
output(2, 3) <= input(1);
output(2, 4) <= input(2);
output(2, 5) <= input(3);
output(2, 6) <= input(4);
output(2, 7) <= input(5);
output(2, 8) <= input(6);
output(2, 9) <= input(7);
output(2, 10) <= input(8);
output(2, 11) <= input(9);
output(2, 12) <= input(10);
output(2, 13) <= input(11);
output(2, 14) <= input(12);
output(2, 15) <= input(13);
output(2, 16) <= input(34);
output(2, 17) <= input(32);
output(2, 18) <= input(0);
output(2, 19) <= input(1);
output(2, 20) <= input(2);
output(2, 21) <= input(3);
output(2, 22) <= input(4);
output(2, 23) <= input(5);
output(2, 24) <= input(6);
output(2, 25) <= input(7);
output(2, 26) <= input(8);
output(2, 27) <= input(9);
output(2, 28) <= input(10);
output(2, 29) <= input(11);
output(2, 30) <= input(12);
output(2, 31) <= input(13);
output(2, 32) <= input(35);
output(2, 33) <= input(33);
output(2, 34) <= input(16);
output(2, 35) <= input(17);
output(2, 36) <= input(18);
output(2, 37) <= input(19);
output(2, 38) <= input(20);
output(2, 39) <= input(21);
output(2, 40) <= input(22);
output(2, 41) <= input(23);
output(2, 42) <= input(24);
output(2, 43) <= input(25);
output(2, 44) <= input(26);
output(2, 45) <= input(27);
output(2, 46) <= input(28);
output(2, 47) <= input(29);
output(2, 48) <= input(35);
output(2, 49) <= input(33);
output(2, 50) <= input(16);
output(2, 51) <= input(17);
output(2, 52) <= input(18);
output(2, 53) <= input(19);
output(2, 54) <= input(20);
output(2, 55) <= input(21);
output(2, 56) <= input(22);
output(2, 57) <= input(23);
output(2, 58) <= input(24);
output(2, 59) <= input(25);
output(2, 60) <= input(26);
output(2, 61) <= input(27);
output(2, 62) <= input(28);
output(2, 63) <= input(29);
output(2, 64) <= input(36);
output(2, 65) <= input(34);
output(2, 66) <= input(32);
output(2, 67) <= input(0);
output(2, 68) <= input(1);
output(2, 69) <= input(2);
output(2, 70) <= input(3);
output(2, 71) <= input(4);
output(2, 72) <= input(5);
output(2, 73) <= input(6);
output(2, 74) <= input(7);
output(2, 75) <= input(8);
output(2, 76) <= input(9);
output(2, 77) <= input(10);
output(2, 78) <= input(11);
output(2, 79) <= input(12);
output(2, 80) <= input(36);
output(2, 81) <= input(34);
output(2, 82) <= input(32);
output(2, 83) <= input(0);
output(2, 84) <= input(1);
output(2, 85) <= input(2);
output(2, 86) <= input(3);
output(2, 87) <= input(4);
output(2, 88) <= input(5);
output(2, 89) <= input(6);
output(2, 90) <= input(7);
output(2, 91) <= input(8);
output(2, 92) <= input(9);
output(2, 93) <= input(10);
output(2, 94) <= input(11);
output(2, 95) <= input(12);
output(2, 96) <= input(37);
output(2, 97) <= input(35);
output(2, 98) <= input(33);
output(2, 99) <= input(16);
output(2, 100) <= input(17);
output(2, 101) <= input(18);
output(2, 102) <= input(19);
output(2, 103) <= input(20);
output(2, 104) <= input(21);
output(2, 105) <= input(22);
output(2, 106) <= input(23);
output(2, 107) <= input(24);
output(2, 108) <= input(25);
output(2, 109) <= input(26);
output(2, 110) <= input(27);
output(2, 111) <= input(28);
output(2, 112) <= input(37);
output(2, 113) <= input(35);
output(2, 114) <= input(33);
output(2, 115) <= input(16);
output(2, 116) <= input(17);
output(2, 117) <= input(18);
output(2, 118) <= input(19);
output(2, 119) <= input(20);
output(2, 120) <= input(21);
output(2, 121) <= input(22);
output(2, 122) <= input(23);
output(2, 123) <= input(24);
output(2, 124) <= input(25);
output(2, 125) <= input(26);
output(2, 126) <= input(27);
output(2, 127) <= input(28);
output(2, 128) <= input(38);
output(2, 129) <= input(36);
output(2, 130) <= input(34);
output(2, 131) <= input(32);
output(2, 132) <= input(0);
output(2, 133) <= input(1);
output(2, 134) <= input(2);
output(2, 135) <= input(3);
output(2, 136) <= input(4);
output(2, 137) <= input(5);
output(2, 138) <= input(6);
output(2, 139) <= input(7);
output(2, 140) <= input(8);
output(2, 141) <= input(9);
output(2, 142) <= input(10);
output(2, 143) <= input(11);
output(2, 144) <= input(38);
output(2, 145) <= input(36);
output(2, 146) <= input(34);
output(2, 147) <= input(32);
output(2, 148) <= input(0);
output(2, 149) <= input(1);
output(2, 150) <= input(2);
output(2, 151) <= input(3);
output(2, 152) <= input(4);
output(2, 153) <= input(5);
output(2, 154) <= input(6);
output(2, 155) <= input(7);
output(2, 156) <= input(8);
output(2, 157) <= input(9);
output(2, 158) <= input(10);
output(2, 159) <= input(11);
output(2, 160) <= input(39);
output(2, 161) <= input(37);
output(2, 162) <= input(35);
output(2, 163) <= input(33);
output(2, 164) <= input(16);
output(2, 165) <= input(17);
output(2, 166) <= input(18);
output(2, 167) <= input(19);
output(2, 168) <= input(20);
output(2, 169) <= input(21);
output(2, 170) <= input(22);
output(2, 171) <= input(23);
output(2, 172) <= input(24);
output(2, 173) <= input(25);
output(2, 174) <= input(26);
output(2, 175) <= input(27);
output(2, 176) <= input(39);
output(2, 177) <= input(37);
output(2, 178) <= input(35);
output(2, 179) <= input(33);
output(2, 180) <= input(16);
output(2, 181) <= input(17);
output(2, 182) <= input(18);
output(2, 183) <= input(19);
output(2, 184) <= input(20);
output(2, 185) <= input(21);
output(2, 186) <= input(22);
output(2, 187) <= input(23);
output(2, 188) <= input(24);
output(2, 189) <= input(25);
output(2, 190) <= input(26);
output(2, 191) <= input(27);
output(2, 192) <= input(40);
output(2, 193) <= input(38);
output(2, 194) <= input(36);
output(2, 195) <= input(34);
output(2, 196) <= input(32);
output(2, 197) <= input(0);
output(2, 198) <= input(1);
output(2, 199) <= input(2);
output(2, 200) <= input(3);
output(2, 201) <= input(4);
output(2, 202) <= input(5);
output(2, 203) <= input(6);
output(2, 204) <= input(7);
output(2, 205) <= input(8);
output(2, 206) <= input(9);
output(2, 207) <= input(10);
output(2, 208) <= input(40);
output(2, 209) <= input(38);
output(2, 210) <= input(36);
output(2, 211) <= input(34);
output(2, 212) <= input(32);
output(2, 213) <= input(0);
output(2, 214) <= input(1);
output(2, 215) <= input(2);
output(2, 216) <= input(3);
output(2, 217) <= input(4);
output(2, 218) <= input(5);
output(2, 219) <= input(6);
output(2, 220) <= input(7);
output(2, 221) <= input(8);
output(2, 222) <= input(9);
output(2, 223) <= input(10);
output(2, 224) <= input(41);
output(2, 225) <= input(39);
output(2, 226) <= input(37);
output(2, 227) <= input(35);
output(2, 228) <= input(33);
output(2, 229) <= input(16);
output(2, 230) <= input(17);
output(2, 231) <= input(18);
output(2, 232) <= input(19);
output(2, 233) <= input(20);
output(2, 234) <= input(21);
output(2, 235) <= input(22);
output(2, 236) <= input(23);
output(2, 237) <= input(24);
output(2, 238) <= input(25);
output(2, 239) <= input(26);
output(2, 240) <= input(41);
output(2, 241) <= input(39);
output(2, 242) <= input(37);
output(2, 243) <= input(35);
output(2, 244) <= input(33);
output(2, 245) <= input(16);
output(2, 246) <= input(17);
output(2, 247) <= input(18);
output(2, 248) <= input(19);
output(2, 249) <= input(20);
output(2, 250) <= input(21);
output(2, 251) <= input(22);
output(2, 252) <= input(23);
output(2, 253) <= input(24);
output(2, 254) <= input(25);
output(2, 255) <= input(26);
when "0100" =>
output(0, 0) <= input(0);
output(0, 1) <= input(1);
output(0, 2) <= input(2);
output(0, 3) <= input(3);
output(0, 4) <= input(4);
output(0, 5) <= input(5);
output(0, 6) <= input(6);
output(0, 7) <= input(7);
output(0, 8) <= input(8);
output(0, 9) <= input(9);
output(0, 10) <= input(10);
output(0, 11) <= input(11);
output(0, 12) <= input(12);
output(0, 13) <= input(13);
output(0, 14) <= input(14);
output(0, 15) <= input(15);
output(0, 16) <= input(16);
output(0, 17) <= input(17);
output(0, 18) <= input(18);
output(0, 19) <= input(19);
output(0, 20) <= input(20);
output(0, 21) <= input(21);
output(0, 22) <= input(22);
output(0, 23) <= input(23);
output(0, 24) <= input(24);
output(0, 25) <= input(25);
output(0, 26) <= input(26);
output(0, 27) <= input(27);
output(0, 28) <= input(28);
output(0, 29) <= input(29);
output(0, 30) <= input(30);
output(0, 31) <= input(31);
output(0, 32) <= input(16);
output(0, 33) <= input(17);
output(0, 34) <= input(18);
output(0, 35) <= input(19);
output(0, 36) <= input(20);
output(0, 37) <= input(21);
output(0, 38) <= input(22);
output(0, 39) <= input(23);
output(0, 40) <= input(24);
output(0, 41) <= input(25);
output(0, 42) <= input(26);
output(0, 43) <= input(27);
output(0, 44) <= input(28);
output(0, 45) <= input(29);
output(0, 46) <= input(30);
output(0, 47) <= input(31);
output(0, 48) <= input(32);
output(0, 49) <= input(0);
output(0, 50) <= input(1);
output(0, 51) <= input(2);
output(0, 52) <= input(3);
output(0, 53) <= input(4);
output(0, 54) <= input(5);
output(0, 55) <= input(6);
output(0, 56) <= input(7);
output(0, 57) <= input(8);
output(0, 58) <= input(9);
output(0, 59) <= input(10);
output(0, 60) <= input(11);
output(0, 61) <= input(12);
output(0, 62) <= input(13);
output(0, 63) <= input(14);
output(0, 64) <= input(33);
output(0, 65) <= input(16);
output(0, 66) <= input(17);
output(0, 67) <= input(18);
output(0, 68) <= input(19);
output(0, 69) <= input(20);
output(0, 70) <= input(21);
output(0, 71) <= input(22);
output(0, 72) <= input(23);
output(0, 73) <= input(24);
output(0, 74) <= input(25);
output(0, 75) <= input(26);
output(0, 76) <= input(27);
output(0, 77) <= input(28);
output(0, 78) <= input(29);
output(0, 79) <= input(30);
output(0, 80) <= input(33);
output(0, 81) <= input(16);
output(0, 82) <= input(17);
output(0, 83) <= input(18);
output(0, 84) <= input(19);
output(0, 85) <= input(20);
output(0, 86) <= input(21);
output(0, 87) <= input(22);
output(0, 88) <= input(23);
output(0, 89) <= input(24);
output(0, 90) <= input(25);
output(0, 91) <= input(26);
output(0, 92) <= input(27);
output(0, 93) <= input(28);
output(0, 94) <= input(29);
output(0, 95) <= input(30);
output(0, 96) <= input(34);
output(0, 97) <= input(32);
output(0, 98) <= input(0);
output(0, 99) <= input(1);
output(0, 100) <= input(2);
output(0, 101) <= input(3);
output(0, 102) <= input(4);
output(0, 103) <= input(5);
output(0, 104) <= input(6);
output(0, 105) <= input(7);
output(0, 106) <= input(8);
output(0, 107) <= input(9);
output(0, 108) <= input(10);
output(0, 109) <= input(11);
output(0, 110) <= input(12);
output(0, 111) <= input(13);
output(0, 112) <= input(34);
output(0, 113) <= input(32);
output(0, 114) <= input(0);
output(0, 115) <= input(1);
output(0, 116) <= input(2);
output(0, 117) <= input(3);
output(0, 118) <= input(4);
output(0, 119) <= input(5);
output(0, 120) <= input(6);
output(0, 121) <= input(7);
output(0, 122) <= input(8);
output(0, 123) <= input(9);
output(0, 124) <= input(10);
output(0, 125) <= input(11);
output(0, 126) <= input(12);
output(0, 127) <= input(13);
output(0, 128) <= input(35);
output(0, 129) <= input(33);
output(0, 130) <= input(16);
output(0, 131) <= input(17);
output(0, 132) <= input(18);
output(0, 133) <= input(19);
output(0, 134) <= input(20);
output(0, 135) <= input(21);
output(0, 136) <= input(22);
output(0, 137) <= input(23);
output(0, 138) <= input(24);
output(0, 139) <= input(25);
output(0, 140) <= input(26);
output(0, 141) <= input(27);
output(0, 142) <= input(28);
output(0, 143) <= input(29);
output(0, 144) <= input(36);
output(0, 145) <= input(34);
output(0, 146) <= input(32);
output(0, 147) <= input(0);
output(0, 148) <= input(1);
output(0, 149) <= input(2);
output(0, 150) <= input(3);
output(0, 151) <= input(4);
output(0, 152) <= input(5);
output(0, 153) <= input(6);
output(0, 154) <= input(7);
output(0, 155) <= input(8);
output(0, 156) <= input(9);
output(0, 157) <= input(10);
output(0, 158) <= input(11);
output(0, 159) <= input(12);
output(0, 160) <= input(36);
output(0, 161) <= input(34);
output(0, 162) <= input(32);
output(0, 163) <= input(0);
output(0, 164) <= input(1);
output(0, 165) <= input(2);
output(0, 166) <= input(3);
output(0, 167) <= input(4);
output(0, 168) <= input(5);
output(0, 169) <= input(6);
output(0, 170) <= input(7);
output(0, 171) <= input(8);
output(0, 172) <= input(9);
output(0, 173) <= input(10);
output(0, 174) <= input(11);
output(0, 175) <= input(12);
output(0, 176) <= input(37);
output(0, 177) <= input(35);
output(0, 178) <= input(33);
output(0, 179) <= input(16);
output(0, 180) <= input(17);
output(0, 181) <= input(18);
output(0, 182) <= input(19);
output(0, 183) <= input(20);
output(0, 184) <= input(21);
output(0, 185) <= input(22);
output(0, 186) <= input(23);
output(0, 187) <= input(24);
output(0, 188) <= input(25);
output(0, 189) <= input(26);
output(0, 190) <= input(27);
output(0, 191) <= input(28);
output(0, 192) <= input(38);
output(0, 193) <= input(36);
output(0, 194) <= input(34);
output(0, 195) <= input(32);
output(0, 196) <= input(0);
output(0, 197) <= input(1);
output(0, 198) <= input(2);
output(0, 199) <= input(3);
output(0, 200) <= input(4);
output(0, 201) <= input(5);
output(0, 202) <= input(6);
output(0, 203) <= input(7);
output(0, 204) <= input(8);
output(0, 205) <= input(9);
output(0, 206) <= input(10);
output(0, 207) <= input(11);
output(0, 208) <= input(38);
output(0, 209) <= input(36);
output(0, 210) <= input(34);
output(0, 211) <= input(32);
output(0, 212) <= input(0);
output(0, 213) <= input(1);
output(0, 214) <= input(2);
output(0, 215) <= input(3);
output(0, 216) <= input(4);
output(0, 217) <= input(5);
output(0, 218) <= input(6);
output(0, 219) <= input(7);
output(0, 220) <= input(8);
output(0, 221) <= input(9);
output(0, 222) <= input(10);
output(0, 223) <= input(11);
output(0, 224) <= input(39);
output(0, 225) <= input(37);
output(0, 226) <= input(35);
output(0, 227) <= input(33);
output(0, 228) <= input(16);
output(0, 229) <= input(17);
output(0, 230) <= input(18);
output(0, 231) <= input(19);
output(0, 232) <= input(20);
output(0, 233) <= input(21);
output(0, 234) <= input(22);
output(0, 235) <= input(23);
output(0, 236) <= input(24);
output(0, 237) <= input(25);
output(0, 238) <= input(26);
output(0, 239) <= input(27);
output(0, 240) <= input(39);
output(0, 241) <= input(37);
output(0, 242) <= input(35);
output(0, 243) <= input(33);
output(0, 244) <= input(16);
output(0, 245) <= input(17);
output(0, 246) <= input(18);
output(0, 247) <= input(19);
output(0, 248) <= input(20);
output(0, 249) <= input(21);
output(0, 250) <= input(22);
output(0, 251) <= input(23);
output(0, 252) <= input(24);
output(0, 253) <= input(25);
output(0, 254) <= input(26);
output(0, 255) <= input(27);
output(1, 0) <= input(32);
output(1, 1) <= input(0);
output(1, 2) <= input(1);
output(1, 3) <= input(2);
output(1, 4) <= input(3);
output(1, 5) <= input(4);
output(1, 6) <= input(5);
output(1, 7) <= input(6);
output(1, 8) <= input(7);
output(1, 9) <= input(8);
output(1, 10) <= input(9);
output(1, 11) <= input(10);
output(1, 12) <= input(11);
output(1, 13) <= input(12);
output(1, 14) <= input(13);
output(1, 15) <= input(14);
output(1, 16) <= input(33);
output(1, 17) <= input(16);
output(1, 18) <= input(17);
output(1, 19) <= input(18);
output(1, 20) <= input(19);
output(1, 21) <= input(20);
output(1, 22) <= input(21);
output(1, 23) <= input(22);
output(1, 24) <= input(23);
output(1, 25) <= input(24);
output(1, 26) <= input(25);
output(1, 27) <= input(26);
output(1, 28) <= input(27);
output(1, 29) <= input(28);
output(1, 30) <= input(29);
output(1, 31) <= input(30);
output(1, 32) <= input(34);
output(1, 33) <= input(32);
output(1, 34) <= input(0);
output(1, 35) <= input(1);
output(1, 36) <= input(2);
output(1, 37) <= input(3);
output(1, 38) <= input(4);
output(1, 39) <= input(5);
output(1, 40) <= input(6);
output(1, 41) <= input(7);
output(1, 42) <= input(8);
output(1, 43) <= input(9);
output(1, 44) <= input(10);
output(1, 45) <= input(11);
output(1, 46) <= input(12);
output(1, 47) <= input(13);
output(1, 48) <= input(34);
output(1, 49) <= input(32);
output(1, 50) <= input(0);
output(1, 51) <= input(1);
output(1, 52) <= input(2);
output(1, 53) <= input(3);
output(1, 54) <= input(4);
output(1, 55) <= input(5);
output(1, 56) <= input(6);
output(1, 57) <= input(7);
output(1, 58) <= input(8);
output(1, 59) <= input(9);
output(1, 60) <= input(10);
output(1, 61) <= input(11);
output(1, 62) <= input(12);
output(1, 63) <= input(13);
output(1, 64) <= input(35);
output(1, 65) <= input(33);
output(1, 66) <= input(16);
output(1, 67) <= input(17);
output(1, 68) <= input(18);
output(1, 69) <= input(19);
output(1, 70) <= input(20);
output(1, 71) <= input(21);
output(1, 72) <= input(22);
output(1, 73) <= input(23);
output(1, 74) <= input(24);
output(1, 75) <= input(25);
output(1, 76) <= input(26);
output(1, 77) <= input(27);
output(1, 78) <= input(28);
output(1, 79) <= input(29);
output(1, 80) <= input(36);
output(1, 81) <= input(34);
output(1, 82) <= input(32);
output(1, 83) <= input(0);
output(1, 84) <= input(1);
output(1, 85) <= input(2);
output(1, 86) <= input(3);
output(1, 87) <= input(4);
output(1, 88) <= input(5);
output(1, 89) <= input(6);
output(1, 90) <= input(7);
output(1, 91) <= input(8);
output(1, 92) <= input(9);
output(1, 93) <= input(10);
output(1, 94) <= input(11);
output(1, 95) <= input(12);
output(1, 96) <= input(37);
output(1, 97) <= input(35);
output(1, 98) <= input(33);
output(1, 99) <= input(16);
output(1, 100) <= input(17);
output(1, 101) <= input(18);
output(1, 102) <= input(19);
output(1, 103) <= input(20);
output(1, 104) <= input(21);
output(1, 105) <= input(22);
output(1, 106) <= input(23);
output(1, 107) <= input(24);
output(1, 108) <= input(25);
output(1, 109) <= input(26);
output(1, 110) <= input(27);
output(1, 111) <= input(28);
output(1, 112) <= input(37);
output(1, 113) <= input(35);
output(1, 114) <= input(33);
output(1, 115) <= input(16);
output(1, 116) <= input(17);
output(1, 117) <= input(18);
output(1, 118) <= input(19);
output(1, 119) <= input(20);
output(1, 120) <= input(21);
output(1, 121) <= input(22);
output(1, 122) <= input(23);
output(1, 123) <= input(24);
output(1, 124) <= input(25);
output(1, 125) <= input(26);
output(1, 126) <= input(27);
output(1, 127) <= input(28);
output(1, 128) <= input(38);
output(1, 129) <= input(36);
output(1, 130) <= input(34);
output(1, 131) <= input(32);
output(1, 132) <= input(0);
output(1, 133) <= input(1);
output(1, 134) <= input(2);
output(1, 135) <= input(3);
output(1, 136) <= input(4);
output(1, 137) <= input(5);
output(1, 138) <= input(6);
output(1, 139) <= input(7);
output(1, 140) <= input(8);
output(1, 141) <= input(9);
output(1, 142) <= input(10);
output(1, 143) <= input(11);
output(1, 144) <= input(39);
output(1, 145) <= input(37);
output(1, 146) <= input(35);
output(1, 147) <= input(33);
output(1, 148) <= input(16);
output(1, 149) <= input(17);
output(1, 150) <= input(18);
output(1, 151) <= input(19);
output(1, 152) <= input(20);
output(1, 153) <= input(21);
output(1, 154) <= input(22);
output(1, 155) <= input(23);
output(1, 156) <= input(24);
output(1, 157) <= input(25);
output(1, 158) <= input(26);
output(1, 159) <= input(27);
output(1, 160) <= input(40);
output(1, 161) <= input(38);
output(1, 162) <= input(36);
output(1, 163) <= input(34);
output(1, 164) <= input(32);
output(1, 165) <= input(0);
output(1, 166) <= input(1);
output(1, 167) <= input(2);
output(1, 168) <= input(3);
output(1, 169) <= input(4);
output(1, 170) <= input(5);
output(1, 171) <= input(6);
output(1, 172) <= input(7);
output(1, 173) <= input(8);
output(1, 174) <= input(9);
output(1, 175) <= input(10);
output(1, 176) <= input(40);
output(1, 177) <= input(38);
output(1, 178) <= input(36);
output(1, 179) <= input(34);
output(1, 180) <= input(32);
output(1, 181) <= input(0);
output(1, 182) <= input(1);
output(1, 183) <= input(2);
output(1, 184) <= input(3);
output(1, 185) <= input(4);
output(1, 186) <= input(5);
output(1, 187) <= input(6);
output(1, 188) <= input(7);
output(1, 189) <= input(8);
output(1, 190) <= input(9);
output(1, 191) <= input(10);
output(1, 192) <= input(41);
output(1, 193) <= input(39);
output(1, 194) <= input(37);
output(1, 195) <= input(35);
output(1, 196) <= input(33);
output(1, 197) <= input(16);
output(1, 198) <= input(17);
output(1, 199) <= input(18);
output(1, 200) <= input(19);
output(1, 201) <= input(20);
output(1, 202) <= input(21);
output(1, 203) <= input(22);
output(1, 204) <= input(23);
output(1, 205) <= input(24);
output(1, 206) <= input(25);
output(1, 207) <= input(26);
output(1, 208) <= input(42);
output(1, 209) <= input(40);
output(1, 210) <= input(38);
output(1, 211) <= input(36);
output(1, 212) <= input(34);
output(1, 213) <= input(32);
output(1, 214) <= input(0);
output(1, 215) <= input(1);
output(1, 216) <= input(2);
output(1, 217) <= input(3);
output(1, 218) <= input(4);
output(1, 219) <= input(5);
output(1, 220) <= input(6);
output(1, 221) <= input(7);
output(1, 222) <= input(8);
output(1, 223) <= input(9);
output(1, 224) <= input(43);
output(1, 225) <= input(41);
output(1, 226) <= input(39);
output(1, 227) <= input(37);
output(1, 228) <= input(35);
output(1, 229) <= input(33);
output(1, 230) <= input(16);
output(1, 231) <= input(17);
output(1, 232) <= input(18);
output(1, 233) <= input(19);
output(1, 234) <= input(20);
output(1, 235) <= input(21);
output(1, 236) <= input(22);
output(1, 237) <= input(23);
output(1, 238) <= input(24);
output(1, 239) <= input(25);
output(1, 240) <= input(43);
output(1, 241) <= input(41);
output(1, 242) <= input(39);
output(1, 243) <= input(37);
output(1, 244) <= input(35);
output(1, 245) <= input(33);
output(1, 246) <= input(16);
output(1, 247) <= input(17);
output(1, 248) <= input(18);
output(1, 249) <= input(19);
output(1, 250) <= input(20);
output(1, 251) <= input(21);
output(1, 252) <= input(22);
output(1, 253) <= input(23);
output(1, 254) <= input(24);
output(1, 255) <= input(25);
output(2, 0) <= input(34);
output(2, 1) <= input(32);
output(2, 2) <= input(0);
output(2, 3) <= input(1);
output(2, 4) <= input(2);
output(2, 5) <= input(3);
output(2, 6) <= input(4);
output(2, 7) <= input(5);
output(2, 8) <= input(6);
output(2, 9) <= input(7);
output(2, 10) <= input(8);
output(2, 11) <= input(9);
output(2, 12) <= input(10);
output(2, 13) <= input(11);
output(2, 14) <= input(12);
output(2, 15) <= input(13);
output(2, 16) <= input(35);
output(2, 17) <= input(33);
output(2, 18) <= input(16);
output(2, 19) <= input(17);
output(2, 20) <= input(18);
output(2, 21) <= input(19);
output(2, 22) <= input(20);
output(2, 23) <= input(21);
output(2, 24) <= input(22);
output(2, 25) <= input(23);
output(2, 26) <= input(24);
output(2, 27) <= input(25);
output(2, 28) <= input(26);
output(2, 29) <= input(27);
output(2, 30) <= input(28);
output(2, 31) <= input(29);
output(2, 32) <= input(36);
output(2, 33) <= input(34);
output(2, 34) <= input(32);
output(2, 35) <= input(0);
output(2, 36) <= input(1);
output(2, 37) <= input(2);
output(2, 38) <= input(3);
output(2, 39) <= input(4);
output(2, 40) <= input(5);
output(2, 41) <= input(6);
output(2, 42) <= input(7);
output(2, 43) <= input(8);
output(2, 44) <= input(9);
output(2, 45) <= input(10);
output(2, 46) <= input(11);
output(2, 47) <= input(12);
output(2, 48) <= input(37);
output(2, 49) <= input(35);
output(2, 50) <= input(33);
output(2, 51) <= input(16);
output(2, 52) <= input(17);
output(2, 53) <= input(18);
output(2, 54) <= input(19);
output(2, 55) <= input(20);
output(2, 56) <= input(21);
output(2, 57) <= input(22);
output(2, 58) <= input(23);
output(2, 59) <= input(24);
output(2, 60) <= input(25);
output(2, 61) <= input(26);
output(2, 62) <= input(27);
output(2, 63) <= input(28);
output(2, 64) <= input(38);
output(2, 65) <= input(36);
output(2, 66) <= input(34);
output(2, 67) <= input(32);
output(2, 68) <= input(0);
output(2, 69) <= input(1);
output(2, 70) <= input(2);
output(2, 71) <= input(3);
output(2, 72) <= input(4);
output(2, 73) <= input(5);
output(2, 74) <= input(6);
output(2, 75) <= input(7);
output(2, 76) <= input(8);
output(2, 77) <= input(9);
output(2, 78) <= input(10);
output(2, 79) <= input(11);
output(2, 80) <= input(39);
output(2, 81) <= input(37);
output(2, 82) <= input(35);
output(2, 83) <= input(33);
output(2, 84) <= input(16);
output(2, 85) <= input(17);
output(2, 86) <= input(18);
output(2, 87) <= input(19);
output(2, 88) <= input(20);
output(2, 89) <= input(21);
output(2, 90) <= input(22);
output(2, 91) <= input(23);
output(2, 92) <= input(24);
output(2, 93) <= input(25);
output(2, 94) <= input(26);
output(2, 95) <= input(27);
output(2, 96) <= input(40);
output(2, 97) <= input(38);
output(2, 98) <= input(36);
output(2, 99) <= input(34);
output(2, 100) <= input(32);
output(2, 101) <= input(0);
output(2, 102) <= input(1);
output(2, 103) <= input(2);
output(2, 104) <= input(3);
output(2, 105) <= input(4);
output(2, 106) <= input(5);
output(2, 107) <= input(6);
output(2, 108) <= input(7);
output(2, 109) <= input(8);
output(2, 110) <= input(9);
output(2, 111) <= input(10);
output(2, 112) <= input(40);
output(2, 113) <= input(38);
output(2, 114) <= input(36);
output(2, 115) <= input(34);
output(2, 116) <= input(32);
output(2, 117) <= input(0);
output(2, 118) <= input(1);
output(2, 119) <= input(2);
output(2, 120) <= input(3);
output(2, 121) <= input(4);
output(2, 122) <= input(5);
output(2, 123) <= input(6);
output(2, 124) <= input(7);
output(2, 125) <= input(8);
output(2, 126) <= input(9);
output(2, 127) <= input(10);
output(2, 128) <= input(41);
output(2, 129) <= input(39);
output(2, 130) <= input(37);
output(2, 131) <= input(35);
output(2, 132) <= input(33);
output(2, 133) <= input(16);
output(2, 134) <= input(17);
output(2, 135) <= input(18);
output(2, 136) <= input(19);
output(2, 137) <= input(20);
output(2, 138) <= input(21);
output(2, 139) <= input(22);
output(2, 140) <= input(23);
output(2, 141) <= input(24);
output(2, 142) <= input(25);
output(2, 143) <= input(26);
output(2, 144) <= input(42);
output(2, 145) <= input(40);
output(2, 146) <= input(38);
output(2, 147) <= input(36);
output(2, 148) <= input(34);
output(2, 149) <= input(32);
output(2, 150) <= input(0);
output(2, 151) <= input(1);
output(2, 152) <= input(2);
output(2, 153) <= input(3);
output(2, 154) <= input(4);
output(2, 155) <= input(5);
output(2, 156) <= input(6);
output(2, 157) <= input(7);
output(2, 158) <= input(8);
output(2, 159) <= input(9);
output(2, 160) <= input(43);
output(2, 161) <= input(41);
output(2, 162) <= input(39);
output(2, 163) <= input(37);
output(2, 164) <= input(35);
output(2, 165) <= input(33);
output(2, 166) <= input(16);
output(2, 167) <= input(17);
output(2, 168) <= input(18);
output(2, 169) <= input(19);
output(2, 170) <= input(20);
output(2, 171) <= input(21);
output(2, 172) <= input(22);
output(2, 173) <= input(23);
output(2, 174) <= input(24);
output(2, 175) <= input(25);
output(2, 176) <= input(44);
output(2, 177) <= input(42);
output(2, 178) <= input(40);
output(2, 179) <= input(38);
output(2, 180) <= input(36);
output(2, 181) <= input(34);
output(2, 182) <= input(32);
output(2, 183) <= input(0);
output(2, 184) <= input(1);
output(2, 185) <= input(2);
output(2, 186) <= input(3);
output(2, 187) <= input(4);
output(2, 188) <= input(5);
output(2, 189) <= input(6);
output(2, 190) <= input(7);
output(2, 191) <= input(8);
output(2, 192) <= input(45);
output(2, 193) <= input(43);
output(2, 194) <= input(41);
output(2, 195) <= input(39);
output(2, 196) <= input(37);
output(2, 197) <= input(35);
output(2, 198) <= input(33);
output(2, 199) <= input(16);
output(2, 200) <= input(17);
output(2, 201) <= input(18);
output(2, 202) <= input(19);
output(2, 203) <= input(20);
output(2, 204) <= input(21);
output(2, 205) <= input(22);
output(2, 206) <= input(23);
output(2, 207) <= input(24);
output(2, 208) <= input(46);
output(2, 209) <= input(44);
output(2, 210) <= input(42);
output(2, 211) <= input(40);
output(2, 212) <= input(38);
output(2, 213) <= input(36);
output(2, 214) <= input(34);
output(2, 215) <= input(32);
output(2, 216) <= input(0);
output(2, 217) <= input(1);
output(2, 218) <= input(2);
output(2, 219) <= input(3);
output(2, 220) <= input(4);
output(2, 221) <= input(5);
output(2, 222) <= input(6);
output(2, 223) <= input(7);
output(2, 224) <= input(47);
output(2, 225) <= input(45);
output(2, 226) <= input(43);
output(2, 227) <= input(41);
output(2, 228) <= input(39);
output(2, 229) <= input(37);
output(2, 230) <= input(35);
output(2, 231) <= input(33);
output(2, 232) <= input(16);
output(2, 233) <= input(17);
output(2, 234) <= input(18);
output(2, 235) <= input(19);
output(2, 236) <= input(20);
output(2, 237) <= input(21);
output(2, 238) <= input(22);
output(2, 239) <= input(23);
output(2, 240) <= input(47);
output(2, 241) <= input(45);
output(2, 242) <= input(43);
output(2, 243) <= input(41);
output(2, 244) <= input(39);
output(2, 245) <= input(37);
output(2, 246) <= input(35);
output(2, 247) <= input(33);
output(2, 248) <= input(16);
output(2, 249) <= input(17);
output(2, 250) <= input(18);
output(2, 251) <= input(19);
output(2, 252) <= input(20);
output(2, 253) <= input(21);
output(2, 254) <= input(22);
output(2, 255) <= input(23);
when "0101" =>
output(0, 0) <= input(0);
output(0, 1) <= input(1);
output(0, 2) <= input(2);
output(0, 3) <= input(3);
output(0, 4) <= input(4);
output(0, 5) <= input(5);
output(0, 6) <= input(6);
output(0, 7) <= input(7);
output(0, 8) <= input(8);
output(0, 9) <= input(9);
output(0, 10) <= input(10);
output(0, 11) <= input(11);
output(0, 12) <= input(12);
output(0, 13) <= input(13);
output(0, 14) <= input(14);
output(0, 15) <= input(15);
output(0, 16) <= input(16);
output(0, 17) <= input(17);
output(0, 18) <= input(18);
output(0, 19) <= input(19);
output(0, 20) <= input(20);
output(0, 21) <= input(21);
output(0, 22) <= input(22);
output(0, 23) <= input(23);
output(0, 24) <= input(24);
output(0, 25) <= input(25);
output(0, 26) <= input(26);
output(0, 27) <= input(27);
output(0, 28) <= input(28);
output(0, 29) <= input(29);
output(0, 30) <= input(30);
output(0, 31) <= input(31);
output(0, 32) <= input(32);
output(0, 33) <= input(0);
output(0, 34) <= input(1);
output(0, 35) <= input(2);
output(0, 36) <= input(3);
output(0, 37) <= input(4);
output(0, 38) <= input(5);
output(0, 39) <= input(6);
output(0, 40) <= input(7);
output(0, 41) <= input(8);
output(0, 42) <= input(9);
output(0, 43) <= input(10);
output(0, 44) <= input(11);
output(0, 45) <= input(12);
output(0, 46) <= input(13);
output(0, 47) <= input(14);
output(0, 48) <= input(33);
output(0, 49) <= input(16);
output(0, 50) <= input(17);
output(0, 51) <= input(18);
output(0, 52) <= input(19);
output(0, 53) <= input(20);
output(0, 54) <= input(21);
output(0, 55) <= input(22);
output(0, 56) <= input(23);
output(0, 57) <= input(24);
output(0, 58) <= input(25);
output(0, 59) <= input(26);
output(0, 60) <= input(27);
output(0, 61) <= input(28);
output(0, 62) <= input(29);
output(0, 63) <= input(30);
output(0, 64) <= input(34);
output(0, 65) <= input(32);
output(0, 66) <= input(0);
output(0, 67) <= input(1);
output(0, 68) <= input(2);
output(0, 69) <= input(3);
output(0, 70) <= input(4);
output(0, 71) <= input(5);
output(0, 72) <= input(6);
output(0, 73) <= input(7);
output(0, 74) <= input(8);
output(0, 75) <= input(9);
output(0, 76) <= input(10);
output(0, 77) <= input(11);
output(0, 78) <= input(12);
output(0, 79) <= input(13);
output(0, 80) <= input(35);
output(0, 81) <= input(33);
output(0, 82) <= input(16);
output(0, 83) <= input(17);
output(0, 84) <= input(18);
output(0, 85) <= input(19);
output(0, 86) <= input(20);
output(0, 87) <= input(21);
output(0, 88) <= input(22);
output(0, 89) <= input(23);
output(0, 90) <= input(24);
output(0, 91) <= input(25);
output(0, 92) <= input(26);
output(0, 93) <= input(27);
output(0, 94) <= input(28);
output(0, 95) <= input(29);
output(0, 96) <= input(36);
output(0, 97) <= input(34);
output(0, 98) <= input(32);
output(0, 99) <= input(0);
output(0, 100) <= input(1);
output(0, 101) <= input(2);
output(0, 102) <= input(3);
output(0, 103) <= input(4);
output(0, 104) <= input(5);
output(0, 105) <= input(6);
output(0, 106) <= input(7);
output(0, 107) <= input(8);
output(0, 108) <= input(9);
output(0, 109) <= input(10);
output(0, 110) <= input(11);
output(0, 111) <= input(12);
output(0, 112) <= input(37);
output(0, 113) <= input(35);
output(0, 114) <= input(33);
output(0, 115) <= input(16);
output(0, 116) <= input(17);
output(0, 117) <= input(18);
output(0, 118) <= input(19);
output(0, 119) <= input(20);
output(0, 120) <= input(21);
output(0, 121) <= input(22);
output(0, 122) <= input(23);
output(0, 123) <= input(24);
output(0, 124) <= input(25);
output(0, 125) <= input(26);
output(0, 126) <= input(27);
output(0, 127) <= input(28);
output(0, 128) <= input(38);
output(0, 129) <= input(36);
output(0, 130) <= input(34);
output(0, 131) <= input(32);
output(0, 132) <= input(0);
output(0, 133) <= input(1);
output(0, 134) <= input(2);
output(0, 135) <= input(3);
output(0, 136) <= input(4);
output(0, 137) <= input(5);
output(0, 138) <= input(6);
output(0, 139) <= input(7);
output(0, 140) <= input(8);
output(0, 141) <= input(9);
output(0, 142) <= input(10);
output(0, 143) <= input(11);
output(0, 144) <= input(39);
output(0, 145) <= input(37);
output(0, 146) <= input(35);
output(0, 147) <= input(33);
output(0, 148) <= input(16);
output(0, 149) <= input(17);
output(0, 150) <= input(18);
output(0, 151) <= input(19);
output(0, 152) <= input(20);
output(0, 153) <= input(21);
output(0, 154) <= input(22);
output(0, 155) <= input(23);
output(0, 156) <= input(24);
output(0, 157) <= input(25);
output(0, 158) <= input(26);
output(0, 159) <= input(27);
output(0, 160) <= input(40);
output(0, 161) <= input(38);
output(0, 162) <= input(36);
output(0, 163) <= input(34);
output(0, 164) <= input(32);
output(0, 165) <= input(0);
output(0, 166) <= input(1);
output(0, 167) <= input(2);
output(0, 168) <= input(3);
output(0, 169) <= input(4);
output(0, 170) <= input(5);
output(0, 171) <= input(6);
output(0, 172) <= input(7);
output(0, 173) <= input(8);
output(0, 174) <= input(9);
output(0, 175) <= input(10);
output(0, 176) <= input(41);
output(0, 177) <= input(39);
output(0, 178) <= input(37);
output(0, 179) <= input(35);
output(0, 180) <= input(33);
output(0, 181) <= input(16);
output(0, 182) <= input(17);
output(0, 183) <= input(18);
output(0, 184) <= input(19);
output(0, 185) <= input(20);
output(0, 186) <= input(21);
output(0, 187) <= input(22);
output(0, 188) <= input(23);
output(0, 189) <= input(24);
output(0, 190) <= input(25);
output(0, 191) <= input(26);
output(0, 192) <= input(42);
output(0, 193) <= input(40);
output(0, 194) <= input(38);
output(0, 195) <= input(36);
output(0, 196) <= input(34);
output(0, 197) <= input(32);
output(0, 198) <= input(0);
output(0, 199) <= input(1);
output(0, 200) <= input(2);
output(0, 201) <= input(3);
output(0, 202) <= input(4);
output(0, 203) <= input(5);
output(0, 204) <= input(6);
output(0, 205) <= input(7);
output(0, 206) <= input(8);
output(0, 207) <= input(9);
output(0, 208) <= input(43);
output(0, 209) <= input(41);
output(0, 210) <= input(39);
output(0, 211) <= input(37);
output(0, 212) <= input(35);
output(0, 213) <= input(33);
output(0, 214) <= input(16);
output(0, 215) <= input(17);
output(0, 216) <= input(18);
output(0, 217) <= input(19);
output(0, 218) <= input(20);
output(0, 219) <= input(21);
output(0, 220) <= input(22);
output(0, 221) <= input(23);
output(0, 222) <= input(24);
output(0, 223) <= input(25);
output(0, 224) <= input(44);
output(0, 225) <= input(42);
output(0, 226) <= input(40);
output(0, 227) <= input(38);
output(0, 228) <= input(36);
output(0, 229) <= input(34);
output(0, 230) <= input(32);
output(0, 231) <= input(0);
output(0, 232) <= input(1);
output(0, 233) <= input(2);
output(0, 234) <= input(3);
output(0, 235) <= input(4);
output(0, 236) <= input(5);
output(0, 237) <= input(6);
output(0, 238) <= input(7);
output(0, 239) <= input(8);
output(0, 240) <= input(45);
output(0, 241) <= input(43);
output(0, 242) <= input(41);
output(0, 243) <= input(39);
output(0, 244) <= input(37);
output(0, 245) <= input(35);
output(0, 246) <= input(33);
output(0, 247) <= input(16);
output(0, 248) <= input(17);
output(0, 249) <= input(18);
output(0, 250) <= input(19);
output(0, 251) <= input(20);
output(0, 252) <= input(21);
output(0, 253) <= input(22);
output(0, 254) <= input(23);
output(0, 255) <= input(24);
output(1, 0) <= input(33);
output(1, 1) <= input(16);
output(1, 2) <= input(17);
output(1, 3) <= input(18);
output(1, 4) <= input(19);
output(1, 5) <= input(20);
output(1, 6) <= input(21);
output(1, 7) <= input(22);
output(1, 8) <= input(23);
output(1, 9) <= input(24);
output(1, 10) <= input(25);
output(1, 11) <= input(26);
output(1, 12) <= input(27);
output(1, 13) <= input(28);
output(1, 14) <= input(29);
output(1, 15) <= input(30);
output(1, 16) <= input(34);
output(1, 17) <= input(32);
output(1, 18) <= input(0);
output(1, 19) <= input(1);
output(1, 20) <= input(2);
output(1, 21) <= input(3);
output(1, 22) <= input(4);
output(1, 23) <= input(5);
output(1, 24) <= input(6);
output(1, 25) <= input(7);
output(1, 26) <= input(8);
output(1, 27) <= input(9);
output(1, 28) <= input(10);
output(1, 29) <= input(11);
output(1, 30) <= input(12);
output(1, 31) <= input(13);
output(1, 32) <= input(35);
output(1, 33) <= input(33);
output(1, 34) <= input(16);
output(1, 35) <= input(17);
output(1, 36) <= input(18);
output(1, 37) <= input(19);
output(1, 38) <= input(20);
output(1, 39) <= input(21);
output(1, 40) <= input(22);
output(1, 41) <= input(23);
output(1, 42) <= input(24);
output(1, 43) <= input(25);
output(1, 44) <= input(26);
output(1, 45) <= input(27);
output(1, 46) <= input(28);
output(1, 47) <= input(29);
output(1, 48) <= input(36);
output(1, 49) <= input(34);
output(1, 50) <= input(32);
output(1, 51) <= input(0);
output(1, 52) <= input(1);
output(1, 53) <= input(2);
output(1, 54) <= input(3);
output(1, 55) <= input(4);
output(1, 56) <= input(5);
output(1, 57) <= input(6);
output(1, 58) <= input(7);
output(1, 59) <= input(8);
output(1, 60) <= input(9);
output(1, 61) <= input(10);
output(1, 62) <= input(11);
output(1, 63) <= input(12);
output(1, 64) <= input(37);
output(1, 65) <= input(35);
output(1, 66) <= input(33);
output(1, 67) <= input(16);
output(1, 68) <= input(17);
output(1, 69) <= input(18);
output(1, 70) <= input(19);
output(1, 71) <= input(20);
output(1, 72) <= input(21);
output(1, 73) <= input(22);
output(1, 74) <= input(23);
output(1, 75) <= input(24);
output(1, 76) <= input(25);
output(1, 77) <= input(26);
output(1, 78) <= input(27);
output(1, 79) <= input(28);
output(1, 80) <= input(38);
output(1, 81) <= input(36);
output(1, 82) <= input(34);
output(1, 83) <= input(32);
output(1, 84) <= input(0);
output(1, 85) <= input(1);
output(1, 86) <= input(2);
output(1, 87) <= input(3);
output(1, 88) <= input(4);
output(1, 89) <= input(5);
output(1, 90) <= input(6);
output(1, 91) <= input(7);
output(1, 92) <= input(8);
output(1, 93) <= input(9);
output(1, 94) <= input(10);
output(1, 95) <= input(11);
output(1, 96) <= input(39);
output(1, 97) <= input(37);
output(1, 98) <= input(35);
output(1, 99) <= input(33);
output(1, 100) <= input(16);
output(1, 101) <= input(17);
output(1, 102) <= input(18);
output(1, 103) <= input(19);
output(1, 104) <= input(20);
output(1, 105) <= input(21);
output(1, 106) <= input(22);
output(1, 107) <= input(23);
output(1, 108) <= input(24);
output(1, 109) <= input(25);
output(1, 110) <= input(26);
output(1, 111) <= input(27);
output(1, 112) <= input(40);
output(1, 113) <= input(38);
output(1, 114) <= input(36);
output(1, 115) <= input(34);
output(1, 116) <= input(32);
output(1, 117) <= input(0);
output(1, 118) <= input(1);
output(1, 119) <= input(2);
output(1, 120) <= input(3);
output(1, 121) <= input(4);
output(1, 122) <= input(5);
output(1, 123) <= input(6);
output(1, 124) <= input(7);
output(1, 125) <= input(8);
output(1, 126) <= input(9);
output(1, 127) <= input(10);
output(1, 128) <= input(42);
output(1, 129) <= input(40);
output(1, 130) <= input(38);
output(1, 131) <= input(36);
output(1, 132) <= input(34);
output(1, 133) <= input(32);
output(1, 134) <= input(0);
output(1, 135) <= input(1);
output(1, 136) <= input(2);
output(1, 137) <= input(3);
output(1, 138) <= input(4);
output(1, 139) <= input(5);
output(1, 140) <= input(6);
output(1, 141) <= input(7);
output(1, 142) <= input(8);
output(1, 143) <= input(9);
output(1, 144) <= input(43);
output(1, 145) <= input(41);
output(1, 146) <= input(39);
output(1, 147) <= input(37);
output(1, 148) <= input(35);
output(1, 149) <= input(33);
output(1, 150) <= input(16);
output(1, 151) <= input(17);
output(1, 152) <= input(18);
output(1, 153) <= input(19);
output(1, 154) <= input(20);
output(1, 155) <= input(21);
output(1, 156) <= input(22);
output(1, 157) <= input(23);
output(1, 158) <= input(24);
output(1, 159) <= input(25);
output(1, 160) <= input(44);
output(1, 161) <= input(42);
output(1, 162) <= input(40);
output(1, 163) <= input(38);
output(1, 164) <= input(36);
output(1, 165) <= input(34);
output(1, 166) <= input(32);
output(1, 167) <= input(0);
output(1, 168) <= input(1);
output(1, 169) <= input(2);
output(1, 170) <= input(3);
output(1, 171) <= input(4);
output(1, 172) <= input(5);
output(1, 173) <= input(6);
output(1, 174) <= input(7);
output(1, 175) <= input(8);
output(1, 176) <= input(45);
output(1, 177) <= input(43);
output(1, 178) <= input(41);
output(1, 179) <= input(39);
output(1, 180) <= input(37);
output(1, 181) <= input(35);
output(1, 182) <= input(33);
output(1, 183) <= input(16);
output(1, 184) <= input(17);
output(1, 185) <= input(18);
output(1, 186) <= input(19);
output(1, 187) <= input(20);
output(1, 188) <= input(21);
output(1, 189) <= input(22);
output(1, 190) <= input(23);
output(1, 191) <= input(24);
output(1, 192) <= input(46);
output(1, 193) <= input(44);
output(1, 194) <= input(42);
output(1, 195) <= input(40);
output(1, 196) <= input(38);
output(1, 197) <= input(36);
output(1, 198) <= input(34);
output(1, 199) <= input(32);
output(1, 200) <= input(0);
output(1, 201) <= input(1);
output(1, 202) <= input(2);
output(1, 203) <= input(3);
output(1, 204) <= input(4);
output(1, 205) <= input(5);
output(1, 206) <= input(6);
output(1, 207) <= input(7);
output(1, 208) <= input(47);
output(1, 209) <= input(45);
output(1, 210) <= input(43);
output(1, 211) <= input(41);
output(1, 212) <= input(39);
output(1, 213) <= input(37);
output(1, 214) <= input(35);
output(1, 215) <= input(33);
output(1, 216) <= input(16);
output(1, 217) <= input(17);
output(1, 218) <= input(18);
output(1, 219) <= input(19);
output(1, 220) <= input(20);
output(1, 221) <= input(21);
output(1, 222) <= input(22);
output(1, 223) <= input(23);
output(1, 224) <= input(48);
output(1, 225) <= input(46);
output(1, 226) <= input(44);
output(1, 227) <= input(42);
output(1, 228) <= input(40);
output(1, 229) <= input(38);
output(1, 230) <= input(36);
output(1, 231) <= input(34);
output(1, 232) <= input(32);
output(1, 233) <= input(0);
output(1, 234) <= input(1);
output(1, 235) <= input(2);
output(1, 236) <= input(3);
output(1, 237) <= input(4);
output(1, 238) <= input(5);
output(1, 239) <= input(6);
output(1, 240) <= input(49);
output(1, 241) <= input(47);
output(1, 242) <= input(45);
output(1, 243) <= input(43);
output(1, 244) <= input(41);
output(1, 245) <= input(39);
output(1, 246) <= input(37);
output(1, 247) <= input(35);
output(1, 248) <= input(33);
output(1, 249) <= input(16);
output(1, 250) <= input(17);
output(1, 251) <= input(18);
output(1, 252) <= input(19);
output(1, 253) <= input(20);
output(1, 254) <= input(21);
output(1, 255) <= input(22);
when "0110" =>
output(0, 0) <= input(0);
output(0, 1) <= input(1);
output(0, 2) <= input(2);
output(0, 3) <= input(3);
output(0, 4) <= input(4);
output(0, 5) <= input(5);
output(0, 6) <= input(6);
output(0, 7) <= input(7);
output(0, 8) <= input(8);
output(0, 9) <= input(9);
output(0, 10) <= input(10);
output(0, 11) <= input(11);
output(0, 12) <= input(12);
output(0, 13) <= input(13);
output(0, 14) <= input(14);
output(0, 15) <= input(15);
output(0, 16) <= input(16);
output(0, 17) <= input(17);
output(0, 18) <= input(18);
output(0, 19) <= input(19);
output(0, 20) <= input(20);
output(0, 21) <= input(21);
output(0, 22) <= input(22);
output(0, 23) <= input(23);
output(0, 24) <= input(24);
output(0, 25) <= input(25);
output(0, 26) <= input(26);
output(0, 27) <= input(27);
output(0, 28) <= input(28);
output(0, 29) <= input(29);
output(0, 30) <= input(30);
output(0, 31) <= input(31);
output(0, 32) <= input(32);
output(0, 33) <= input(0);
output(0, 34) <= input(1);
output(0, 35) <= input(2);
output(0, 36) <= input(3);
output(0, 37) <= input(4);
output(0, 38) <= input(5);
output(0, 39) <= input(6);
output(0, 40) <= input(7);
output(0, 41) <= input(8);
output(0, 42) <= input(9);
output(0, 43) <= input(10);
output(0, 44) <= input(11);
output(0, 45) <= input(12);
output(0, 46) <= input(13);
output(0, 47) <= input(14);
output(0, 48) <= input(33);
output(0, 49) <= input(16);
output(0, 50) <= input(17);
output(0, 51) <= input(18);
output(0, 52) <= input(19);
output(0, 53) <= input(20);
output(0, 54) <= input(21);
output(0, 55) <= input(22);
output(0, 56) <= input(23);
output(0, 57) <= input(24);
output(0, 58) <= input(25);
output(0, 59) <= input(26);
output(0, 60) <= input(27);
output(0, 61) <= input(28);
output(0, 62) <= input(29);
output(0, 63) <= input(30);
output(0, 64) <= input(34);
output(0, 65) <= input(33);
output(0, 66) <= input(16);
output(0, 67) <= input(17);
output(0, 68) <= input(18);
output(0, 69) <= input(19);
output(0, 70) <= input(20);
output(0, 71) <= input(21);
output(0, 72) <= input(22);
output(0, 73) <= input(23);
output(0, 74) <= input(24);
output(0, 75) <= input(25);
output(0, 76) <= input(26);
output(0, 77) <= input(27);
output(0, 78) <= input(28);
output(0, 79) <= input(29);
output(0, 80) <= input(35);
output(0, 81) <= input(36);
output(0, 82) <= input(32);
output(0, 83) <= input(0);
output(0, 84) <= input(1);
output(0, 85) <= input(2);
output(0, 86) <= input(3);
output(0, 87) <= input(4);
output(0, 88) <= input(5);
output(0, 89) <= input(6);
output(0, 90) <= input(7);
output(0, 91) <= input(8);
output(0, 92) <= input(9);
output(0, 93) <= input(10);
output(0, 94) <= input(11);
output(0, 95) <= input(12);
output(0, 96) <= input(37);
output(0, 97) <= input(34);
output(0, 98) <= input(33);
output(0, 99) <= input(16);
output(0, 100) <= input(17);
output(0, 101) <= input(18);
output(0, 102) <= input(19);
output(0, 103) <= input(20);
output(0, 104) <= input(21);
output(0, 105) <= input(22);
output(0, 106) <= input(23);
output(0, 107) <= input(24);
output(0, 108) <= input(25);
output(0, 109) <= input(26);
output(0, 110) <= input(27);
output(0, 111) <= input(28);
output(0, 112) <= input(38);
output(0, 113) <= input(35);
output(0, 114) <= input(36);
output(0, 115) <= input(32);
output(0, 116) <= input(0);
output(0, 117) <= input(1);
output(0, 118) <= input(2);
output(0, 119) <= input(3);
output(0, 120) <= input(4);
output(0, 121) <= input(5);
output(0, 122) <= input(6);
output(0, 123) <= input(7);
output(0, 124) <= input(8);
output(0, 125) <= input(9);
output(0, 126) <= input(10);
output(0, 127) <= input(11);
output(0, 128) <= input(39);
output(0, 129) <= input(38);
output(0, 130) <= input(35);
output(0, 131) <= input(36);
output(0, 132) <= input(32);
output(0, 133) <= input(0);
output(0, 134) <= input(1);
output(0, 135) <= input(2);
output(0, 136) <= input(3);
output(0, 137) <= input(4);
output(0, 138) <= input(5);
output(0, 139) <= input(6);
output(0, 140) <= input(7);
output(0, 141) <= input(8);
output(0, 142) <= input(9);
output(0, 143) <= input(10);
output(0, 144) <= input(40);
output(0, 145) <= input(41);
output(0, 146) <= input(37);
output(0, 147) <= input(34);
output(0, 148) <= input(33);
output(0, 149) <= input(16);
output(0, 150) <= input(17);
output(0, 151) <= input(18);
output(0, 152) <= input(19);
output(0, 153) <= input(20);
output(0, 154) <= input(21);
output(0, 155) <= input(22);
output(0, 156) <= input(23);
output(0, 157) <= input(24);
output(0, 158) <= input(25);
output(0, 159) <= input(26);
output(0, 160) <= input(42);
output(0, 161) <= input(39);
output(0, 162) <= input(38);
output(0, 163) <= input(35);
output(0, 164) <= input(36);
output(0, 165) <= input(32);
output(0, 166) <= input(0);
output(0, 167) <= input(1);
output(0, 168) <= input(2);
output(0, 169) <= input(3);
output(0, 170) <= input(4);
output(0, 171) <= input(5);
output(0, 172) <= input(6);
output(0, 173) <= input(7);
output(0, 174) <= input(8);
output(0, 175) <= input(9);
output(0, 176) <= input(43);
output(0, 177) <= input(40);
output(0, 178) <= input(41);
output(0, 179) <= input(37);
output(0, 180) <= input(34);
output(0, 181) <= input(33);
output(0, 182) <= input(16);
output(0, 183) <= input(17);
output(0, 184) <= input(18);
output(0, 185) <= input(19);
output(0, 186) <= input(20);
output(0, 187) <= input(21);
output(0, 188) <= input(22);
output(0, 189) <= input(23);
output(0, 190) <= input(24);
output(0, 191) <= input(25);
output(0, 192) <= input(44);
output(0, 193) <= input(43);
output(0, 194) <= input(40);
output(0, 195) <= input(41);
output(0, 196) <= input(37);
output(0, 197) <= input(34);
output(0, 198) <= input(33);
output(0, 199) <= input(16);
output(0, 200) <= input(17);
output(0, 201) <= input(18);
output(0, 202) <= input(19);
output(0, 203) <= input(20);
output(0, 204) <= input(21);
output(0, 205) <= input(22);
output(0, 206) <= input(23);
output(0, 207) <= input(24);
output(0, 208) <= input(45);
output(0, 209) <= input(46);
output(0, 210) <= input(42);
output(0, 211) <= input(39);
output(0, 212) <= input(38);
output(0, 213) <= input(35);
output(0, 214) <= input(36);
output(0, 215) <= input(32);
output(0, 216) <= input(0);
output(0, 217) <= input(1);
output(0, 218) <= input(2);
output(0, 219) <= input(3);
output(0, 220) <= input(4);
output(0, 221) <= input(5);
output(0, 222) <= input(6);
output(0, 223) <= input(7);
output(0, 224) <= input(47);
output(0, 225) <= input(44);
output(0, 226) <= input(43);
output(0, 227) <= input(40);
output(0, 228) <= input(41);
output(0, 229) <= input(37);
output(0, 230) <= input(34);
output(0, 231) <= input(33);
output(0, 232) <= input(16);
output(0, 233) <= input(17);
output(0, 234) <= input(18);
output(0, 235) <= input(19);
output(0, 236) <= input(20);
output(0, 237) <= input(21);
output(0, 238) <= input(22);
output(0, 239) <= input(23);
output(0, 240) <= input(48);
output(0, 241) <= input(45);
output(0, 242) <= input(46);
output(0, 243) <= input(42);
output(0, 244) <= input(39);
output(0, 245) <= input(38);
output(0, 246) <= input(35);
output(0, 247) <= input(36);
output(0, 248) <= input(32);
output(0, 249) <= input(0);
output(0, 250) <= input(1);
output(0, 251) <= input(2);
output(0, 252) <= input(3);
output(0, 253) <= input(4);
output(0, 254) <= input(5);
output(0, 255) <= input(6);
output(1, 0) <= input(33);
output(1, 1) <= input(16);
output(1, 2) <= input(17);
output(1, 3) <= input(18);
output(1, 4) <= input(19);
output(1, 5) <= input(20);
output(1, 6) <= input(21);
output(1, 7) <= input(22);
output(1, 8) <= input(23);
output(1, 9) <= input(24);
output(1, 10) <= input(25);
output(1, 11) <= input(26);
output(1, 12) <= input(27);
output(1, 13) <= input(28);
output(1, 14) <= input(29);
output(1, 15) <= input(30);
output(1, 16) <= input(36);
output(1, 17) <= input(32);
output(1, 18) <= input(0);
output(1, 19) <= input(1);
output(1, 20) <= input(2);
output(1, 21) <= input(3);
output(1, 22) <= input(4);
output(1, 23) <= input(5);
output(1, 24) <= input(6);
output(1, 25) <= input(7);
output(1, 26) <= input(8);
output(1, 27) <= input(9);
output(1, 28) <= input(10);
output(1, 29) <= input(11);
output(1, 30) <= input(12);
output(1, 31) <= input(13);
output(1, 32) <= input(35);
output(1, 33) <= input(36);
output(1, 34) <= input(32);
output(1, 35) <= input(0);
output(1, 36) <= input(1);
output(1, 37) <= input(2);
output(1, 38) <= input(3);
output(1, 39) <= input(4);
output(1, 40) <= input(5);
output(1, 41) <= input(6);
output(1, 42) <= input(7);
output(1, 43) <= input(8);
output(1, 44) <= input(9);
output(1, 45) <= input(10);
output(1, 46) <= input(11);
output(1, 47) <= input(12);
output(1, 48) <= input(37);
output(1, 49) <= input(34);
output(1, 50) <= input(33);
output(1, 51) <= input(16);
output(1, 52) <= input(17);
output(1, 53) <= input(18);
output(1, 54) <= input(19);
output(1, 55) <= input(20);
output(1, 56) <= input(21);
output(1, 57) <= input(22);
output(1, 58) <= input(23);
output(1, 59) <= input(24);
output(1, 60) <= input(25);
output(1, 61) <= input(26);
output(1, 62) <= input(27);
output(1, 63) <= input(28);
output(1, 64) <= input(41);
output(1, 65) <= input(37);
output(1, 66) <= input(34);
output(1, 67) <= input(33);
output(1, 68) <= input(16);
output(1, 69) <= input(17);
output(1, 70) <= input(18);
output(1, 71) <= input(19);
output(1, 72) <= input(20);
output(1, 73) <= input(21);
output(1, 74) <= input(22);
output(1, 75) <= input(23);
output(1, 76) <= input(24);
output(1, 77) <= input(25);
output(1, 78) <= input(26);
output(1, 79) <= input(27);
output(1, 80) <= input(39);
output(1, 81) <= input(38);
output(1, 82) <= input(35);
output(1, 83) <= input(36);
output(1, 84) <= input(32);
output(1, 85) <= input(0);
output(1, 86) <= input(1);
output(1, 87) <= input(2);
output(1, 88) <= input(3);
output(1, 89) <= input(4);
output(1, 90) <= input(5);
output(1, 91) <= input(6);
output(1, 92) <= input(7);
output(1, 93) <= input(8);
output(1, 94) <= input(9);
output(1, 95) <= input(10);
output(1, 96) <= input(49);
output(1, 97) <= input(39);
output(1, 98) <= input(38);
output(1, 99) <= input(35);
output(1, 100) <= input(36);
output(1, 101) <= input(32);
output(1, 102) <= input(0);
output(1, 103) <= input(1);
output(1, 104) <= input(2);
output(1, 105) <= input(3);
output(1, 106) <= input(4);
output(1, 107) <= input(5);
output(1, 108) <= input(6);
output(1, 109) <= input(7);
output(1, 110) <= input(8);
output(1, 111) <= input(9);
output(1, 112) <= input(50);
output(1, 113) <= input(51);
output(1, 114) <= input(41);
output(1, 115) <= input(37);
output(1, 116) <= input(34);
output(1, 117) <= input(33);
output(1, 118) <= input(16);
output(1, 119) <= input(17);
output(1, 120) <= input(18);
output(1, 121) <= input(19);
output(1, 122) <= input(20);
output(1, 123) <= input(21);
output(1, 124) <= input(22);
output(1, 125) <= input(23);
output(1, 126) <= input(24);
output(1, 127) <= input(25);
output(1, 128) <= input(52);
output(1, 129) <= input(49);
output(1, 130) <= input(39);
output(1, 131) <= input(38);
output(1, 132) <= input(35);
output(1, 133) <= input(36);
output(1, 134) <= input(32);
output(1, 135) <= input(0);
output(1, 136) <= input(1);
output(1, 137) <= input(2);
output(1, 138) <= input(3);
output(1, 139) <= input(4);
output(1, 140) <= input(5);
output(1, 141) <= input(6);
output(1, 142) <= input(7);
output(1, 143) <= input(8);
output(1, 144) <= input(53);
output(1, 145) <= input(52);
output(1, 146) <= input(49);
output(1, 147) <= input(39);
output(1, 148) <= input(38);
output(1, 149) <= input(35);
output(1, 150) <= input(36);
output(1, 151) <= input(32);
output(1, 152) <= input(0);
output(1, 153) <= input(1);
output(1, 154) <= input(2);
output(1, 155) <= input(3);
output(1, 156) <= input(4);
output(1, 157) <= input(5);
output(1, 158) <= input(6);
output(1, 159) <= input(7);
output(1, 160) <= input(54);
output(1, 161) <= input(55);
output(1, 162) <= input(50);
output(1, 163) <= input(51);
output(1, 164) <= input(41);
output(1, 165) <= input(37);
output(1, 166) <= input(34);
output(1, 167) <= input(33);
output(1, 168) <= input(16);
output(1, 169) <= input(17);
output(1, 170) <= input(18);
output(1, 171) <= input(19);
output(1, 172) <= input(20);
output(1, 173) <= input(21);
output(1, 174) <= input(22);
output(1, 175) <= input(23);
output(1, 176) <= input(56);
output(1, 177) <= input(54);
output(1, 178) <= input(55);
output(1, 179) <= input(50);
output(1, 180) <= input(51);
output(1, 181) <= input(41);
output(1, 182) <= input(37);
output(1, 183) <= input(34);
output(1, 184) <= input(33);
output(1, 185) <= input(16);
output(1, 186) <= input(17);
output(1, 187) <= input(18);
output(1, 188) <= input(19);
output(1, 189) <= input(20);
output(1, 190) <= input(21);
output(1, 191) <= input(22);
output(1, 192) <= input(57);
output(1, 193) <= input(58);
output(1, 194) <= input(53);
output(1, 195) <= input(52);
output(1, 196) <= input(49);
output(1, 197) <= input(39);
output(1, 198) <= input(38);
output(1, 199) <= input(35);
output(1, 200) <= input(36);
output(1, 201) <= input(32);
output(1, 202) <= input(0);
output(1, 203) <= input(1);
output(1, 204) <= input(2);
output(1, 205) <= input(3);
output(1, 206) <= input(4);
output(1, 207) <= input(5);
output(1, 208) <= input(59);
output(1, 209) <= input(57);
output(1, 210) <= input(58);
output(1, 211) <= input(53);
output(1, 212) <= input(52);
output(1, 213) <= input(49);
output(1, 214) <= input(39);
output(1, 215) <= input(38);
output(1, 216) <= input(35);
output(1, 217) <= input(36);
output(1, 218) <= input(32);
output(1, 219) <= input(0);
output(1, 220) <= input(1);
output(1, 221) <= input(2);
output(1, 222) <= input(3);
output(1, 223) <= input(4);
output(1, 224) <= input(60);
output(1, 225) <= input(61);
output(1, 226) <= input(56);
output(1, 227) <= input(54);
output(1, 228) <= input(55);
output(1, 229) <= input(50);
output(1, 230) <= input(51);
output(1, 231) <= input(41);
output(1, 232) <= input(37);
output(1, 233) <= input(34);
output(1, 234) <= input(33);
output(1, 235) <= input(16);
output(1, 236) <= input(17);
output(1, 237) <= input(18);
output(1, 238) <= input(19);
output(1, 239) <= input(20);
output(1, 240) <= input(62);
output(1, 241) <= input(59);
output(1, 242) <= input(57);
output(1, 243) <= input(58);
output(1, 244) <= input(53);
output(1, 245) <= input(52);
output(1, 246) <= input(49);
output(1, 247) <= input(39);
output(1, 248) <= input(38);
output(1, 249) <= input(35);
output(1, 250) <= input(36);
output(1, 251) <= input(32);
output(1, 252) <= input(0);
output(1, 253) <= input(1);
output(1, 254) <= input(2);
output(1, 255) <= input(3);
output(2, 0) <= input(35);
output(2, 1) <= input(36);
output(2, 2) <= input(32);
output(2, 3) <= input(0);
output(2, 4) <= input(1);
output(2, 5) <= input(2);
output(2, 6) <= input(3);
output(2, 7) <= input(4);
output(2, 8) <= input(5);
output(2, 9) <= input(6);
output(2, 10) <= input(7);
output(2, 11) <= input(8);
output(2, 12) <= input(9);
output(2, 13) <= input(10);
output(2, 14) <= input(11);
output(2, 15) <= input(12);
output(2, 16) <= input(38);
output(2, 17) <= input(35);
output(2, 18) <= input(36);
output(2, 19) <= input(32);
output(2, 20) <= input(0);
output(2, 21) <= input(1);
output(2, 22) <= input(2);
output(2, 23) <= input(3);
output(2, 24) <= input(4);
output(2, 25) <= input(5);
output(2, 26) <= input(6);
output(2, 27) <= input(7);
output(2, 28) <= input(8);
output(2, 29) <= input(9);
output(2, 30) <= input(10);
output(2, 31) <= input(11);
output(2, 32) <= input(41);
output(2, 33) <= input(37);
output(2, 34) <= input(34);
output(2, 35) <= input(33);
output(2, 36) <= input(16);
output(2, 37) <= input(17);
output(2, 38) <= input(18);
output(2, 39) <= input(19);
output(2, 40) <= input(20);
output(2, 41) <= input(21);
output(2, 42) <= input(22);
output(2, 43) <= input(23);
output(2, 44) <= input(24);
output(2, 45) <= input(25);
output(2, 46) <= input(26);
output(2, 47) <= input(27);
output(2, 48) <= input(51);
output(2, 49) <= input(41);
output(2, 50) <= input(37);
output(2, 51) <= input(34);
output(2, 52) <= input(33);
output(2, 53) <= input(16);
output(2, 54) <= input(17);
output(2, 55) <= input(18);
output(2, 56) <= input(19);
output(2, 57) <= input(20);
output(2, 58) <= input(21);
output(2, 59) <= input(22);
output(2, 60) <= input(23);
output(2, 61) <= input(24);
output(2, 62) <= input(25);
output(2, 63) <= input(26);
output(2, 64) <= input(63);
output(2, 65) <= input(51);
output(2, 66) <= input(41);
output(2, 67) <= input(37);
output(2, 68) <= input(34);
output(2, 69) <= input(33);
output(2, 70) <= input(16);
output(2, 71) <= input(17);
output(2, 72) <= input(18);
output(2, 73) <= input(19);
output(2, 74) <= input(20);
output(2, 75) <= input(21);
output(2, 76) <= input(22);
output(2, 77) <= input(23);
output(2, 78) <= input(24);
output(2, 79) <= input(25);
output(2, 80) <= input(64);
output(2, 81) <= input(49);
output(2, 82) <= input(39);
output(2, 83) <= input(38);
output(2, 84) <= input(35);
output(2, 85) <= input(36);
output(2, 86) <= input(32);
output(2, 87) <= input(0);
output(2, 88) <= input(1);
output(2, 89) <= input(2);
output(2, 90) <= input(3);
output(2, 91) <= input(4);
output(2, 92) <= input(5);
output(2, 93) <= input(6);
output(2, 94) <= input(7);
output(2, 95) <= input(8);
output(2, 96) <= input(65);
output(2, 97) <= input(64);
output(2, 98) <= input(49);
output(2, 99) <= input(39);
output(2, 100) <= input(38);
output(2, 101) <= input(35);
output(2, 102) <= input(36);
output(2, 103) <= input(32);
output(2, 104) <= input(0);
output(2, 105) <= input(1);
output(2, 106) <= input(2);
output(2, 107) <= input(3);
output(2, 108) <= input(4);
output(2, 109) <= input(5);
output(2, 110) <= input(6);
output(2, 111) <= input(7);
output(2, 112) <= input(66);
output(2, 113) <= input(67);
output(2, 114) <= input(63);
output(2, 115) <= input(51);
output(2, 116) <= input(41);
output(2, 117) <= input(37);
output(2, 118) <= input(34);
output(2, 119) <= input(33);
output(2, 120) <= input(16);
output(2, 121) <= input(17);
output(2, 122) <= input(18);
output(2, 123) <= input(19);
output(2, 124) <= input(20);
output(2, 125) <= input(21);
output(2, 126) <= input(22);
output(2, 127) <= input(23);
output(2, 128) <= input(68);
output(2, 129) <= input(66);
output(2, 130) <= input(67);
output(2, 131) <= input(63);
output(2, 132) <= input(51);
output(2, 133) <= input(41);
output(2, 134) <= input(37);
output(2, 135) <= input(34);
output(2, 136) <= input(33);
output(2, 137) <= input(16);
output(2, 138) <= input(17);
output(2, 139) <= input(18);
output(2, 140) <= input(19);
output(2, 141) <= input(20);
output(2, 142) <= input(21);
output(2, 143) <= input(22);
output(2, 144) <= input(69);
output(2, 145) <= input(68);
output(2, 146) <= input(66);
output(2, 147) <= input(67);
output(2, 148) <= input(63);
output(2, 149) <= input(51);
output(2, 150) <= input(41);
output(2, 151) <= input(37);
output(2, 152) <= input(34);
output(2, 153) <= input(33);
output(2, 154) <= input(16);
output(2, 155) <= input(17);
output(2, 156) <= input(18);
output(2, 157) <= input(19);
output(2, 158) <= input(20);
output(2, 159) <= input(21);
output(2, 160) <= input(70);
output(2, 161) <= input(71);
output(2, 162) <= input(72);
output(2, 163) <= input(65);
output(2, 164) <= input(64);
output(2, 165) <= input(49);
output(2, 166) <= input(39);
output(2, 167) <= input(38);
output(2, 168) <= input(35);
output(2, 169) <= input(36);
output(2, 170) <= input(32);
output(2, 171) <= input(0);
output(2, 172) <= input(1);
output(2, 173) <= input(2);
output(2, 174) <= input(3);
output(2, 175) <= input(4);
output(2, 176) <= input(73);
output(2, 177) <= input(70);
output(2, 178) <= input(71);
output(2, 179) <= input(72);
output(2, 180) <= input(65);
output(2, 181) <= input(64);
output(2, 182) <= input(49);
output(2, 183) <= input(39);
output(2, 184) <= input(38);
output(2, 185) <= input(35);
output(2, 186) <= input(36);
output(2, 187) <= input(32);
output(2, 188) <= input(0);
output(2, 189) <= input(1);
output(2, 190) <= input(2);
output(2, 191) <= input(3);
output(2, 192) <= input(74);
output(2, 193) <= input(73);
output(2, 194) <= input(70);
output(2, 195) <= input(71);
output(2, 196) <= input(72);
output(2, 197) <= input(65);
output(2, 198) <= input(64);
output(2, 199) <= input(49);
output(2, 200) <= input(39);
output(2, 201) <= input(38);
output(2, 202) <= input(35);
output(2, 203) <= input(36);
output(2, 204) <= input(32);
output(2, 205) <= input(0);
output(2, 206) <= input(1);
output(2, 207) <= input(2);
output(2, 208) <= input(75);
output(2, 209) <= input(76);
output(2, 210) <= input(77);
output(2, 211) <= input(69);
output(2, 212) <= input(68);
output(2, 213) <= input(66);
output(2, 214) <= input(67);
output(2, 215) <= input(63);
output(2, 216) <= input(51);
output(2, 217) <= input(41);
output(2, 218) <= input(37);
output(2, 219) <= input(34);
output(2, 220) <= input(33);
output(2, 221) <= input(16);
output(2, 222) <= input(17);
output(2, 223) <= input(18);
output(2, 224) <= input(78);
output(2, 225) <= input(75);
output(2, 226) <= input(76);
output(2, 227) <= input(77);
output(2, 228) <= input(69);
output(2, 229) <= input(68);
output(2, 230) <= input(66);
output(2, 231) <= input(67);
output(2, 232) <= input(63);
output(2, 233) <= input(51);
output(2, 234) <= input(41);
output(2, 235) <= input(37);
output(2, 236) <= input(34);
output(2, 237) <= input(33);
output(2, 238) <= input(16);
output(2, 239) <= input(17);
output(2, 240) <= input(79);
output(2, 241) <= input(80);
output(2, 242) <= input(74);
output(2, 243) <= input(73);
output(2, 244) <= input(70);
output(2, 245) <= input(71);
output(2, 246) <= input(72);
output(2, 247) <= input(65);
output(2, 248) <= input(64);
output(2, 249) <= input(49);
output(2, 250) <= input(39);
output(2, 251) <= input(38);
output(2, 252) <= input(35);
output(2, 253) <= input(36);
output(2, 254) <= input(32);
output(2, 255) <= input(0);
when "0111" =>
output(0, 0) <= input(0);
output(0, 1) <= input(1);
output(0, 2) <= input(2);
output(0, 3) <= input(3);
output(0, 4) <= input(4);
output(0, 5) <= input(5);
output(0, 6) <= input(6);
output(0, 7) <= input(7);
output(0, 8) <= input(8);
output(0, 9) <= input(9);
output(0, 10) <= input(10);
output(0, 11) <= input(11);
output(0, 12) <= input(12);
output(0, 13) <= input(13);
output(0, 14) <= input(14);
output(0, 15) <= input(15);
output(0, 16) <= input(16);
output(0, 17) <= input(0);
output(0, 18) <= input(1);
output(0, 19) <= input(2);
output(0, 20) <= input(3);
output(0, 21) <= input(4);
output(0, 22) <= input(5);
output(0, 23) <= input(6);
output(0, 24) <= input(7);
output(0, 25) <= input(8);
output(0, 26) <= input(9);
output(0, 27) <= input(10);
output(0, 28) <= input(11);
output(0, 29) <= input(12);
output(0, 30) <= input(13);
output(0, 31) <= input(14);
output(0, 32) <= input(17);
output(0, 33) <= input(16);
output(0, 34) <= input(0);
output(0, 35) <= input(1);
output(0, 36) <= input(2);
output(0, 37) <= input(3);
output(0, 38) <= input(4);
output(0, 39) <= input(5);
output(0, 40) <= input(6);
output(0, 41) <= input(7);
output(0, 42) <= input(8);
output(0, 43) <= input(9);
output(0, 44) <= input(10);
output(0, 45) <= input(11);
output(0, 46) <= input(12);
output(0, 47) <= input(13);
output(0, 48) <= input(18);
output(0, 49) <= input(17);
output(0, 50) <= input(16);
output(0, 51) <= input(0);
output(0, 52) <= input(1);
output(0, 53) <= input(2);
output(0, 54) <= input(3);
output(0, 55) <= input(4);
output(0, 56) <= input(5);
output(0, 57) <= input(6);
output(0, 58) <= input(7);
output(0, 59) <= input(8);
output(0, 60) <= input(9);
output(0, 61) <= input(10);
output(0, 62) <= input(11);
output(0, 63) <= input(12);
output(0, 64) <= input(19);
output(0, 65) <= input(18);
output(0, 66) <= input(17);
output(0, 67) <= input(16);
output(0, 68) <= input(0);
output(0, 69) <= input(1);
output(0, 70) <= input(2);
output(0, 71) <= input(3);
output(0, 72) <= input(4);
output(0, 73) <= input(5);
output(0, 74) <= input(6);
output(0, 75) <= input(7);
output(0, 76) <= input(8);
output(0, 77) <= input(9);
output(0, 78) <= input(10);
output(0, 79) <= input(11);
output(0, 80) <= input(20);
output(0, 81) <= input(21);
output(0, 82) <= input(22);
output(0, 83) <= input(23);
output(0, 84) <= input(24);
output(0, 85) <= input(25);
output(0, 86) <= input(26);
output(0, 87) <= input(27);
output(0, 88) <= input(28);
output(0, 89) <= input(29);
output(0, 90) <= input(30);
output(0, 91) <= input(31);
output(0, 92) <= input(32);
output(0, 93) <= input(33);
output(0, 94) <= input(34);
output(0, 95) <= input(35);
output(0, 96) <= input(36);
output(0, 97) <= input(20);
output(0, 98) <= input(21);
output(0, 99) <= input(22);
output(0, 100) <= input(23);
output(0, 101) <= input(24);
output(0, 102) <= input(25);
output(0, 103) <= input(26);
output(0, 104) <= input(27);
output(0, 105) <= input(28);
output(0, 106) <= input(29);
output(0, 107) <= input(30);
output(0, 108) <= input(31);
output(0, 109) <= input(32);
output(0, 110) <= input(33);
output(0, 111) <= input(34);
output(0, 112) <= input(37);
output(0, 113) <= input(36);
output(0, 114) <= input(20);
output(0, 115) <= input(21);
output(0, 116) <= input(22);
output(0, 117) <= input(23);
output(0, 118) <= input(24);
output(0, 119) <= input(25);
output(0, 120) <= input(26);
output(0, 121) <= input(27);
output(0, 122) <= input(28);
output(0, 123) <= input(29);
output(0, 124) <= input(30);
output(0, 125) <= input(31);
output(0, 126) <= input(32);
output(0, 127) <= input(33);
output(0, 128) <= input(38);
output(0, 129) <= input(37);
output(0, 130) <= input(36);
output(0, 131) <= input(20);
output(0, 132) <= input(21);
output(0, 133) <= input(22);
output(0, 134) <= input(23);
output(0, 135) <= input(24);
output(0, 136) <= input(25);
output(0, 137) <= input(26);
output(0, 138) <= input(27);
output(0, 139) <= input(28);
output(0, 140) <= input(29);
output(0, 141) <= input(30);
output(0, 142) <= input(31);
output(0, 143) <= input(32);
output(0, 144) <= input(39);
output(0, 145) <= input(38);
output(0, 146) <= input(37);
output(0, 147) <= input(36);
output(0, 148) <= input(20);
output(0, 149) <= input(21);
output(0, 150) <= input(22);
output(0, 151) <= input(23);
output(0, 152) <= input(24);
output(0, 153) <= input(25);
output(0, 154) <= input(26);
output(0, 155) <= input(27);
output(0, 156) <= input(28);
output(0, 157) <= input(29);
output(0, 158) <= input(30);
output(0, 159) <= input(31);
output(0, 160) <= input(40);
output(0, 161) <= input(41);
output(0, 162) <= input(42);
output(0, 163) <= input(43);
output(0, 164) <= input(44);
output(0, 165) <= input(19);
output(0, 166) <= input(18);
output(0, 167) <= input(17);
output(0, 168) <= input(16);
output(0, 169) <= input(0);
output(0, 170) <= input(1);
output(0, 171) <= input(2);
output(0, 172) <= input(3);
output(0, 173) <= input(4);
output(0, 174) <= input(5);
output(0, 175) <= input(6);
output(0, 176) <= input(45);
output(0, 177) <= input(40);
output(0, 178) <= input(41);
output(0, 179) <= input(42);
output(0, 180) <= input(43);
output(0, 181) <= input(44);
output(0, 182) <= input(19);
output(0, 183) <= input(18);
output(0, 184) <= input(17);
output(0, 185) <= input(16);
output(0, 186) <= input(0);
output(0, 187) <= input(1);
output(0, 188) <= input(2);
output(0, 189) <= input(3);
output(0, 190) <= input(4);
output(0, 191) <= input(5);
output(0, 192) <= input(46);
output(0, 193) <= input(45);
output(0, 194) <= input(40);
output(0, 195) <= input(41);
output(0, 196) <= input(42);
output(0, 197) <= input(43);
output(0, 198) <= input(44);
output(0, 199) <= input(19);
output(0, 200) <= input(18);
output(0, 201) <= input(17);
output(0, 202) <= input(16);
output(0, 203) <= input(0);
output(0, 204) <= input(1);
output(0, 205) <= input(2);
output(0, 206) <= input(3);
output(0, 207) <= input(4);
output(0, 208) <= input(47);
output(0, 209) <= input(46);
output(0, 210) <= input(45);
output(0, 211) <= input(40);
output(0, 212) <= input(41);
output(0, 213) <= input(42);
output(0, 214) <= input(43);
output(0, 215) <= input(44);
output(0, 216) <= input(19);
output(0, 217) <= input(18);
output(0, 218) <= input(17);
output(0, 219) <= input(16);
output(0, 220) <= input(0);
output(0, 221) <= input(1);
output(0, 222) <= input(2);
output(0, 223) <= input(3);
output(0, 224) <= input(48);
output(0, 225) <= input(47);
output(0, 226) <= input(46);
output(0, 227) <= input(45);
output(0, 228) <= input(40);
output(0, 229) <= input(41);
output(0, 230) <= input(42);
output(0, 231) <= input(43);
output(0, 232) <= input(44);
output(0, 233) <= input(19);
output(0, 234) <= input(18);
output(0, 235) <= input(17);
output(0, 236) <= input(16);
output(0, 237) <= input(0);
output(0, 238) <= input(1);
output(0, 239) <= input(2);
output(0, 240) <= input(49);
output(0, 241) <= input(50);
output(0, 242) <= input(51);
output(0, 243) <= input(52);
output(0, 244) <= input(53);
output(0, 245) <= input(39);
output(0, 246) <= input(38);
output(0, 247) <= input(37);
output(0, 248) <= input(36);
output(0, 249) <= input(20);
output(0, 250) <= input(21);
output(0, 251) <= input(22);
output(0, 252) <= input(23);
output(0, 253) <= input(24);
output(0, 254) <= input(25);
output(0, 255) <= input(26);
output(1, 0) <= input(54);
output(1, 1) <= input(55);
output(1, 2) <= input(56);
output(1, 3) <= input(57);
output(1, 4) <= input(58);
output(1, 5) <= input(59);
output(1, 6) <= input(60);
output(1, 7) <= input(61);
output(1, 8) <= input(62);
output(1, 9) <= input(63);
output(1, 10) <= input(64);
output(1, 11) <= input(65);
output(1, 12) <= input(66);
output(1, 13) <= input(67);
output(1, 14) <= input(68);
output(1, 15) <= input(69);
output(1, 16) <= input(70);
output(1, 17) <= input(54);
output(1, 18) <= input(55);
output(1, 19) <= input(56);
output(1, 20) <= input(57);
output(1, 21) <= input(58);
output(1, 22) <= input(59);
output(1, 23) <= input(60);
output(1, 24) <= input(61);
output(1, 25) <= input(62);
output(1, 26) <= input(63);
output(1, 27) <= input(64);
output(1, 28) <= input(65);
output(1, 29) <= input(66);
output(1, 30) <= input(67);
output(1, 31) <= input(68);
output(1, 32) <= input(71);
output(1, 33) <= input(70);
output(1, 34) <= input(54);
output(1, 35) <= input(55);
output(1, 36) <= input(56);
output(1, 37) <= input(57);
output(1, 38) <= input(58);
output(1, 39) <= input(59);
output(1, 40) <= input(60);
output(1, 41) <= input(61);
output(1, 42) <= input(62);
output(1, 43) <= input(63);
output(1, 44) <= input(64);
output(1, 45) <= input(65);
output(1, 46) <= input(66);
output(1, 47) <= input(67);
output(1, 48) <= input(72);
output(1, 49) <= input(71);
output(1, 50) <= input(70);
output(1, 51) <= input(54);
output(1, 52) <= input(55);
output(1, 53) <= input(56);
output(1, 54) <= input(57);
output(1, 55) <= input(58);
output(1, 56) <= input(59);
output(1, 57) <= input(60);
output(1, 58) <= input(61);
output(1, 59) <= input(62);
output(1, 60) <= input(63);
output(1, 61) <= input(64);
output(1, 62) <= input(65);
output(1, 63) <= input(66);
output(1, 64) <= input(73);
output(1, 65) <= input(72);
output(1, 66) <= input(71);
output(1, 67) <= input(70);
output(1, 68) <= input(54);
output(1, 69) <= input(55);
output(1, 70) <= input(56);
output(1, 71) <= input(57);
output(1, 72) <= input(58);
output(1, 73) <= input(59);
output(1, 74) <= input(60);
output(1, 75) <= input(61);
output(1, 76) <= input(62);
output(1, 77) <= input(63);
output(1, 78) <= input(64);
output(1, 79) <= input(65);
output(1, 80) <= input(74);
output(1, 81) <= input(73);
output(1, 82) <= input(72);
output(1, 83) <= input(71);
output(1, 84) <= input(70);
output(1, 85) <= input(54);
output(1, 86) <= input(55);
output(1, 87) <= input(56);
output(1, 88) <= input(57);
output(1, 89) <= input(58);
output(1, 90) <= input(59);
output(1, 91) <= input(60);
output(1, 92) <= input(61);
output(1, 93) <= input(62);
output(1, 94) <= input(63);
output(1, 95) <= input(64);
output(1, 96) <= input(75);
output(1, 97) <= input(74);
output(1, 98) <= input(73);
output(1, 99) <= input(72);
output(1, 100) <= input(71);
output(1, 101) <= input(70);
output(1, 102) <= input(54);
output(1, 103) <= input(55);
output(1, 104) <= input(56);
output(1, 105) <= input(57);
output(1, 106) <= input(58);
output(1, 107) <= input(59);
output(1, 108) <= input(60);
output(1, 109) <= input(61);
output(1, 110) <= input(62);
output(1, 111) <= input(63);
output(1, 112) <= input(76);
output(1, 113) <= input(75);
output(1, 114) <= input(74);
output(1, 115) <= input(73);
output(1, 116) <= input(72);
output(1, 117) <= input(71);
output(1, 118) <= input(70);
output(1, 119) <= input(54);
output(1, 120) <= input(55);
output(1, 121) <= input(56);
output(1, 122) <= input(57);
output(1, 123) <= input(58);
output(1, 124) <= input(59);
output(1, 125) <= input(60);
output(1, 126) <= input(61);
output(1, 127) <= input(62);
output(1, 128) <= input(77);
output(1, 129) <= input(76);
output(1, 130) <= input(75);
output(1, 131) <= input(74);
output(1, 132) <= input(73);
output(1, 133) <= input(72);
output(1, 134) <= input(71);
output(1, 135) <= input(70);
output(1, 136) <= input(54);
output(1, 137) <= input(55);
output(1, 138) <= input(56);
output(1, 139) <= input(57);
output(1, 140) <= input(58);
output(1, 141) <= input(59);
output(1, 142) <= input(60);
output(1, 143) <= input(61);
output(1, 144) <= input(78);
output(1, 145) <= input(77);
output(1, 146) <= input(76);
output(1, 147) <= input(75);
output(1, 148) <= input(74);
output(1, 149) <= input(73);
output(1, 150) <= input(72);
output(1, 151) <= input(71);
output(1, 152) <= input(70);
output(1, 153) <= input(54);
output(1, 154) <= input(55);
output(1, 155) <= input(56);
output(1, 156) <= input(57);
output(1, 157) <= input(58);
output(1, 158) <= input(59);
output(1, 159) <= input(60);
output(1, 160) <= input(79);
output(1, 161) <= input(78);
output(1, 162) <= input(77);
output(1, 163) <= input(76);
output(1, 164) <= input(75);
output(1, 165) <= input(74);
output(1, 166) <= input(73);
output(1, 167) <= input(72);
output(1, 168) <= input(71);
output(1, 169) <= input(70);
output(1, 170) <= input(54);
output(1, 171) <= input(55);
output(1, 172) <= input(56);
output(1, 173) <= input(57);
output(1, 174) <= input(58);
output(1, 175) <= input(59);
output(1, 176) <= input(80);
output(1, 177) <= input(79);
output(1, 178) <= input(78);
output(1, 179) <= input(77);
output(1, 180) <= input(76);
output(1, 181) <= input(75);
output(1, 182) <= input(74);
output(1, 183) <= input(73);
output(1, 184) <= input(72);
output(1, 185) <= input(71);
output(1, 186) <= input(70);
output(1, 187) <= input(54);
output(1, 188) <= input(55);
output(1, 189) <= input(56);
output(1, 190) <= input(57);
output(1, 191) <= input(58);
output(1, 192) <= input(81);
output(1, 193) <= input(80);
output(1, 194) <= input(79);
output(1, 195) <= input(78);
output(1, 196) <= input(77);
output(1, 197) <= input(76);
output(1, 198) <= input(75);
output(1, 199) <= input(74);
output(1, 200) <= input(73);
output(1, 201) <= input(72);
output(1, 202) <= input(71);
output(1, 203) <= input(70);
output(1, 204) <= input(54);
output(1, 205) <= input(55);
output(1, 206) <= input(56);
output(1, 207) <= input(57);
output(1, 208) <= input(82);
output(1, 209) <= input(81);
output(1, 210) <= input(80);
output(1, 211) <= input(79);
output(1, 212) <= input(78);
output(1, 213) <= input(77);
output(1, 214) <= input(76);
output(1, 215) <= input(75);
output(1, 216) <= input(74);
output(1, 217) <= input(73);
output(1, 218) <= input(72);
output(1, 219) <= input(71);
output(1, 220) <= input(70);
output(1, 221) <= input(54);
output(1, 222) <= input(55);
output(1, 223) <= input(56);
output(1, 224) <= input(83);
output(1, 225) <= input(82);
output(1, 226) <= input(81);
output(1, 227) <= input(80);
output(1, 228) <= input(79);
output(1, 229) <= input(78);
output(1, 230) <= input(77);
output(1, 231) <= input(76);
output(1, 232) <= input(75);
output(1, 233) <= input(74);
output(1, 234) <= input(73);
output(1, 235) <= input(72);
output(1, 236) <= input(71);
output(1, 237) <= input(70);
output(1, 238) <= input(54);
output(1, 239) <= input(55);
output(1, 240) <= input(84);
output(1, 241) <= input(83);
output(1, 242) <= input(82);
output(1, 243) <= input(81);
output(1, 244) <= input(80);
output(1, 245) <= input(79);
output(1, 246) <= input(78);
output(1, 247) <= input(77);
output(1, 248) <= input(76);
output(1, 249) <= input(75);
output(1, 250) <= input(74);
output(1, 251) <= input(73);
output(1, 252) <= input(72);
output(1, 253) <= input(71);
output(1, 254) <= input(70);
output(1, 255) <= input(54);
when "1000" =>
output(0, 0) <= input(0);
output(0, 1) <= input(1);
output(0, 2) <= input(2);
output(0, 3) <= input(3);
output(0, 4) <= input(4);
output(0, 5) <= input(5);
output(0, 6) <= input(6);
output(0, 7) <= input(7);
output(0, 8) <= input(8);
output(0, 9) <= input(9);
output(0, 10) <= input(10);
output(0, 11) <= input(11);
output(0, 12) <= input(12);
output(0, 13) <= input(13);
output(0, 14) <= input(14);
output(0, 15) <= input(15);
output(0, 16) <= input(16);
output(0, 17) <= input(0);
output(0, 18) <= input(1);
output(0, 19) <= input(2);
output(0, 20) <= input(3);
output(0, 21) <= input(4);
output(0, 22) <= input(5);
output(0, 23) <= input(6);
output(0, 24) <= input(7);
output(0, 25) <= input(8);
output(0, 26) <= input(9);
output(0, 27) <= input(10);
output(0, 28) <= input(11);
output(0, 29) <= input(12);
output(0, 30) <= input(13);
output(0, 31) <= input(14);
output(0, 32) <= input(17);
output(0, 33) <= input(16);
output(0, 34) <= input(0);
output(0, 35) <= input(1);
output(0, 36) <= input(2);
output(0, 37) <= input(3);
output(0, 38) <= input(4);
output(0, 39) <= input(5);
output(0, 40) <= input(6);
output(0, 41) <= input(7);
output(0, 42) <= input(8);
output(0, 43) <= input(9);
output(0, 44) <= input(10);
output(0, 45) <= input(11);
output(0, 46) <= input(12);
output(0, 47) <= input(13);
output(0, 48) <= input(18);
output(0, 49) <= input(17);
output(0, 50) <= input(16);
output(0, 51) <= input(0);
output(0, 52) <= input(1);
output(0, 53) <= input(2);
output(0, 54) <= input(3);
output(0, 55) <= input(4);
output(0, 56) <= input(5);
output(0, 57) <= input(6);
output(0, 58) <= input(7);
output(0, 59) <= input(8);
output(0, 60) <= input(9);
output(0, 61) <= input(10);
output(0, 62) <= input(11);
output(0, 63) <= input(12);
output(0, 64) <= input(19);
output(0, 65) <= input(18);
output(0, 66) <= input(17);
output(0, 67) <= input(16);
output(0, 68) <= input(0);
output(0, 69) <= input(1);
output(0, 70) <= input(2);
output(0, 71) <= input(3);
output(0, 72) <= input(4);
output(0, 73) <= input(5);
output(0, 74) <= input(6);
output(0, 75) <= input(7);
output(0, 76) <= input(8);
output(0, 77) <= input(9);
output(0, 78) <= input(10);
output(0, 79) <= input(11);
output(0, 80) <= input(20);
output(0, 81) <= input(21);
output(0, 82) <= input(22);
output(0, 83) <= input(23);
output(0, 84) <= input(24);
output(0, 85) <= input(25);
output(0, 86) <= input(26);
output(0, 87) <= input(27);
output(0, 88) <= input(28);
output(0, 89) <= input(29);
output(0, 90) <= input(30);
output(0, 91) <= input(31);
output(0, 92) <= input(32);
output(0, 93) <= input(33);
output(0, 94) <= input(34);
output(0, 95) <= input(35);
output(0, 96) <= input(36);
output(0, 97) <= input(20);
output(0, 98) <= input(21);
output(0, 99) <= input(22);
output(0, 100) <= input(23);
output(0, 101) <= input(24);
output(0, 102) <= input(25);
output(0, 103) <= input(26);
output(0, 104) <= input(27);
output(0, 105) <= input(28);
output(0, 106) <= input(29);
output(0, 107) <= input(30);
output(0, 108) <= input(31);
output(0, 109) <= input(32);
output(0, 110) <= input(33);
output(0, 111) <= input(34);
output(0, 112) <= input(37);
output(0, 113) <= input(36);
output(0, 114) <= input(20);
output(0, 115) <= input(21);
output(0, 116) <= input(22);
output(0, 117) <= input(23);
output(0, 118) <= input(24);
output(0, 119) <= input(25);
output(0, 120) <= input(26);
output(0, 121) <= input(27);
output(0, 122) <= input(28);
output(0, 123) <= input(29);
output(0, 124) <= input(30);
output(0, 125) <= input(31);
output(0, 126) <= input(32);
output(0, 127) <= input(33);
output(0, 128) <= input(38);
output(0, 129) <= input(37);
output(0, 130) <= input(36);
output(0, 131) <= input(20);
output(0, 132) <= input(21);
output(0, 133) <= input(22);
output(0, 134) <= input(23);
output(0, 135) <= input(24);
output(0, 136) <= input(25);
output(0, 137) <= input(26);
output(0, 138) <= input(27);
output(0, 139) <= input(28);
output(0, 140) <= input(29);
output(0, 141) <= input(30);
output(0, 142) <= input(31);
output(0, 143) <= input(32);
output(0, 144) <= input(39);
output(0, 145) <= input(38);
output(0, 146) <= input(37);
output(0, 147) <= input(36);
output(0, 148) <= input(20);
output(0, 149) <= input(21);
output(0, 150) <= input(22);
output(0, 151) <= input(23);
output(0, 152) <= input(24);
output(0, 153) <= input(25);
output(0, 154) <= input(26);
output(0, 155) <= input(27);
output(0, 156) <= input(28);
output(0, 157) <= input(29);
output(0, 158) <= input(30);
output(0, 159) <= input(31);
output(0, 160) <= input(40);
output(0, 161) <= input(41);
output(0, 162) <= input(42);
output(0, 163) <= input(43);
output(0, 164) <= input(44);
output(0, 165) <= input(19);
output(0, 166) <= input(18);
output(0, 167) <= input(17);
output(0, 168) <= input(16);
output(0, 169) <= input(0);
output(0, 170) <= input(1);
output(0, 171) <= input(2);
output(0, 172) <= input(3);
output(0, 173) <= input(4);
output(0, 174) <= input(5);
output(0, 175) <= input(6);
output(0, 176) <= input(45);
output(0, 177) <= input(40);
output(0, 178) <= input(41);
output(0, 179) <= input(42);
output(0, 180) <= input(43);
output(0, 181) <= input(44);
output(0, 182) <= input(19);
output(0, 183) <= input(18);
output(0, 184) <= input(17);
output(0, 185) <= input(16);
output(0, 186) <= input(0);
output(0, 187) <= input(1);
output(0, 188) <= input(2);
output(0, 189) <= input(3);
output(0, 190) <= input(4);
output(0, 191) <= input(5);
output(0, 192) <= input(46);
output(0, 193) <= input(45);
output(0, 194) <= input(40);
output(0, 195) <= input(41);
output(0, 196) <= input(42);
output(0, 197) <= input(43);
output(0, 198) <= input(44);
output(0, 199) <= input(19);
output(0, 200) <= input(18);
output(0, 201) <= input(17);
output(0, 202) <= input(16);
output(0, 203) <= input(0);
output(0, 204) <= input(1);
output(0, 205) <= input(2);
output(0, 206) <= input(3);
output(0, 207) <= input(4);
output(0, 208) <= input(47);
output(0, 209) <= input(46);
output(0, 210) <= input(45);
output(0, 211) <= input(40);
output(0, 212) <= input(41);
output(0, 213) <= input(42);
output(0, 214) <= input(43);
output(0, 215) <= input(44);
output(0, 216) <= input(19);
output(0, 217) <= input(18);
output(0, 218) <= input(17);
output(0, 219) <= input(16);
output(0, 220) <= input(0);
output(0, 221) <= input(1);
output(0, 222) <= input(2);
output(0, 223) <= input(3);
output(0, 224) <= input(48);
output(0, 225) <= input(47);
output(0, 226) <= input(46);
output(0, 227) <= input(45);
output(0, 228) <= input(40);
output(0, 229) <= input(41);
output(0, 230) <= input(42);
output(0, 231) <= input(43);
output(0, 232) <= input(44);
output(0, 233) <= input(19);
output(0, 234) <= input(18);
output(0, 235) <= input(17);
output(0, 236) <= input(16);
output(0, 237) <= input(0);
output(0, 238) <= input(1);
output(0, 239) <= input(2);
output(0, 240) <= input(49);
output(0, 241) <= input(50);
output(0, 242) <= input(51);
output(0, 243) <= input(52);
output(0, 244) <= input(53);
output(0, 245) <= input(39);
output(0, 246) <= input(38);
output(0, 247) <= input(37);
output(0, 248) <= input(36);
output(0, 249) <= input(20);
output(0, 250) <= input(21);
output(0, 251) <= input(22);
output(0, 252) <= input(23);
output(0, 253) <= input(24);
output(0, 254) <= input(25);
output(0, 255) <= input(26);
when "1001" =>
output(0, 0) <= input(0);
output(0, 1) <= input(1);
output(0, 2) <= input(2);
output(0, 3) <= input(3);
output(0, 4) <= input(4);
output(0, 5) <= input(5);
output(0, 6) <= input(6);
output(0, 7) <= input(7);
output(0, 8) <= input(8);
output(0, 9) <= input(9);
output(0, 10) <= input(10);
output(0, 11) <= input(11);
output(0, 12) <= input(12);
output(0, 13) <= input(13);
output(0, 14) <= input(14);
output(0, 15) <= input(15);
output(0, 16) <= input(16);
output(0, 17) <= input(0);
output(0, 18) <= input(1);
output(0, 19) <= input(2);
output(0, 20) <= input(3);
output(0, 21) <= input(4);
output(0, 22) <= input(5);
output(0, 23) <= input(6);
output(0, 24) <= input(7);
output(0, 25) <= input(8);
output(0, 26) <= input(9);
output(0, 27) <= input(10);
output(0, 28) <= input(11);
output(0, 29) <= input(12);
output(0, 30) <= input(13);
output(0, 31) <= input(14);
output(0, 32) <= input(17);
output(0, 33) <= input(18);
output(0, 34) <= input(19);
output(0, 35) <= input(20);
output(0, 36) <= input(21);
output(0, 37) <= input(22);
output(0, 38) <= input(23);
output(0, 39) <= input(24);
output(0, 40) <= input(25);
output(0, 41) <= input(26);
output(0, 42) <= input(27);
output(0, 43) <= input(28);
output(0, 44) <= input(29);
output(0, 45) <= input(30);
output(0, 46) <= input(31);
output(0, 47) <= input(32);
output(0, 48) <= input(33);
output(0, 49) <= input(17);
output(0, 50) <= input(18);
output(0, 51) <= input(19);
output(0, 52) <= input(20);
output(0, 53) <= input(21);
output(0, 54) <= input(22);
output(0, 55) <= input(23);
output(0, 56) <= input(24);
output(0, 57) <= input(25);
output(0, 58) <= input(26);
output(0, 59) <= input(27);
output(0, 60) <= input(28);
output(0, 61) <= input(29);
output(0, 62) <= input(30);
output(0, 63) <= input(31);
output(0, 64) <= input(34);
output(0, 65) <= input(33);
output(0, 66) <= input(17);
output(0, 67) <= input(18);
output(0, 68) <= input(19);
output(0, 69) <= input(20);
output(0, 70) <= input(21);
output(0, 71) <= input(22);
output(0, 72) <= input(23);
output(0, 73) <= input(24);
output(0, 74) <= input(25);
output(0, 75) <= input(26);
output(0, 76) <= input(27);
output(0, 77) <= input(28);
output(0, 78) <= input(29);
output(0, 79) <= input(30);
output(0, 80) <= input(35);
output(0, 81) <= input(36);
output(0, 82) <= input(37);
output(0, 83) <= input(16);
output(0, 84) <= input(0);
output(0, 85) <= input(1);
output(0, 86) <= input(2);
output(0, 87) <= input(3);
output(0, 88) <= input(4);
output(0, 89) <= input(5);
output(0, 90) <= input(6);
output(0, 91) <= input(7);
output(0, 92) <= input(8);
output(0, 93) <= input(9);
output(0, 94) <= input(10);
output(0, 95) <= input(11);
output(0, 96) <= input(38);
output(0, 97) <= input(35);
output(0, 98) <= input(36);
output(0, 99) <= input(37);
output(0, 100) <= input(16);
output(0, 101) <= input(0);
output(0, 102) <= input(1);
output(0, 103) <= input(2);
output(0, 104) <= input(3);
output(0, 105) <= input(4);
output(0, 106) <= input(5);
output(0, 107) <= input(6);
output(0, 108) <= input(7);
output(0, 109) <= input(8);
output(0, 110) <= input(9);
output(0, 111) <= input(10);
output(0, 112) <= input(39);
output(0, 113) <= input(40);
output(0, 114) <= input(34);
output(0, 115) <= input(33);
output(0, 116) <= input(17);
output(0, 117) <= input(18);
output(0, 118) <= input(19);
output(0, 119) <= input(20);
output(0, 120) <= input(21);
output(0, 121) <= input(22);
output(0, 122) <= input(23);
output(0, 123) <= input(24);
output(0, 124) <= input(25);
output(0, 125) <= input(26);
output(0, 126) <= input(27);
output(0, 127) <= input(28);
output(0, 128) <= input(41);
output(0, 129) <= input(39);
output(0, 130) <= input(40);
output(0, 131) <= input(34);
output(0, 132) <= input(33);
output(0, 133) <= input(17);
output(0, 134) <= input(18);
output(0, 135) <= input(19);
output(0, 136) <= input(20);
output(0, 137) <= input(21);
output(0, 138) <= input(22);
output(0, 139) <= input(23);
output(0, 140) <= input(24);
output(0, 141) <= input(25);
output(0, 142) <= input(26);
output(0, 143) <= input(27);
output(0, 144) <= input(42);
output(0, 145) <= input(41);
output(0, 146) <= input(39);
output(0, 147) <= input(40);
output(0, 148) <= input(34);
output(0, 149) <= input(33);
output(0, 150) <= input(17);
output(0, 151) <= input(18);
output(0, 152) <= input(19);
output(0, 153) <= input(20);
output(0, 154) <= input(21);
output(0, 155) <= input(22);
output(0, 156) <= input(23);
output(0, 157) <= input(24);
output(0, 158) <= input(25);
output(0, 159) <= input(26);
output(0, 160) <= input(43);
output(0, 161) <= input(44);
output(0, 162) <= input(45);
output(0, 163) <= input(38);
output(0, 164) <= input(35);
output(0, 165) <= input(36);
output(0, 166) <= input(37);
output(0, 167) <= input(16);
output(0, 168) <= input(0);
output(0, 169) <= input(1);
output(0, 170) <= input(2);
output(0, 171) <= input(3);
output(0, 172) <= input(4);
output(0, 173) <= input(5);
output(0, 174) <= input(6);
output(0, 175) <= input(7);
output(0, 176) <= input(46);
output(0, 177) <= input(43);
output(0, 178) <= input(44);
output(0, 179) <= input(45);
output(0, 180) <= input(38);
output(0, 181) <= input(35);
output(0, 182) <= input(36);
output(0, 183) <= input(37);
output(0, 184) <= input(16);
output(0, 185) <= input(0);
output(0, 186) <= input(1);
output(0, 187) <= input(2);
output(0, 188) <= input(3);
output(0, 189) <= input(4);
output(0, 190) <= input(5);
output(0, 191) <= input(6);
output(0, 192) <= input(47);
output(0, 193) <= input(46);
output(0, 194) <= input(43);
output(0, 195) <= input(44);
output(0, 196) <= input(45);
output(0, 197) <= input(38);
output(0, 198) <= input(35);
output(0, 199) <= input(36);
output(0, 200) <= input(37);
output(0, 201) <= input(16);
output(0, 202) <= input(0);
output(0, 203) <= input(1);
output(0, 204) <= input(2);
output(0, 205) <= input(3);
output(0, 206) <= input(4);
output(0, 207) <= input(5);
output(0, 208) <= input(48);
output(0, 209) <= input(49);
output(0, 210) <= input(50);
output(0, 211) <= input(42);
output(0, 212) <= input(41);
output(0, 213) <= input(39);
output(0, 214) <= input(40);
output(0, 215) <= input(34);
output(0, 216) <= input(33);
output(0, 217) <= input(17);
output(0, 218) <= input(18);
output(0, 219) <= input(19);
output(0, 220) <= input(20);
output(0, 221) <= input(21);
output(0, 222) <= input(22);
output(0, 223) <= input(23);
output(0, 224) <= input(51);
output(0, 225) <= input(48);
output(0, 226) <= input(49);
output(0, 227) <= input(50);
output(0, 228) <= input(42);
output(0, 229) <= input(41);
output(0, 230) <= input(39);
output(0, 231) <= input(40);
output(0, 232) <= input(34);
output(0, 233) <= input(33);
output(0, 234) <= input(17);
output(0, 235) <= input(18);
output(0, 236) <= input(19);
output(0, 237) <= input(20);
output(0, 238) <= input(21);
output(0, 239) <= input(22);
output(0, 240) <= input(52);
output(0, 241) <= input(53);
output(0, 242) <= input(47);
output(0, 243) <= input(46);
output(0, 244) <= input(43);
output(0, 245) <= input(44);
output(0, 246) <= input(45);
output(0, 247) <= input(38);
output(0, 248) <= input(35);
output(0, 249) <= input(36);
output(0, 250) <= input(37);
output(0, 251) <= input(16);
output(0, 252) <= input(0);
output(0, 253) <= input(1);
output(0, 254) <= input(2);
output(0, 255) <= input(3);
output(1, 0) <= input(20);
output(1, 1) <= input(21);
output(1, 2) <= input(22);
output(1, 3) <= input(23);
output(1, 4) <= input(24);
output(1, 5) <= input(25);
output(1, 6) <= input(26);
output(1, 7) <= input(27);
output(1, 8) <= input(28);
output(1, 9) <= input(29);
output(1, 10) <= input(30);
output(1, 11) <= input(31);
output(1, 12) <= input(32);
output(1, 13) <= input(54);
output(1, 14) <= input(55);
output(1, 15) <= input(56);
output(1, 16) <= input(1);
output(1, 17) <= input(2);
output(1, 18) <= input(3);
output(1, 19) <= input(4);
output(1, 20) <= input(5);
output(1, 21) <= input(6);
output(1, 22) <= input(7);
output(1, 23) <= input(8);
output(1, 24) <= input(9);
output(1, 25) <= input(10);
output(1, 26) <= input(11);
output(1, 27) <= input(12);
output(1, 28) <= input(13);
output(1, 29) <= input(14);
output(1, 30) <= input(15);
output(1, 31) <= input(57);
output(1, 32) <= input(0);
output(1, 33) <= input(1);
output(1, 34) <= input(2);
output(1, 35) <= input(3);
output(1, 36) <= input(4);
output(1, 37) <= input(5);
output(1, 38) <= input(6);
output(1, 39) <= input(7);
output(1, 40) <= input(8);
output(1, 41) <= input(9);
output(1, 42) <= input(10);
output(1, 43) <= input(11);
output(1, 44) <= input(12);
output(1, 45) <= input(13);
output(1, 46) <= input(14);
output(1, 47) <= input(15);
output(1, 48) <= input(18);
output(1, 49) <= input(19);
output(1, 50) <= input(20);
output(1, 51) <= input(21);
output(1, 52) <= input(22);
output(1, 53) <= input(23);
output(1, 54) <= input(24);
output(1, 55) <= input(25);
output(1, 56) <= input(26);
output(1, 57) <= input(27);
output(1, 58) <= input(28);
output(1, 59) <= input(29);
output(1, 60) <= input(30);
output(1, 61) <= input(31);
output(1, 62) <= input(32);
output(1, 63) <= input(54);
output(1, 64) <= input(17);
output(1, 65) <= input(18);
output(1, 66) <= input(19);
output(1, 67) <= input(20);
output(1, 68) <= input(21);
output(1, 69) <= input(22);
output(1, 70) <= input(23);
output(1, 71) <= input(24);
output(1, 72) <= input(25);
output(1, 73) <= input(26);
output(1, 74) <= input(27);
output(1, 75) <= input(28);
output(1, 76) <= input(29);
output(1, 77) <= input(30);
output(1, 78) <= input(31);
output(1, 79) <= input(32);
output(1, 80) <= input(37);
output(1, 81) <= input(16);
output(1, 82) <= input(0);
output(1, 83) <= input(1);
output(1, 84) <= input(2);
output(1, 85) <= input(3);
output(1, 86) <= input(4);
output(1, 87) <= input(5);
output(1, 88) <= input(6);
output(1, 89) <= input(7);
output(1, 90) <= input(8);
output(1, 91) <= input(9);
output(1, 92) <= input(10);
output(1, 93) <= input(11);
output(1, 94) <= input(12);
output(1, 95) <= input(13);
output(1, 96) <= input(36);
output(1, 97) <= input(37);
output(1, 98) <= input(16);
output(1, 99) <= input(0);
output(1, 100) <= input(1);
output(1, 101) <= input(2);
output(1, 102) <= input(3);
output(1, 103) <= input(4);
output(1, 104) <= input(5);
output(1, 105) <= input(6);
output(1, 106) <= input(7);
output(1, 107) <= input(8);
output(1, 108) <= input(9);
output(1, 109) <= input(10);
output(1, 110) <= input(11);
output(1, 111) <= input(12);
output(1, 112) <= input(58);
output(1, 113) <= input(33);
output(1, 114) <= input(17);
output(1, 115) <= input(18);
output(1, 116) <= input(19);
output(1, 117) <= input(20);
output(1, 118) <= input(21);
output(1, 119) <= input(22);
output(1, 120) <= input(23);
output(1, 121) <= input(24);
output(1, 122) <= input(25);
output(1, 123) <= input(26);
output(1, 124) <= input(27);
output(1, 125) <= input(28);
output(1, 126) <= input(29);
output(1, 127) <= input(30);
output(1, 128) <= input(59);
output(1, 129) <= input(36);
output(1, 130) <= input(37);
output(1, 131) <= input(16);
output(1, 132) <= input(0);
output(1, 133) <= input(1);
output(1, 134) <= input(2);
output(1, 135) <= input(3);
output(1, 136) <= input(4);
output(1, 137) <= input(5);
output(1, 138) <= input(6);
output(1, 139) <= input(7);
output(1, 140) <= input(8);
output(1, 141) <= input(9);
output(1, 142) <= input(10);
output(1, 143) <= input(11);
output(1, 144) <= input(60);
output(1, 145) <= input(59);
output(1, 146) <= input(36);
output(1, 147) <= input(37);
output(1, 148) <= input(16);
output(1, 149) <= input(0);
output(1, 150) <= input(1);
output(1, 151) <= input(2);
output(1, 152) <= input(3);
output(1, 153) <= input(4);
output(1, 154) <= input(5);
output(1, 155) <= input(6);
output(1, 156) <= input(7);
output(1, 157) <= input(8);
output(1, 158) <= input(9);
output(1, 159) <= input(10);
output(1, 160) <= input(61);
output(1, 161) <= input(62);
output(1, 162) <= input(58);
output(1, 163) <= input(33);
output(1, 164) <= input(17);
output(1, 165) <= input(18);
output(1, 166) <= input(19);
output(1, 167) <= input(20);
output(1, 168) <= input(21);
output(1, 169) <= input(22);
output(1, 170) <= input(23);
output(1, 171) <= input(24);
output(1, 172) <= input(25);
output(1, 173) <= input(26);
output(1, 174) <= input(27);
output(1, 175) <= input(28);
output(1, 176) <= input(63);
output(1, 177) <= input(61);
output(1, 178) <= input(62);
output(1, 179) <= input(58);
output(1, 180) <= input(33);
output(1, 181) <= input(17);
output(1, 182) <= input(18);
output(1, 183) <= input(19);
output(1, 184) <= input(20);
output(1, 185) <= input(21);
output(1, 186) <= input(22);
output(1, 187) <= input(23);
output(1, 188) <= input(24);
output(1, 189) <= input(25);
output(1, 190) <= input(26);
output(1, 191) <= input(27);
output(1, 192) <= input(64);
output(1, 193) <= input(65);
output(1, 194) <= input(60);
output(1, 195) <= input(59);
output(1, 196) <= input(36);
output(1, 197) <= input(37);
output(1, 198) <= input(16);
output(1, 199) <= input(0);
output(1, 200) <= input(1);
output(1, 201) <= input(2);
output(1, 202) <= input(3);
output(1, 203) <= input(4);
output(1, 204) <= input(5);
output(1, 205) <= input(6);
output(1, 206) <= input(7);
output(1, 207) <= input(8);
output(1, 208) <= input(66);
output(1, 209) <= input(64);
output(1, 210) <= input(65);
output(1, 211) <= input(60);
output(1, 212) <= input(59);
output(1, 213) <= input(36);
output(1, 214) <= input(37);
output(1, 215) <= input(16);
output(1, 216) <= input(0);
output(1, 217) <= input(1);
output(1, 218) <= input(2);
output(1, 219) <= input(3);
output(1, 220) <= input(4);
output(1, 221) <= input(5);
output(1, 222) <= input(6);
output(1, 223) <= input(7);
output(1, 224) <= input(67);
output(1, 225) <= input(68);
output(1, 226) <= input(63);
output(1, 227) <= input(61);
output(1, 228) <= input(62);
output(1, 229) <= input(58);
output(1, 230) <= input(33);
output(1, 231) <= input(17);
output(1, 232) <= input(18);
output(1, 233) <= input(19);
output(1, 234) <= input(20);
output(1, 235) <= input(21);
output(1, 236) <= input(22);
output(1, 237) <= input(23);
output(1, 238) <= input(24);
output(1, 239) <= input(25);
output(1, 240) <= input(69);
output(1, 241) <= input(66);
output(1, 242) <= input(64);
output(1, 243) <= input(65);
output(1, 244) <= input(60);
output(1, 245) <= input(59);
output(1, 246) <= input(36);
output(1, 247) <= input(37);
output(1, 248) <= input(16);
output(1, 249) <= input(0);
output(1, 250) <= input(1);
output(1, 251) <= input(2);
output(1, 252) <= input(3);
output(1, 253) <= input(4);
output(1, 254) <= input(5);
output(1, 255) <= input(6);
output(2, 0) <= input(3);
output(2, 1) <= input(4);
output(2, 2) <= input(5);
output(2, 3) <= input(6);
output(2, 4) <= input(7);
output(2, 5) <= input(8);
output(2, 6) <= input(9);
output(2, 7) <= input(10);
output(2, 8) <= input(11);
output(2, 9) <= input(12);
output(2, 10) <= input(13);
output(2, 11) <= input(14);
output(2, 12) <= input(15);
output(2, 13) <= input(57);
output(2, 14) <= input(70);
output(2, 15) <= input(71);
output(2, 16) <= input(21);
output(2, 17) <= input(22);
output(2, 18) <= input(23);
output(2, 19) <= input(24);
output(2, 20) <= input(25);
output(2, 21) <= input(26);
output(2, 22) <= input(27);
output(2, 23) <= input(28);
output(2, 24) <= input(29);
output(2, 25) <= input(30);
output(2, 26) <= input(31);
output(2, 27) <= input(32);
output(2, 28) <= input(54);
output(2, 29) <= input(55);
output(2, 30) <= input(56);
output(2, 31) <= input(72);
output(2, 32) <= input(2);
output(2, 33) <= input(3);
output(2, 34) <= input(4);
output(2, 35) <= input(5);
output(2, 36) <= input(6);
output(2, 37) <= input(7);
output(2, 38) <= input(8);
output(2, 39) <= input(9);
output(2, 40) <= input(10);
output(2, 41) <= input(11);
output(2, 42) <= input(12);
output(2, 43) <= input(13);
output(2, 44) <= input(14);
output(2, 45) <= input(15);
output(2, 46) <= input(57);
output(2, 47) <= input(70);
output(2, 48) <= input(20);
output(2, 49) <= input(21);
output(2, 50) <= input(22);
output(2, 51) <= input(23);
output(2, 52) <= input(24);
output(2, 53) <= input(25);
output(2, 54) <= input(26);
output(2, 55) <= input(27);
output(2, 56) <= input(28);
output(2, 57) <= input(29);
output(2, 58) <= input(30);
output(2, 59) <= input(31);
output(2, 60) <= input(32);
output(2, 61) <= input(54);
output(2, 62) <= input(55);
output(2, 63) <= input(56);
output(2, 64) <= input(19);
output(2, 65) <= input(20);
output(2, 66) <= input(21);
output(2, 67) <= input(22);
output(2, 68) <= input(23);
output(2, 69) <= input(24);
output(2, 70) <= input(25);
output(2, 71) <= input(26);
output(2, 72) <= input(27);
output(2, 73) <= input(28);
output(2, 74) <= input(29);
output(2, 75) <= input(30);
output(2, 76) <= input(31);
output(2, 77) <= input(32);
output(2, 78) <= input(54);
output(2, 79) <= input(55);
output(2, 80) <= input(0);
output(2, 81) <= input(1);
output(2, 82) <= input(2);
output(2, 83) <= input(3);
output(2, 84) <= input(4);
output(2, 85) <= input(5);
output(2, 86) <= input(6);
output(2, 87) <= input(7);
output(2, 88) <= input(8);
output(2, 89) <= input(9);
output(2, 90) <= input(10);
output(2, 91) <= input(11);
output(2, 92) <= input(12);
output(2, 93) <= input(13);
output(2, 94) <= input(14);
output(2, 95) <= input(15);
output(2, 96) <= input(18);
output(2, 97) <= input(19);
output(2, 98) <= input(20);
output(2, 99) <= input(21);
output(2, 100) <= input(22);
output(2, 101) <= input(23);
output(2, 102) <= input(24);
output(2, 103) <= input(25);
output(2, 104) <= input(26);
output(2, 105) <= input(27);
output(2, 106) <= input(28);
output(2, 107) <= input(29);
output(2, 108) <= input(30);
output(2, 109) <= input(31);
output(2, 110) <= input(32);
output(2, 111) <= input(54);
output(2, 112) <= input(16);
output(2, 113) <= input(0);
output(2, 114) <= input(1);
output(2, 115) <= input(2);
output(2, 116) <= input(3);
output(2, 117) <= input(4);
output(2, 118) <= input(5);
output(2, 119) <= input(6);
output(2, 120) <= input(7);
output(2, 121) <= input(8);
output(2, 122) <= input(9);
output(2, 123) <= input(10);
output(2, 124) <= input(11);
output(2, 125) <= input(12);
output(2, 126) <= input(13);
output(2, 127) <= input(14);
output(2, 128) <= input(37);
output(2, 129) <= input(16);
output(2, 130) <= input(0);
output(2, 131) <= input(1);
output(2, 132) <= input(2);
output(2, 133) <= input(3);
output(2, 134) <= input(4);
output(2, 135) <= input(5);
output(2, 136) <= input(6);
output(2, 137) <= input(7);
output(2, 138) <= input(8);
output(2, 139) <= input(9);
output(2, 140) <= input(10);
output(2, 141) <= input(11);
output(2, 142) <= input(12);
output(2, 143) <= input(13);
output(2, 144) <= input(73);
output(2, 145) <= input(17);
output(2, 146) <= input(18);
output(2, 147) <= input(19);
output(2, 148) <= input(20);
output(2, 149) <= input(21);
output(2, 150) <= input(22);
output(2, 151) <= input(23);
output(2, 152) <= input(24);
output(2, 153) <= input(25);
output(2, 154) <= input(26);
output(2, 155) <= input(27);
output(2, 156) <= input(28);
output(2, 157) <= input(29);
output(2, 158) <= input(30);
output(2, 159) <= input(31);
output(2, 160) <= input(74);
output(2, 161) <= input(37);
output(2, 162) <= input(16);
output(2, 163) <= input(0);
output(2, 164) <= input(1);
output(2, 165) <= input(2);
output(2, 166) <= input(3);
output(2, 167) <= input(4);
output(2, 168) <= input(5);
output(2, 169) <= input(6);
output(2, 170) <= input(7);
output(2, 171) <= input(8);
output(2, 172) <= input(9);
output(2, 173) <= input(10);
output(2, 174) <= input(11);
output(2, 175) <= input(12);
output(2, 176) <= input(75);
output(2, 177) <= input(73);
output(2, 178) <= input(17);
output(2, 179) <= input(18);
output(2, 180) <= input(19);
output(2, 181) <= input(20);
output(2, 182) <= input(21);
output(2, 183) <= input(22);
output(2, 184) <= input(23);
output(2, 185) <= input(24);
output(2, 186) <= input(25);
output(2, 187) <= input(26);
output(2, 188) <= input(27);
output(2, 189) <= input(28);
output(2, 190) <= input(29);
output(2, 191) <= input(30);
output(2, 192) <= input(76);
output(2, 193) <= input(75);
output(2, 194) <= input(73);
output(2, 195) <= input(17);
output(2, 196) <= input(18);
output(2, 197) <= input(19);
output(2, 198) <= input(20);
output(2, 199) <= input(21);
output(2, 200) <= input(22);
output(2, 201) <= input(23);
output(2, 202) <= input(24);
output(2, 203) <= input(25);
output(2, 204) <= input(26);
output(2, 205) <= input(27);
output(2, 206) <= input(28);
output(2, 207) <= input(29);
output(2, 208) <= input(77);
output(2, 209) <= input(78);
output(2, 210) <= input(74);
output(2, 211) <= input(37);
output(2, 212) <= input(16);
output(2, 213) <= input(0);
output(2, 214) <= input(1);
output(2, 215) <= input(2);
output(2, 216) <= input(3);
output(2, 217) <= input(4);
output(2, 218) <= input(5);
output(2, 219) <= input(6);
output(2, 220) <= input(7);
output(2, 221) <= input(8);
output(2, 222) <= input(9);
output(2, 223) <= input(10);
output(2, 224) <= input(79);
output(2, 225) <= input(76);
output(2, 226) <= input(75);
output(2, 227) <= input(73);
output(2, 228) <= input(17);
output(2, 229) <= input(18);
output(2, 230) <= input(19);
output(2, 231) <= input(20);
output(2, 232) <= input(21);
output(2, 233) <= input(22);
output(2, 234) <= input(23);
output(2, 235) <= input(24);
output(2, 236) <= input(25);
output(2, 237) <= input(26);
output(2, 238) <= input(27);
output(2, 239) <= input(28);
output(2, 240) <= input(80);
output(2, 241) <= input(77);
output(2, 242) <= input(78);
output(2, 243) <= input(74);
output(2, 244) <= input(37);
output(2, 245) <= input(16);
output(2, 246) <= input(0);
output(2, 247) <= input(1);
output(2, 248) <= input(2);
output(2, 249) <= input(3);
output(2, 250) <= input(4);
output(2, 251) <= input(5);
output(2, 252) <= input(6);
output(2, 253) <= input(7);
output(2, 254) <= input(8);
output(2, 255) <= input(9);
when "1010" =>
output(0, 0) <= input(0);
output(0, 1) <= input(1);
output(0, 2) <= input(2);
output(0, 3) <= input(3);
output(0, 4) <= input(4);
output(0, 5) <= input(5);
output(0, 6) <= input(6);
output(0, 7) <= input(7);
output(0, 8) <= input(8);
output(0, 9) <= input(9);
output(0, 10) <= input(10);
output(0, 11) <= input(11);
output(0, 12) <= input(12);
output(0, 13) <= input(13);
output(0, 14) <= input(14);
output(0, 15) <= input(15);
output(0, 16) <= input(16);
output(0, 17) <= input(17);
output(0, 18) <= input(18);
output(0, 19) <= input(19);
output(0, 20) <= input(20);
output(0, 21) <= input(21);
output(0, 22) <= input(22);
output(0, 23) <= input(23);
output(0, 24) <= input(24);
output(0, 25) <= input(25);
output(0, 26) <= input(26);
output(0, 27) <= input(27);
output(0, 28) <= input(28);
output(0, 29) <= input(29);
output(0, 30) <= input(30);
output(0, 31) <= input(31);
output(0, 32) <= input(32);
output(0, 33) <= input(0);
output(0, 34) <= input(1);
output(0, 35) <= input(2);
output(0, 36) <= input(3);
output(0, 37) <= input(4);
output(0, 38) <= input(5);
output(0, 39) <= input(6);
output(0, 40) <= input(7);
output(0, 41) <= input(8);
output(0, 42) <= input(9);
output(0, 43) <= input(10);
output(0, 44) <= input(11);
output(0, 45) <= input(12);
output(0, 46) <= input(13);
output(0, 47) <= input(14);
output(0, 48) <= input(33);
output(0, 49) <= input(16);
output(0, 50) <= input(17);
output(0, 51) <= input(18);
output(0, 52) <= input(19);
output(0, 53) <= input(20);
output(0, 54) <= input(21);
output(0, 55) <= input(22);
output(0, 56) <= input(23);
output(0, 57) <= input(24);
output(0, 58) <= input(25);
output(0, 59) <= input(26);
output(0, 60) <= input(27);
output(0, 61) <= input(28);
output(0, 62) <= input(29);
output(0, 63) <= input(30);
output(0, 64) <= input(34);
output(0, 65) <= input(32);
output(0, 66) <= input(0);
output(0, 67) <= input(1);
output(0, 68) <= input(2);
output(0, 69) <= input(3);
output(0, 70) <= input(4);
output(0, 71) <= input(5);
output(0, 72) <= input(6);
output(0, 73) <= input(7);
output(0, 74) <= input(8);
output(0, 75) <= input(9);
output(0, 76) <= input(10);
output(0, 77) <= input(11);
output(0, 78) <= input(12);
output(0, 79) <= input(13);
output(0, 80) <= input(35);
output(0, 81) <= input(33);
output(0, 82) <= input(16);
output(0, 83) <= input(17);
output(0, 84) <= input(18);
output(0, 85) <= input(19);
output(0, 86) <= input(20);
output(0, 87) <= input(21);
output(0, 88) <= input(22);
output(0, 89) <= input(23);
output(0, 90) <= input(24);
output(0, 91) <= input(25);
output(0, 92) <= input(26);
output(0, 93) <= input(27);
output(0, 94) <= input(28);
output(0, 95) <= input(29);
output(0, 96) <= input(36);
output(0, 97) <= input(34);
output(0, 98) <= input(32);
output(0, 99) <= input(0);
output(0, 100) <= input(1);
output(0, 101) <= input(2);
output(0, 102) <= input(3);
output(0, 103) <= input(4);
output(0, 104) <= input(5);
output(0, 105) <= input(6);
output(0, 106) <= input(7);
output(0, 107) <= input(8);
output(0, 108) <= input(9);
output(0, 109) <= input(10);
output(0, 110) <= input(11);
output(0, 111) <= input(12);
output(0, 112) <= input(37);
output(0, 113) <= input(35);
output(0, 114) <= input(33);
output(0, 115) <= input(16);
output(0, 116) <= input(17);
output(0, 117) <= input(18);
output(0, 118) <= input(19);
output(0, 119) <= input(20);
output(0, 120) <= input(21);
output(0, 121) <= input(22);
output(0, 122) <= input(23);
output(0, 123) <= input(24);
output(0, 124) <= input(25);
output(0, 125) <= input(26);
output(0, 126) <= input(27);
output(0, 127) <= input(28);
output(0, 128) <= input(38);
output(0, 129) <= input(37);
output(0, 130) <= input(35);
output(0, 131) <= input(33);
output(0, 132) <= input(16);
output(0, 133) <= input(17);
output(0, 134) <= input(18);
output(0, 135) <= input(19);
output(0, 136) <= input(20);
output(0, 137) <= input(21);
output(0, 138) <= input(22);
output(0, 139) <= input(23);
output(0, 140) <= input(24);
output(0, 141) <= input(25);
output(0, 142) <= input(26);
output(0, 143) <= input(27);
output(0, 144) <= input(39);
output(0, 145) <= input(40);
output(0, 146) <= input(36);
output(0, 147) <= input(34);
output(0, 148) <= input(32);
output(0, 149) <= input(0);
output(0, 150) <= input(1);
output(0, 151) <= input(2);
output(0, 152) <= input(3);
output(0, 153) <= input(4);
output(0, 154) <= input(5);
output(0, 155) <= input(6);
output(0, 156) <= input(7);
output(0, 157) <= input(8);
output(0, 158) <= input(9);
output(0, 159) <= input(10);
output(0, 160) <= input(41);
output(0, 161) <= input(38);
output(0, 162) <= input(37);
output(0, 163) <= input(35);
output(0, 164) <= input(33);
output(0, 165) <= input(16);
output(0, 166) <= input(17);
output(0, 167) <= input(18);
output(0, 168) <= input(19);
output(0, 169) <= input(20);
output(0, 170) <= input(21);
output(0, 171) <= input(22);
output(0, 172) <= input(23);
output(0, 173) <= input(24);
output(0, 174) <= input(25);
output(0, 175) <= input(26);
output(0, 176) <= input(42);
output(0, 177) <= input(39);
output(0, 178) <= input(40);
output(0, 179) <= input(36);
output(0, 180) <= input(34);
output(0, 181) <= input(32);
output(0, 182) <= input(0);
output(0, 183) <= input(1);
output(0, 184) <= input(2);
output(0, 185) <= input(3);
output(0, 186) <= input(4);
output(0, 187) <= input(5);
output(0, 188) <= input(6);
output(0, 189) <= input(7);
output(0, 190) <= input(8);
output(0, 191) <= input(9);
output(0, 192) <= input(43);
output(0, 193) <= input(41);
output(0, 194) <= input(38);
output(0, 195) <= input(37);
output(0, 196) <= input(35);
output(0, 197) <= input(33);
output(0, 198) <= input(16);
output(0, 199) <= input(17);
output(0, 200) <= input(18);
output(0, 201) <= input(19);
output(0, 202) <= input(20);
output(0, 203) <= input(21);
output(0, 204) <= input(22);
output(0, 205) <= input(23);
output(0, 206) <= input(24);
output(0, 207) <= input(25);
output(0, 208) <= input(44);
output(0, 209) <= input(42);
output(0, 210) <= input(39);
output(0, 211) <= input(40);
output(0, 212) <= input(36);
output(0, 213) <= input(34);
output(0, 214) <= input(32);
output(0, 215) <= input(0);
output(0, 216) <= input(1);
output(0, 217) <= input(2);
output(0, 218) <= input(3);
output(0, 219) <= input(4);
output(0, 220) <= input(5);
output(0, 221) <= input(6);
output(0, 222) <= input(7);
output(0, 223) <= input(8);
output(0, 224) <= input(45);
output(0, 225) <= input(43);
output(0, 226) <= input(41);
output(0, 227) <= input(38);
output(0, 228) <= input(37);
output(0, 229) <= input(35);
output(0, 230) <= input(33);
output(0, 231) <= input(16);
output(0, 232) <= input(17);
output(0, 233) <= input(18);
output(0, 234) <= input(19);
output(0, 235) <= input(20);
output(0, 236) <= input(21);
output(0, 237) <= input(22);
output(0, 238) <= input(23);
output(0, 239) <= input(24);
output(0, 240) <= input(46);
output(0, 241) <= input(44);
output(0, 242) <= input(42);
output(0, 243) <= input(39);
output(0, 244) <= input(40);
output(0, 245) <= input(36);
output(0, 246) <= input(34);
output(0, 247) <= input(32);
output(0, 248) <= input(0);
output(0, 249) <= input(1);
output(0, 250) <= input(2);
output(0, 251) <= input(3);
output(0, 252) <= input(4);
output(0, 253) <= input(5);
output(0, 254) <= input(6);
output(0, 255) <= input(7);
output(1, 0) <= input(18);
output(1, 1) <= input(19);
output(1, 2) <= input(20);
output(1, 3) <= input(21);
output(1, 4) <= input(22);
output(1, 5) <= input(23);
output(1, 6) <= input(24);
output(1, 7) <= input(25);
output(1, 8) <= input(26);
output(1, 9) <= input(27);
output(1, 10) <= input(28);
output(1, 11) <= input(29);
output(1, 12) <= input(30);
output(1, 13) <= input(31);
output(1, 14) <= input(47);
output(1, 15) <= input(48);
output(1, 16) <= input(1);
output(1, 17) <= input(2);
output(1, 18) <= input(3);
output(1, 19) <= input(4);
output(1, 20) <= input(5);
output(1, 21) <= input(6);
output(1, 22) <= input(7);
output(1, 23) <= input(8);
output(1, 24) <= input(9);
output(1, 25) <= input(10);
output(1, 26) <= input(11);
output(1, 27) <= input(12);
output(1, 28) <= input(13);
output(1, 29) <= input(14);
output(1, 30) <= input(15);
output(1, 31) <= input(49);
output(1, 32) <= input(17);
output(1, 33) <= input(18);
output(1, 34) <= input(19);
output(1, 35) <= input(20);
output(1, 36) <= input(21);
output(1, 37) <= input(22);
output(1, 38) <= input(23);
output(1, 39) <= input(24);
output(1, 40) <= input(25);
output(1, 41) <= input(26);
output(1, 42) <= input(27);
output(1, 43) <= input(28);
output(1, 44) <= input(29);
output(1, 45) <= input(30);
output(1, 46) <= input(31);
output(1, 47) <= input(47);
output(1, 48) <= input(0);
output(1, 49) <= input(1);
output(1, 50) <= input(2);
output(1, 51) <= input(3);
output(1, 52) <= input(4);
output(1, 53) <= input(5);
output(1, 54) <= input(6);
output(1, 55) <= input(7);
output(1, 56) <= input(8);
output(1, 57) <= input(9);
output(1, 58) <= input(10);
output(1, 59) <= input(11);
output(1, 60) <= input(12);
output(1, 61) <= input(13);
output(1, 62) <= input(14);
output(1, 63) <= input(15);
output(1, 64) <= input(16);
output(1, 65) <= input(17);
output(1, 66) <= input(18);
output(1, 67) <= input(19);
output(1, 68) <= input(20);
output(1, 69) <= input(21);
output(1, 70) <= input(22);
output(1, 71) <= input(23);
output(1, 72) <= input(24);
output(1, 73) <= input(25);
output(1, 74) <= input(26);
output(1, 75) <= input(27);
output(1, 76) <= input(28);
output(1, 77) <= input(29);
output(1, 78) <= input(30);
output(1, 79) <= input(31);
output(1, 80) <= input(32);
output(1, 81) <= input(0);
output(1, 82) <= input(1);
output(1, 83) <= input(2);
output(1, 84) <= input(3);
output(1, 85) <= input(4);
output(1, 86) <= input(5);
output(1, 87) <= input(6);
output(1, 88) <= input(7);
output(1, 89) <= input(8);
output(1, 90) <= input(9);
output(1, 91) <= input(10);
output(1, 92) <= input(11);
output(1, 93) <= input(12);
output(1, 94) <= input(13);
output(1, 95) <= input(14);
output(1, 96) <= input(33);
output(1, 97) <= input(16);
output(1, 98) <= input(17);
output(1, 99) <= input(18);
output(1, 100) <= input(19);
output(1, 101) <= input(20);
output(1, 102) <= input(21);
output(1, 103) <= input(22);
output(1, 104) <= input(23);
output(1, 105) <= input(24);
output(1, 106) <= input(25);
output(1, 107) <= input(26);
output(1, 108) <= input(27);
output(1, 109) <= input(28);
output(1, 110) <= input(29);
output(1, 111) <= input(30);
output(1, 112) <= input(34);
output(1, 113) <= input(32);
output(1, 114) <= input(0);
output(1, 115) <= input(1);
output(1, 116) <= input(2);
output(1, 117) <= input(3);
output(1, 118) <= input(4);
output(1, 119) <= input(5);
output(1, 120) <= input(6);
output(1, 121) <= input(7);
output(1, 122) <= input(8);
output(1, 123) <= input(9);
output(1, 124) <= input(10);
output(1, 125) <= input(11);
output(1, 126) <= input(12);
output(1, 127) <= input(13);
output(1, 128) <= input(35);
output(1, 129) <= input(33);
output(1, 130) <= input(16);
output(1, 131) <= input(17);
output(1, 132) <= input(18);
output(1, 133) <= input(19);
output(1, 134) <= input(20);
output(1, 135) <= input(21);
output(1, 136) <= input(22);
output(1, 137) <= input(23);
output(1, 138) <= input(24);
output(1, 139) <= input(25);
output(1, 140) <= input(26);
output(1, 141) <= input(27);
output(1, 142) <= input(28);
output(1, 143) <= input(29);
output(1, 144) <= input(36);
output(1, 145) <= input(34);
output(1, 146) <= input(32);
output(1, 147) <= input(0);
output(1, 148) <= input(1);
output(1, 149) <= input(2);
output(1, 150) <= input(3);
output(1, 151) <= input(4);
output(1, 152) <= input(5);
output(1, 153) <= input(6);
output(1, 154) <= input(7);
output(1, 155) <= input(8);
output(1, 156) <= input(9);
output(1, 157) <= input(10);
output(1, 158) <= input(11);
output(1, 159) <= input(12);
output(1, 160) <= input(37);
output(1, 161) <= input(35);
output(1, 162) <= input(33);
output(1, 163) <= input(16);
output(1, 164) <= input(17);
output(1, 165) <= input(18);
output(1, 166) <= input(19);
output(1, 167) <= input(20);
output(1, 168) <= input(21);
output(1, 169) <= input(22);
output(1, 170) <= input(23);
output(1, 171) <= input(24);
output(1, 172) <= input(25);
output(1, 173) <= input(26);
output(1, 174) <= input(27);
output(1, 175) <= input(28);
output(1, 176) <= input(40);
output(1, 177) <= input(36);
output(1, 178) <= input(34);
output(1, 179) <= input(32);
output(1, 180) <= input(0);
output(1, 181) <= input(1);
output(1, 182) <= input(2);
output(1, 183) <= input(3);
output(1, 184) <= input(4);
output(1, 185) <= input(5);
output(1, 186) <= input(6);
output(1, 187) <= input(7);
output(1, 188) <= input(8);
output(1, 189) <= input(9);
output(1, 190) <= input(10);
output(1, 191) <= input(11);
output(1, 192) <= input(38);
output(1, 193) <= input(37);
output(1, 194) <= input(35);
output(1, 195) <= input(33);
output(1, 196) <= input(16);
output(1, 197) <= input(17);
output(1, 198) <= input(18);
output(1, 199) <= input(19);
output(1, 200) <= input(20);
output(1, 201) <= input(21);
output(1, 202) <= input(22);
output(1, 203) <= input(23);
output(1, 204) <= input(24);
output(1, 205) <= input(25);
output(1, 206) <= input(26);
output(1, 207) <= input(27);
output(1, 208) <= input(39);
output(1, 209) <= input(40);
output(1, 210) <= input(36);
output(1, 211) <= input(34);
output(1, 212) <= input(32);
output(1, 213) <= input(0);
output(1, 214) <= input(1);
output(1, 215) <= input(2);
output(1, 216) <= input(3);
output(1, 217) <= input(4);
output(1, 218) <= input(5);
output(1, 219) <= input(6);
output(1, 220) <= input(7);
output(1, 221) <= input(8);
output(1, 222) <= input(9);
output(1, 223) <= input(10);
output(1, 224) <= input(41);
output(1, 225) <= input(38);
output(1, 226) <= input(37);
output(1, 227) <= input(35);
output(1, 228) <= input(33);
output(1, 229) <= input(16);
output(1, 230) <= input(17);
output(1, 231) <= input(18);
output(1, 232) <= input(19);
output(1, 233) <= input(20);
output(1, 234) <= input(21);
output(1, 235) <= input(22);
output(1, 236) <= input(23);
output(1, 237) <= input(24);
output(1, 238) <= input(25);
output(1, 239) <= input(26);
output(1, 240) <= input(42);
output(1, 241) <= input(39);
output(1, 242) <= input(40);
output(1, 243) <= input(36);
output(1, 244) <= input(34);
output(1, 245) <= input(32);
output(1, 246) <= input(0);
output(1, 247) <= input(1);
output(1, 248) <= input(2);
output(1, 249) <= input(3);
output(1, 250) <= input(4);
output(1, 251) <= input(5);
output(1, 252) <= input(6);
output(1, 253) <= input(7);
output(1, 254) <= input(8);
output(1, 255) <= input(9);
when "1011" =>
output(0, 0) <= input(0);
output(0, 1) <= input(1);
output(0, 2) <= input(2);
output(0, 3) <= input(3);
output(0, 4) <= input(4);
output(0, 5) <= input(5);
output(0, 6) <= input(6);
output(0, 7) <= input(7);
output(0, 8) <= input(8);
output(0, 9) <= input(9);
output(0, 10) <= input(10);
output(0, 11) <= input(11);
output(0, 12) <= input(12);
output(0, 13) <= input(13);
output(0, 14) <= input(14);
output(0, 15) <= input(15);
output(0, 16) <= input(16);
output(0, 17) <= input(17);
output(0, 18) <= input(18);
output(0, 19) <= input(19);
output(0, 20) <= input(20);
output(0, 21) <= input(21);
output(0, 22) <= input(22);
output(0, 23) <= input(23);
output(0, 24) <= input(24);
output(0, 25) <= input(25);
output(0, 26) <= input(26);
output(0, 27) <= input(27);
output(0, 28) <= input(28);
output(0, 29) <= input(29);
output(0, 30) <= input(30);
output(0, 31) <= input(31);
output(0, 32) <= input(32);
output(0, 33) <= input(0);
output(0, 34) <= input(1);
output(0, 35) <= input(2);
output(0, 36) <= input(3);
output(0, 37) <= input(4);
output(0, 38) <= input(5);
output(0, 39) <= input(6);
output(0, 40) <= input(7);
output(0, 41) <= input(8);
output(0, 42) <= input(9);
output(0, 43) <= input(10);
output(0, 44) <= input(11);
output(0, 45) <= input(12);
output(0, 46) <= input(13);
output(0, 47) <= input(14);
output(0, 48) <= input(33);
output(0, 49) <= input(16);
output(0, 50) <= input(17);
output(0, 51) <= input(18);
output(0, 52) <= input(19);
output(0, 53) <= input(20);
output(0, 54) <= input(21);
output(0, 55) <= input(22);
output(0, 56) <= input(23);
output(0, 57) <= input(24);
output(0, 58) <= input(25);
output(0, 59) <= input(26);
output(0, 60) <= input(27);
output(0, 61) <= input(28);
output(0, 62) <= input(29);
output(0, 63) <= input(30);
output(0, 64) <= input(34);
output(0, 65) <= input(32);
output(0, 66) <= input(0);
output(0, 67) <= input(1);
output(0, 68) <= input(2);
output(0, 69) <= input(3);
output(0, 70) <= input(4);
output(0, 71) <= input(5);
output(0, 72) <= input(6);
output(0, 73) <= input(7);
output(0, 74) <= input(8);
output(0, 75) <= input(9);
output(0, 76) <= input(10);
output(0, 77) <= input(11);
output(0, 78) <= input(12);
output(0, 79) <= input(13);
output(0, 80) <= input(35);
output(0, 81) <= input(33);
output(0, 82) <= input(16);
output(0, 83) <= input(17);
output(0, 84) <= input(18);
output(0, 85) <= input(19);
output(0, 86) <= input(20);
output(0, 87) <= input(21);
output(0, 88) <= input(22);
output(0, 89) <= input(23);
output(0, 90) <= input(24);
output(0, 91) <= input(25);
output(0, 92) <= input(26);
output(0, 93) <= input(27);
output(0, 94) <= input(28);
output(0, 95) <= input(29);
output(0, 96) <= input(36);
output(0, 97) <= input(34);
output(0, 98) <= input(32);
output(0, 99) <= input(0);
output(0, 100) <= input(1);
output(0, 101) <= input(2);
output(0, 102) <= input(3);
output(0, 103) <= input(4);
output(0, 104) <= input(5);
output(0, 105) <= input(6);
output(0, 106) <= input(7);
output(0, 107) <= input(8);
output(0, 108) <= input(9);
output(0, 109) <= input(10);
output(0, 110) <= input(11);
output(0, 111) <= input(12);
output(0, 112) <= input(36);
output(0, 113) <= input(34);
output(0, 114) <= input(32);
output(0, 115) <= input(0);
output(0, 116) <= input(1);
output(0, 117) <= input(2);
output(0, 118) <= input(3);
output(0, 119) <= input(4);
output(0, 120) <= input(5);
output(0, 121) <= input(6);
output(0, 122) <= input(7);
output(0, 123) <= input(8);
output(0, 124) <= input(9);
output(0, 125) <= input(10);
output(0, 126) <= input(11);
output(0, 127) <= input(12);
output(0, 128) <= input(37);
output(0, 129) <= input(35);
output(0, 130) <= input(33);
output(0, 131) <= input(16);
output(0, 132) <= input(17);
output(0, 133) <= input(18);
output(0, 134) <= input(19);
output(0, 135) <= input(20);
output(0, 136) <= input(21);
output(0, 137) <= input(22);
output(0, 138) <= input(23);
output(0, 139) <= input(24);
output(0, 140) <= input(25);
output(0, 141) <= input(26);
output(0, 142) <= input(27);
output(0, 143) <= input(28);
output(0, 144) <= input(38);
output(0, 145) <= input(36);
output(0, 146) <= input(34);
output(0, 147) <= input(32);
output(0, 148) <= input(0);
output(0, 149) <= input(1);
output(0, 150) <= input(2);
output(0, 151) <= input(3);
output(0, 152) <= input(4);
output(0, 153) <= input(5);
output(0, 154) <= input(6);
output(0, 155) <= input(7);
output(0, 156) <= input(8);
output(0, 157) <= input(9);
output(0, 158) <= input(10);
output(0, 159) <= input(11);
output(0, 160) <= input(39);
output(0, 161) <= input(37);
output(0, 162) <= input(35);
output(0, 163) <= input(33);
output(0, 164) <= input(16);
output(0, 165) <= input(17);
output(0, 166) <= input(18);
output(0, 167) <= input(19);
output(0, 168) <= input(20);
output(0, 169) <= input(21);
output(0, 170) <= input(22);
output(0, 171) <= input(23);
output(0, 172) <= input(24);
output(0, 173) <= input(25);
output(0, 174) <= input(26);
output(0, 175) <= input(27);
output(0, 176) <= input(40);
output(0, 177) <= input(38);
output(0, 178) <= input(36);
output(0, 179) <= input(34);
output(0, 180) <= input(32);
output(0, 181) <= input(0);
output(0, 182) <= input(1);
output(0, 183) <= input(2);
output(0, 184) <= input(3);
output(0, 185) <= input(4);
output(0, 186) <= input(5);
output(0, 187) <= input(6);
output(0, 188) <= input(7);
output(0, 189) <= input(8);
output(0, 190) <= input(9);
output(0, 191) <= input(10);
output(0, 192) <= input(41);
output(0, 193) <= input(39);
output(0, 194) <= input(37);
output(0, 195) <= input(35);
output(0, 196) <= input(33);
output(0, 197) <= input(16);
output(0, 198) <= input(17);
output(0, 199) <= input(18);
output(0, 200) <= input(19);
output(0, 201) <= input(20);
output(0, 202) <= input(21);
output(0, 203) <= input(22);
output(0, 204) <= input(23);
output(0, 205) <= input(24);
output(0, 206) <= input(25);
output(0, 207) <= input(26);
output(0, 208) <= input(42);
output(0, 209) <= input(40);
output(0, 210) <= input(38);
output(0, 211) <= input(36);
output(0, 212) <= input(34);
output(0, 213) <= input(32);
output(0, 214) <= input(0);
output(0, 215) <= input(1);
output(0, 216) <= input(2);
output(0, 217) <= input(3);
output(0, 218) <= input(4);
output(0, 219) <= input(5);
output(0, 220) <= input(6);
output(0, 221) <= input(7);
output(0, 222) <= input(8);
output(0, 223) <= input(9);
output(0, 224) <= input(43);
output(0, 225) <= input(41);
output(0, 226) <= input(39);
output(0, 227) <= input(37);
output(0, 228) <= input(35);
output(0, 229) <= input(33);
output(0, 230) <= input(16);
output(0, 231) <= input(17);
output(0, 232) <= input(18);
output(0, 233) <= input(19);
output(0, 234) <= input(20);
output(0, 235) <= input(21);
output(0, 236) <= input(22);
output(0, 237) <= input(23);
output(0, 238) <= input(24);
output(0, 239) <= input(25);
output(0, 240) <= input(43);
output(0, 241) <= input(41);
output(0, 242) <= input(39);
output(0, 243) <= input(37);
output(0, 244) <= input(35);
output(0, 245) <= input(33);
output(0, 246) <= input(16);
output(0, 247) <= input(17);
output(0, 248) <= input(18);
output(0, 249) <= input(19);
output(0, 250) <= input(20);
output(0, 251) <= input(21);
output(0, 252) <= input(22);
output(0, 253) <= input(23);
output(0, 254) <= input(24);
output(0, 255) <= input(25);
output(1, 0) <= input(1);
output(1, 1) <= input(2);
output(1, 2) <= input(3);
output(1, 3) <= input(4);
output(1, 4) <= input(5);
output(1, 5) <= input(6);
output(1, 6) <= input(7);
output(1, 7) <= input(8);
output(1, 8) <= input(9);
output(1, 9) <= input(10);
output(1, 10) <= input(11);
output(1, 11) <= input(12);
output(1, 12) <= input(13);
output(1, 13) <= input(14);
output(1, 14) <= input(15);
output(1, 15) <= input(44);
output(1, 16) <= input(17);
output(1, 17) <= input(18);
output(1, 18) <= input(19);
output(1, 19) <= input(20);
output(1, 20) <= input(21);
output(1, 21) <= input(22);
output(1, 22) <= input(23);
output(1, 23) <= input(24);
output(1, 24) <= input(25);
output(1, 25) <= input(26);
output(1, 26) <= input(27);
output(1, 27) <= input(28);
output(1, 28) <= input(29);
output(1, 29) <= input(30);
output(1, 30) <= input(31);
output(1, 31) <= input(45);
output(1, 32) <= input(0);
output(1, 33) <= input(1);
output(1, 34) <= input(2);
output(1, 35) <= input(3);
output(1, 36) <= input(4);
output(1, 37) <= input(5);
output(1, 38) <= input(6);
output(1, 39) <= input(7);
output(1, 40) <= input(8);
output(1, 41) <= input(9);
output(1, 42) <= input(10);
output(1, 43) <= input(11);
output(1, 44) <= input(12);
output(1, 45) <= input(13);
output(1, 46) <= input(14);
output(1, 47) <= input(15);
output(1, 48) <= input(0);
output(1, 49) <= input(1);
output(1, 50) <= input(2);
output(1, 51) <= input(3);
output(1, 52) <= input(4);
output(1, 53) <= input(5);
output(1, 54) <= input(6);
output(1, 55) <= input(7);
output(1, 56) <= input(8);
output(1, 57) <= input(9);
output(1, 58) <= input(10);
output(1, 59) <= input(11);
output(1, 60) <= input(12);
output(1, 61) <= input(13);
output(1, 62) <= input(14);
output(1, 63) <= input(15);
output(1, 64) <= input(16);
output(1, 65) <= input(17);
output(1, 66) <= input(18);
output(1, 67) <= input(19);
output(1, 68) <= input(20);
output(1, 69) <= input(21);
output(1, 70) <= input(22);
output(1, 71) <= input(23);
output(1, 72) <= input(24);
output(1, 73) <= input(25);
output(1, 74) <= input(26);
output(1, 75) <= input(27);
output(1, 76) <= input(28);
output(1, 77) <= input(29);
output(1, 78) <= input(30);
output(1, 79) <= input(31);
output(1, 80) <= input(32);
output(1, 81) <= input(0);
output(1, 82) <= input(1);
output(1, 83) <= input(2);
output(1, 84) <= input(3);
output(1, 85) <= input(4);
output(1, 86) <= input(5);
output(1, 87) <= input(6);
output(1, 88) <= input(7);
output(1, 89) <= input(8);
output(1, 90) <= input(9);
output(1, 91) <= input(10);
output(1, 92) <= input(11);
output(1, 93) <= input(12);
output(1, 94) <= input(13);
output(1, 95) <= input(14);
output(1, 96) <= input(33);
output(1, 97) <= input(16);
output(1, 98) <= input(17);
output(1, 99) <= input(18);
output(1, 100) <= input(19);
output(1, 101) <= input(20);
output(1, 102) <= input(21);
output(1, 103) <= input(22);
output(1, 104) <= input(23);
output(1, 105) <= input(24);
output(1, 106) <= input(25);
output(1, 107) <= input(26);
output(1, 108) <= input(27);
output(1, 109) <= input(28);
output(1, 110) <= input(29);
output(1, 111) <= input(30);
output(1, 112) <= input(33);
output(1, 113) <= input(16);
output(1, 114) <= input(17);
output(1, 115) <= input(18);
output(1, 116) <= input(19);
output(1, 117) <= input(20);
output(1, 118) <= input(21);
output(1, 119) <= input(22);
output(1, 120) <= input(23);
output(1, 121) <= input(24);
output(1, 122) <= input(25);
output(1, 123) <= input(26);
output(1, 124) <= input(27);
output(1, 125) <= input(28);
output(1, 126) <= input(29);
output(1, 127) <= input(30);
output(1, 128) <= input(34);
output(1, 129) <= input(32);
output(1, 130) <= input(0);
output(1, 131) <= input(1);
output(1, 132) <= input(2);
output(1, 133) <= input(3);
output(1, 134) <= input(4);
output(1, 135) <= input(5);
output(1, 136) <= input(6);
output(1, 137) <= input(7);
output(1, 138) <= input(8);
output(1, 139) <= input(9);
output(1, 140) <= input(10);
output(1, 141) <= input(11);
output(1, 142) <= input(12);
output(1, 143) <= input(13);
output(1, 144) <= input(35);
output(1, 145) <= input(33);
output(1, 146) <= input(16);
output(1, 147) <= input(17);
output(1, 148) <= input(18);
output(1, 149) <= input(19);
output(1, 150) <= input(20);
output(1, 151) <= input(21);
output(1, 152) <= input(22);
output(1, 153) <= input(23);
output(1, 154) <= input(24);
output(1, 155) <= input(25);
output(1, 156) <= input(26);
output(1, 157) <= input(27);
output(1, 158) <= input(28);
output(1, 159) <= input(29);
output(1, 160) <= input(36);
output(1, 161) <= input(34);
output(1, 162) <= input(32);
output(1, 163) <= input(0);
output(1, 164) <= input(1);
output(1, 165) <= input(2);
output(1, 166) <= input(3);
output(1, 167) <= input(4);
output(1, 168) <= input(5);
output(1, 169) <= input(6);
output(1, 170) <= input(7);
output(1, 171) <= input(8);
output(1, 172) <= input(9);
output(1, 173) <= input(10);
output(1, 174) <= input(11);
output(1, 175) <= input(12);
output(1, 176) <= input(36);
output(1, 177) <= input(34);
output(1, 178) <= input(32);
output(1, 179) <= input(0);
output(1, 180) <= input(1);
output(1, 181) <= input(2);
output(1, 182) <= input(3);
output(1, 183) <= input(4);
output(1, 184) <= input(5);
output(1, 185) <= input(6);
output(1, 186) <= input(7);
output(1, 187) <= input(8);
output(1, 188) <= input(9);
output(1, 189) <= input(10);
output(1, 190) <= input(11);
output(1, 191) <= input(12);
output(1, 192) <= input(37);
output(1, 193) <= input(35);
output(1, 194) <= input(33);
output(1, 195) <= input(16);
output(1, 196) <= input(17);
output(1, 197) <= input(18);
output(1, 198) <= input(19);
output(1, 199) <= input(20);
output(1, 200) <= input(21);
output(1, 201) <= input(22);
output(1, 202) <= input(23);
output(1, 203) <= input(24);
output(1, 204) <= input(25);
output(1, 205) <= input(26);
output(1, 206) <= input(27);
output(1, 207) <= input(28);
output(1, 208) <= input(38);
output(1, 209) <= input(36);
output(1, 210) <= input(34);
output(1, 211) <= input(32);
output(1, 212) <= input(0);
output(1, 213) <= input(1);
output(1, 214) <= input(2);
output(1, 215) <= input(3);
output(1, 216) <= input(4);
output(1, 217) <= input(5);
output(1, 218) <= input(6);
output(1, 219) <= input(7);
output(1, 220) <= input(8);
output(1, 221) <= input(9);
output(1, 222) <= input(10);
output(1, 223) <= input(11);
output(1, 224) <= input(39);
output(1, 225) <= input(37);
output(1, 226) <= input(35);
output(1, 227) <= input(33);
output(1, 228) <= input(16);
output(1, 229) <= input(17);
output(1, 230) <= input(18);
output(1, 231) <= input(19);
output(1, 232) <= input(20);
output(1, 233) <= input(21);
output(1, 234) <= input(22);
output(1, 235) <= input(23);
output(1, 236) <= input(24);
output(1, 237) <= input(25);
output(1, 238) <= input(26);
output(1, 239) <= input(27);
output(1, 240) <= input(39);
output(1, 241) <= input(37);
output(1, 242) <= input(35);
output(1, 243) <= input(33);
output(1, 244) <= input(16);
output(1, 245) <= input(17);
output(1, 246) <= input(18);
output(1, 247) <= input(19);
output(1, 248) <= input(20);
output(1, 249) <= input(21);
output(1, 250) <= input(22);
output(1, 251) <= input(23);
output(1, 252) <= input(24);
output(1, 253) <= input(25);
output(1, 254) <= input(26);
output(1, 255) <= input(27);
output(2, 0) <= input(2);
output(2, 1) <= input(3);
output(2, 2) <= input(4);
output(2, 3) <= input(5);
output(2, 4) <= input(6);
output(2, 5) <= input(7);
output(2, 6) <= input(8);
output(2, 7) <= input(9);
output(2, 8) <= input(10);
output(2, 9) <= input(11);
output(2, 10) <= input(12);
output(2, 11) <= input(13);
output(2, 12) <= input(14);
output(2, 13) <= input(15);
output(2, 14) <= input(44);
output(2, 15) <= input(46);
output(2, 16) <= input(18);
output(2, 17) <= input(19);
output(2, 18) <= input(20);
output(2, 19) <= input(21);
output(2, 20) <= input(22);
output(2, 21) <= input(23);
output(2, 22) <= input(24);
output(2, 23) <= input(25);
output(2, 24) <= input(26);
output(2, 25) <= input(27);
output(2, 26) <= input(28);
output(2, 27) <= input(29);
output(2, 28) <= input(30);
output(2, 29) <= input(31);
output(2, 30) <= input(45);
output(2, 31) <= input(47);
output(2, 32) <= input(18);
output(2, 33) <= input(19);
output(2, 34) <= input(20);
output(2, 35) <= input(21);
output(2, 36) <= input(22);
output(2, 37) <= input(23);
output(2, 38) <= input(24);
output(2, 39) <= input(25);
output(2, 40) <= input(26);
output(2, 41) <= input(27);
output(2, 42) <= input(28);
output(2, 43) <= input(29);
output(2, 44) <= input(30);
output(2, 45) <= input(31);
output(2, 46) <= input(45);
output(2, 47) <= input(47);
output(2, 48) <= input(1);
output(2, 49) <= input(2);
output(2, 50) <= input(3);
output(2, 51) <= input(4);
output(2, 52) <= input(5);
output(2, 53) <= input(6);
output(2, 54) <= input(7);
output(2, 55) <= input(8);
output(2, 56) <= input(9);
output(2, 57) <= input(10);
output(2, 58) <= input(11);
output(2, 59) <= input(12);
output(2, 60) <= input(13);
output(2, 61) <= input(14);
output(2, 62) <= input(15);
output(2, 63) <= input(44);
output(2, 64) <= input(17);
output(2, 65) <= input(18);
output(2, 66) <= input(19);
output(2, 67) <= input(20);
output(2, 68) <= input(21);
output(2, 69) <= input(22);
output(2, 70) <= input(23);
output(2, 71) <= input(24);
output(2, 72) <= input(25);
output(2, 73) <= input(26);
output(2, 74) <= input(27);
output(2, 75) <= input(28);
output(2, 76) <= input(29);
output(2, 77) <= input(30);
output(2, 78) <= input(31);
output(2, 79) <= input(45);
output(2, 80) <= input(17);
output(2, 81) <= input(18);
output(2, 82) <= input(19);
output(2, 83) <= input(20);
output(2, 84) <= input(21);
output(2, 85) <= input(22);
output(2, 86) <= input(23);
output(2, 87) <= input(24);
output(2, 88) <= input(25);
output(2, 89) <= input(26);
output(2, 90) <= input(27);
output(2, 91) <= input(28);
output(2, 92) <= input(29);
output(2, 93) <= input(30);
output(2, 94) <= input(31);
output(2, 95) <= input(45);
output(2, 96) <= input(0);
output(2, 97) <= input(1);
output(2, 98) <= input(2);
output(2, 99) <= input(3);
output(2, 100) <= input(4);
output(2, 101) <= input(5);
output(2, 102) <= input(6);
output(2, 103) <= input(7);
output(2, 104) <= input(8);
output(2, 105) <= input(9);
output(2, 106) <= input(10);
output(2, 107) <= input(11);
output(2, 108) <= input(12);
output(2, 109) <= input(13);
output(2, 110) <= input(14);
output(2, 111) <= input(15);
output(2, 112) <= input(0);
output(2, 113) <= input(1);
output(2, 114) <= input(2);
output(2, 115) <= input(3);
output(2, 116) <= input(4);
output(2, 117) <= input(5);
output(2, 118) <= input(6);
output(2, 119) <= input(7);
output(2, 120) <= input(8);
output(2, 121) <= input(9);
output(2, 122) <= input(10);
output(2, 123) <= input(11);
output(2, 124) <= input(12);
output(2, 125) <= input(13);
output(2, 126) <= input(14);
output(2, 127) <= input(15);
output(2, 128) <= input(16);
output(2, 129) <= input(17);
output(2, 130) <= input(18);
output(2, 131) <= input(19);
output(2, 132) <= input(20);
output(2, 133) <= input(21);
output(2, 134) <= input(22);
output(2, 135) <= input(23);
output(2, 136) <= input(24);
output(2, 137) <= input(25);
output(2, 138) <= input(26);
output(2, 139) <= input(27);
output(2, 140) <= input(28);
output(2, 141) <= input(29);
output(2, 142) <= input(30);
output(2, 143) <= input(31);
output(2, 144) <= input(32);
output(2, 145) <= input(0);
output(2, 146) <= input(1);
output(2, 147) <= input(2);
output(2, 148) <= input(3);
output(2, 149) <= input(4);
output(2, 150) <= input(5);
output(2, 151) <= input(6);
output(2, 152) <= input(7);
output(2, 153) <= input(8);
output(2, 154) <= input(9);
output(2, 155) <= input(10);
output(2, 156) <= input(11);
output(2, 157) <= input(12);
output(2, 158) <= input(13);
output(2, 159) <= input(14);
output(2, 160) <= input(32);
output(2, 161) <= input(0);
output(2, 162) <= input(1);
output(2, 163) <= input(2);
output(2, 164) <= input(3);
output(2, 165) <= input(4);
output(2, 166) <= input(5);
output(2, 167) <= input(6);
output(2, 168) <= input(7);
output(2, 169) <= input(8);
output(2, 170) <= input(9);
output(2, 171) <= input(10);
output(2, 172) <= input(11);
output(2, 173) <= input(12);
output(2, 174) <= input(13);
output(2, 175) <= input(14);
output(2, 176) <= input(33);
output(2, 177) <= input(16);
output(2, 178) <= input(17);
output(2, 179) <= input(18);
output(2, 180) <= input(19);
output(2, 181) <= input(20);
output(2, 182) <= input(21);
output(2, 183) <= input(22);
output(2, 184) <= input(23);
output(2, 185) <= input(24);
output(2, 186) <= input(25);
output(2, 187) <= input(26);
output(2, 188) <= input(27);
output(2, 189) <= input(28);
output(2, 190) <= input(29);
output(2, 191) <= input(30);
output(2, 192) <= input(34);
output(2, 193) <= input(32);
output(2, 194) <= input(0);
output(2, 195) <= input(1);
output(2, 196) <= input(2);
output(2, 197) <= input(3);
output(2, 198) <= input(4);
output(2, 199) <= input(5);
output(2, 200) <= input(6);
output(2, 201) <= input(7);
output(2, 202) <= input(8);
output(2, 203) <= input(9);
output(2, 204) <= input(10);
output(2, 205) <= input(11);
output(2, 206) <= input(12);
output(2, 207) <= input(13);
output(2, 208) <= input(34);
output(2, 209) <= input(32);
output(2, 210) <= input(0);
output(2, 211) <= input(1);
output(2, 212) <= input(2);
output(2, 213) <= input(3);
output(2, 214) <= input(4);
output(2, 215) <= input(5);
output(2, 216) <= input(6);
output(2, 217) <= input(7);
output(2, 218) <= input(8);
output(2, 219) <= input(9);
output(2, 220) <= input(10);
output(2, 221) <= input(11);
output(2, 222) <= input(12);
output(2, 223) <= input(13);
output(2, 224) <= input(35);
output(2, 225) <= input(33);
output(2, 226) <= input(16);
output(2, 227) <= input(17);
output(2, 228) <= input(18);
output(2, 229) <= input(19);
output(2, 230) <= input(20);
output(2, 231) <= input(21);
output(2, 232) <= input(22);
output(2, 233) <= input(23);
output(2, 234) <= input(24);
output(2, 235) <= input(25);
output(2, 236) <= input(26);
output(2, 237) <= input(27);
output(2, 238) <= input(28);
output(2, 239) <= input(29);
output(2, 240) <= input(35);
output(2, 241) <= input(33);
output(2, 242) <= input(16);
output(2, 243) <= input(17);
output(2, 244) <= input(18);
output(2, 245) <= input(19);
output(2, 246) <= input(20);
output(2, 247) <= input(21);
output(2, 248) <= input(22);
output(2, 249) <= input(23);
output(2, 250) <= input(24);
output(2, 251) <= input(25);
output(2, 252) <= input(26);
output(2, 253) <= input(27);
output(2, 254) <= input(28);
output(2, 255) <= input(29);
when "1100" =>
output(0, 0) <= input(0);
output(0, 1) <= input(1);
output(0, 2) <= input(2);
output(0, 3) <= input(3);
output(0, 4) <= input(4);
output(0, 5) <= input(5);
output(0, 6) <= input(6);
output(0, 7) <= input(7);
output(0, 8) <= input(8);
output(0, 9) <= input(9);
output(0, 10) <= input(10);
output(0, 11) <= input(11);
output(0, 12) <= input(12);
output(0, 13) <= input(13);
output(0, 14) <= input(14);
output(0, 15) <= input(15);
output(0, 16) <= input(0);
output(0, 17) <= input(1);
output(0, 18) <= input(2);
output(0, 19) <= input(3);
output(0, 20) <= input(4);
output(0, 21) <= input(5);
output(0, 22) <= input(6);
output(0, 23) <= input(7);
output(0, 24) <= input(8);
output(0, 25) <= input(9);
output(0, 26) <= input(10);
output(0, 27) <= input(11);
output(0, 28) <= input(12);
output(0, 29) <= input(13);
output(0, 30) <= input(14);
output(0, 31) <= input(15);
output(0, 32) <= input(16);
output(0, 33) <= input(17);
output(0, 34) <= input(18);
output(0, 35) <= input(19);
output(0, 36) <= input(20);
output(0, 37) <= input(21);
output(0, 38) <= input(22);
output(0, 39) <= input(23);
output(0, 40) <= input(24);
output(0, 41) <= input(25);
output(0, 42) <= input(26);
output(0, 43) <= input(27);
output(0, 44) <= input(28);
output(0, 45) <= input(29);
output(0, 46) <= input(30);
output(0, 47) <= input(31);
output(0, 48) <= input(16);
output(0, 49) <= input(17);
output(0, 50) <= input(18);
output(0, 51) <= input(19);
output(0, 52) <= input(20);
output(0, 53) <= input(21);
output(0, 54) <= input(22);
output(0, 55) <= input(23);
output(0, 56) <= input(24);
output(0, 57) <= input(25);
output(0, 58) <= input(26);
output(0, 59) <= input(27);
output(0, 60) <= input(28);
output(0, 61) <= input(29);
output(0, 62) <= input(30);
output(0, 63) <= input(31);
output(0, 64) <= input(32);
output(0, 65) <= input(0);
output(0, 66) <= input(1);
output(0, 67) <= input(2);
output(0, 68) <= input(3);
output(0, 69) <= input(4);
output(0, 70) <= input(5);
output(0, 71) <= input(6);
output(0, 72) <= input(7);
output(0, 73) <= input(8);
output(0, 74) <= input(9);
output(0, 75) <= input(10);
output(0, 76) <= input(11);
output(0, 77) <= input(12);
output(0, 78) <= input(13);
output(0, 79) <= input(14);
output(0, 80) <= input(32);
output(0, 81) <= input(0);
output(0, 82) <= input(1);
output(0, 83) <= input(2);
output(0, 84) <= input(3);
output(0, 85) <= input(4);
output(0, 86) <= input(5);
output(0, 87) <= input(6);
output(0, 88) <= input(7);
output(0, 89) <= input(8);
output(0, 90) <= input(9);
output(0, 91) <= input(10);
output(0, 92) <= input(11);
output(0, 93) <= input(12);
output(0, 94) <= input(13);
output(0, 95) <= input(14);
output(0, 96) <= input(33);
output(0, 97) <= input(16);
output(0, 98) <= input(17);
output(0, 99) <= input(18);
output(0, 100) <= input(19);
output(0, 101) <= input(20);
output(0, 102) <= input(21);
output(0, 103) <= input(22);
output(0, 104) <= input(23);
output(0, 105) <= input(24);
output(0, 106) <= input(25);
output(0, 107) <= input(26);
output(0, 108) <= input(27);
output(0, 109) <= input(28);
output(0, 110) <= input(29);
output(0, 111) <= input(30);
output(0, 112) <= input(33);
output(0, 113) <= input(16);
output(0, 114) <= input(17);
output(0, 115) <= input(18);
output(0, 116) <= input(19);
output(0, 117) <= input(20);
output(0, 118) <= input(21);
output(0, 119) <= input(22);
output(0, 120) <= input(23);
output(0, 121) <= input(24);
output(0, 122) <= input(25);
output(0, 123) <= input(26);
output(0, 124) <= input(27);
output(0, 125) <= input(28);
output(0, 126) <= input(29);
output(0, 127) <= input(30);
output(0, 128) <= input(34);
output(0, 129) <= input(32);
output(0, 130) <= input(0);
output(0, 131) <= input(1);
output(0, 132) <= input(2);
output(0, 133) <= input(3);
output(0, 134) <= input(4);
output(0, 135) <= input(5);
output(0, 136) <= input(6);
output(0, 137) <= input(7);
output(0, 138) <= input(8);
output(0, 139) <= input(9);
output(0, 140) <= input(10);
output(0, 141) <= input(11);
output(0, 142) <= input(12);
output(0, 143) <= input(13);
output(0, 144) <= input(34);
output(0, 145) <= input(32);
output(0, 146) <= input(0);
output(0, 147) <= input(1);
output(0, 148) <= input(2);
output(0, 149) <= input(3);
output(0, 150) <= input(4);
output(0, 151) <= input(5);
output(0, 152) <= input(6);
output(0, 153) <= input(7);
output(0, 154) <= input(8);
output(0, 155) <= input(9);
output(0, 156) <= input(10);
output(0, 157) <= input(11);
output(0, 158) <= input(12);
output(0, 159) <= input(13);
output(0, 160) <= input(35);
output(0, 161) <= input(33);
output(0, 162) <= input(16);
output(0, 163) <= input(17);
output(0, 164) <= input(18);
output(0, 165) <= input(19);
output(0, 166) <= input(20);
output(0, 167) <= input(21);
output(0, 168) <= input(22);
output(0, 169) <= input(23);
output(0, 170) <= input(24);
output(0, 171) <= input(25);
output(0, 172) <= input(26);
output(0, 173) <= input(27);
output(0, 174) <= input(28);
output(0, 175) <= input(29);
output(0, 176) <= input(35);
output(0, 177) <= input(33);
output(0, 178) <= input(16);
output(0, 179) <= input(17);
output(0, 180) <= input(18);
output(0, 181) <= input(19);
output(0, 182) <= input(20);
output(0, 183) <= input(21);
output(0, 184) <= input(22);
output(0, 185) <= input(23);
output(0, 186) <= input(24);
output(0, 187) <= input(25);
output(0, 188) <= input(26);
output(0, 189) <= input(27);
output(0, 190) <= input(28);
output(0, 191) <= input(29);
output(0, 192) <= input(36);
output(0, 193) <= input(34);
output(0, 194) <= input(32);
output(0, 195) <= input(0);
output(0, 196) <= input(1);
output(0, 197) <= input(2);
output(0, 198) <= input(3);
output(0, 199) <= input(4);
output(0, 200) <= input(5);
output(0, 201) <= input(6);
output(0, 202) <= input(7);
output(0, 203) <= input(8);
output(0, 204) <= input(9);
output(0, 205) <= input(10);
output(0, 206) <= input(11);
output(0, 207) <= input(12);
output(0, 208) <= input(36);
output(0, 209) <= input(34);
output(0, 210) <= input(32);
output(0, 211) <= input(0);
output(0, 212) <= input(1);
output(0, 213) <= input(2);
output(0, 214) <= input(3);
output(0, 215) <= input(4);
output(0, 216) <= input(5);
output(0, 217) <= input(6);
output(0, 218) <= input(7);
output(0, 219) <= input(8);
output(0, 220) <= input(9);
output(0, 221) <= input(10);
output(0, 222) <= input(11);
output(0, 223) <= input(12);
output(0, 224) <= input(37);
output(0, 225) <= input(35);
output(0, 226) <= input(33);
output(0, 227) <= input(16);
output(0, 228) <= input(17);
output(0, 229) <= input(18);
output(0, 230) <= input(19);
output(0, 231) <= input(20);
output(0, 232) <= input(21);
output(0, 233) <= input(22);
output(0, 234) <= input(23);
output(0, 235) <= input(24);
output(0, 236) <= input(25);
output(0, 237) <= input(26);
output(0, 238) <= input(27);
output(0, 239) <= input(28);
output(0, 240) <= input(37);
output(0, 241) <= input(35);
output(0, 242) <= input(33);
output(0, 243) <= input(16);
output(0, 244) <= input(17);
output(0, 245) <= input(18);
output(0, 246) <= input(19);
output(0, 247) <= input(20);
output(0, 248) <= input(21);
output(0, 249) <= input(22);
output(0, 250) <= input(23);
output(0, 251) <= input(24);
output(0, 252) <= input(25);
output(0, 253) <= input(26);
output(0, 254) <= input(27);
output(0, 255) <= input(28);
output(1, 0) <= input(1);
output(1, 1) <= input(2);
output(1, 2) <= input(3);
output(1, 3) <= input(4);
output(1, 4) <= input(5);
output(1, 5) <= input(6);
output(1, 6) <= input(7);
output(1, 7) <= input(8);
output(1, 8) <= input(9);
output(1, 9) <= input(10);
output(1, 10) <= input(11);
output(1, 11) <= input(12);
output(1, 12) <= input(13);
output(1, 13) <= input(14);
output(1, 14) <= input(15);
output(1, 15) <= input(38);
output(1, 16) <= input(1);
output(1, 17) <= input(2);
output(1, 18) <= input(3);
output(1, 19) <= input(4);
output(1, 20) <= input(5);
output(1, 21) <= input(6);
output(1, 22) <= input(7);
output(1, 23) <= input(8);
output(1, 24) <= input(9);
output(1, 25) <= input(10);
output(1, 26) <= input(11);
output(1, 27) <= input(12);
output(1, 28) <= input(13);
output(1, 29) <= input(14);
output(1, 30) <= input(15);
output(1, 31) <= input(38);
output(1, 32) <= input(17);
output(1, 33) <= input(18);
output(1, 34) <= input(19);
output(1, 35) <= input(20);
output(1, 36) <= input(21);
output(1, 37) <= input(22);
output(1, 38) <= input(23);
output(1, 39) <= input(24);
output(1, 40) <= input(25);
output(1, 41) <= input(26);
output(1, 42) <= input(27);
output(1, 43) <= input(28);
output(1, 44) <= input(29);
output(1, 45) <= input(30);
output(1, 46) <= input(31);
output(1, 47) <= input(39);
output(1, 48) <= input(17);
output(1, 49) <= input(18);
output(1, 50) <= input(19);
output(1, 51) <= input(20);
output(1, 52) <= input(21);
output(1, 53) <= input(22);
output(1, 54) <= input(23);
output(1, 55) <= input(24);
output(1, 56) <= input(25);
output(1, 57) <= input(26);
output(1, 58) <= input(27);
output(1, 59) <= input(28);
output(1, 60) <= input(29);
output(1, 61) <= input(30);
output(1, 62) <= input(31);
output(1, 63) <= input(39);
output(1, 64) <= input(17);
output(1, 65) <= input(18);
output(1, 66) <= input(19);
output(1, 67) <= input(20);
output(1, 68) <= input(21);
output(1, 69) <= input(22);
output(1, 70) <= input(23);
output(1, 71) <= input(24);
output(1, 72) <= input(25);
output(1, 73) <= input(26);
output(1, 74) <= input(27);
output(1, 75) <= input(28);
output(1, 76) <= input(29);
output(1, 77) <= input(30);
output(1, 78) <= input(31);
output(1, 79) <= input(39);
output(1, 80) <= input(0);
output(1, 81) <= input(1);
output(1, 82) <= input(2);
output(1, 83) <= input(3);
output(1, 84) <= input(4);
output(1, 85) <= input(5);
output(1, 86) <= input(6);
output(1, 87) <= input(7);
output(1, 88) <= input(8);
output(1, 89) <= input(9);
output(1, 90) <= input(10);
output(1, 91) <= input(11);
output(1, 92) <= input(12);
output(1, 93) <= input(13);
output(1, 94) <= input(14);
output(1, 95) <= input(15);
output(1, 96) <= input(0);
output(1, 97) <= input(1);
output(1, 98) <= input(2);
output(1, 99) <= input(3);
output(1, 100) <= input(4);
output(1, 101) <= input(5);
output(1, 102) <= input(6);
output(1, 103) <= input(7);
output(1, 104) <= input(8);
output(1, 105) <= input(9);
output(1, 106) <= input(10);
output(1, 107) <= input(11);
output(1, 108) <= input(12);
output(1, 109) <= input(13);
output(1, 110) <= input(14);
output(1, 111) <= input(15);
output(1, 112) <= input(0);
output(1, 113) <= input(1);
output(1, 114) <= input(2);
output(1, 115) <= input(3);
output(1, 116) <= input(4);
output(1, 117) <= input(5);
output(1, 118) <= input(6);
output(1, 119) <= input(7);
output(1, 120) <= input(8);
output(1, 121) <= input(9);
output(1, 122) <= input(10);
output(1, 123) <= input(11);
output(1, 124) <= input(12);
output(1, 125) <= input(13);
output(1, 126) <= input(14);
output(1, 127) <= input(15);
output(1, 128) <= input(16);
output(1, 129) <= input(17);
output(1, 130) <= input(18);
output(1, 131) <= input(19);
output(1, 132) <= input(20);
output(1, 133) <= input(21);
output(1, 134) <= input(22);
output(1, 135) <= input(23);
output(1, 136) <= input(24);
output(1, 137) <= input(25);
output(1, 138) <= input(26);
output(1, 139) <= input(27);
output(1, 140) <= input(28);
output(1, 141) <= input(29);
output(1, 142) <= input(30);
output(1, 143) <= input(31);
output(1, 144) <= input(16);
output(1, 145) <= input(17);
output(1, 146) <= input(18);
output(1, 147) <= input(19);
output(1, 148) <= input(20);
output(1, 149) <= input(21);
output(1, 150) <= input(22);
output(1, 151) <= input(23);
output(1, 152) <= input(24);
output(1, 153) <= input(25);
output(1, 154) <= input(26);
output(1, 155) <= input(27);
output(1, 156) <= input(28);
output(1, 157) <= input(29);
output(1, 158) <= input(30);
output(1, 159) <= input(31);
output(1, 160) <= input(32);
output(1, 161) <= input(0);
output(1, 162) <= input(1);
output(1, 163) <= input(2);
output(1, 164) <= input(3);
output(1, 165) <= input(4);
output(1, 166) <= input(5);
output(1, 167) <= input(6);
output(1, 168) <= input(7);
output(1, 169) <= input(8);
output(1, 170) <= input(9);
output(1, 171) <= input(10);
output(1, 172) <= input(11);
output(1, 173) <= input(12);
output(1, 174) <= input(13);
output(1, 175) <= input(14);
output(1, 176) <= input(32);
output(1, 177) <= input(0);
output(1, 178) <= input(1);
output(1, 179) <= input(2);
output(1, 180) <= input(3);
output(1, 181) <= input(4);
output(1, 182) <= input(5);
output(1, 183) <= input(6);
output(1, 184) <= input(7);
output(1, 185) <= input(8);
output(1, 186) <= input(9);
output(1, 187) <= input(10);
output(1, 188) <= input(11);
output(1, 189) <= input(12);
output(1, 190) <= input(13);
output(1, 191) <= input(14);
output(1, 192) <= input(32);
output(1, 193) <= input(0);
output(1, 194) <= input(1);
output(1, 195) <= input(2);
output(1, 196) <= input(3);
output(1, 197) <= input(4);
output(1, 198) <= input(5);
output(1, 199) <= input(6);
output(1, 200) <= input(7);
output(1, 201) <= input(8);
output(1, 202) <= input(9);
output(1, 203) <= input(10);
output(1, 204) <= input(11);
output(1, 205) <= input(12);
output(1, 206) <= input(13);
output(1, 207) <= input(14);
output(1, 208) <= input(33);
output(1, 209) <= input(16);
output(1, 210) <= input(17);
output(1, 211) <= input(18);
output(1, 212) <= input(19);
output(1, 213) <= input(20);
output(1, 214) <= input(21);
output(1, 215) <= input(22);
output(1, 216) <= input(23);
output(1, 217) <= input(24);
output(1, 218) <= input(25);
output(1, 219) <= input(26);
output(1, 220) <= input(27);
output(1, 221) <= input(28);
output(1, 222) <= input(29);
output(1, 223) <= input(30);
output(1, 224) <= input(33);
output(1, 225) <= input(16);
output(1, 226) <= input(17);
output(1, 227) <= input(18);
output(1, 228) <= input(19);
output(1, 229) <= input(20);
output(1, 230) <= input(21);
output(1, 231) <= input(22);
output(1, 232) <= input(23);
output(1, 233) <= input(24);
output(1, 234) <= input(25);
output(1, 235) <= input(26);
output(1, 236) <= input(27);
output(1, 237) <= input(28);
output(1, 238) <= input(29);
output(1, 239) <= input(30);
output(1, 240) <= input(33);
output(1, 241) <= input(16);
output(1, 242) <= input(17);
output(1, 243) <= input(18);
output(1, 244) <= input(19);
output(1, 245) <= input(20);
output(1, 246) <= input(21);
output(1, 247) <= input(22);
output(1, 248) <= input(23);
output(1, 249) <= input(24);
output(1, 250) <= input(25);
output(1, 251) <= input(26);
output(1, 252) <= input(27);
output(1, 253) <= input(28);
output(1, 254) <= input(29);
output(1, 255) <= input(30);
output(2, 0) <= input(2);
output(2, 1) <= input(3);
output(2, 2) <= input(4);
output(2, 3) <= input(5);
output(2, 4) <= input(6);
output(2, 5) <= input(7);
output(2, 6) <= input(8);
output(2, 7) <= input(9);
output(2, 8) <= input(10);
output(2, 9) <= input(11);
output(2, 10) <= input(12);
output(2, 11) <= input(13);
output(2, 12) <= input(14);
output(2, 13) <= input(15);
output(2, 14) <= input(38);
output(2, 15) <= input(40);
output(2, 16) <= input(2);
output(2, 17) <= input(3);
output(2, 18) <= input(4);
output(2, 19) <= input(5);
output(2, 20) <= input(6);
output(2, 21) <= input(7);
output(2, 22) <= input(8);
output(2, 23) <= input(9);
output(2, 24) <= input(10);
output(2, 25) <= input(11);
output(2, 26) <= input(12);
output(2, 27) <= input(13);
output(2, 28) <= input(14);
output(2, 29) <= input(15);
output(2, 30) <= input(38);
output(2, 31) <= input(40);
output(2, 32) <= input(2);
output(2, 33) <= input(3);
output(2, 34) <= input(4);
output(2, 35) <= input(5);
output(2, 36) <= input(6);
output(2, 37) <= input(7);
output(2, 38) <= input(8);
output(2, 39) <= input(9);
output(2, 40) <= input(10);
output(2, 41) <= input(11);
output(2, 42) <= input(12);
output(2, 43) <= input(13);
output(2, 44) <= input(14);
output(2, 45) <= input(15);
output(2, 46) <= input(38);
output(2, 47) <= input(40);
output(2, 48) <= input(2);
output(2, 49) <= input(3);
output(2, 50) <= input(4);
output(2, 51) <= input(5);
output(2, 52) <= input(6);
output(2, 53) <= input(7);
output(2, 54) <= input(8);
output(2, 55) <= input(9);
output(2, 56) <= input(10);
output(2, 57) <= input(11);
output(2, 58) <= input(12);
output(2, 59) <= input(13);
output(2, 60) <= input(14);
output(2, 61) <= input(15);
output(2, 62) <= input(38);
output(2, 63) <= input(40);
output(2, 64) <= input(18);
output(2, 65) <= input(19);
output(2, 66) <= input(20);
output(2, 67) <= input(21);
output(2, 68) <= input(22);
output(2, 69) <= input(23);
output(2, 70) <= input(24);
output(2, 71) <= input(25);
output(2, 72) <= input(26);
output(2, 73) <= input(27);
output(2, 74) <= input(28);
output(2, 75) <= input(29);
output(2, 76) <= input(30);
output(2, 77) <= input(31);
output(2, 78) <= input(39);
output(2, 79) <= input(41);
output(2, 80) <= input(18);
output(2, 81) <= input(19);
output(2, 82) <= input(20);
output(2, 83) <= input(21);
output(2, 84) <= input(22);
output(2, 85) <= input(23);
output(2, 86) <= input(24);
output(2, 87) <= input(25);
output(2, 88) <= input(26);
output(2, 89) <= input(27);
output(2, 90) <= input(28);
output(2, 91) <= input(29);
output(2, 92) <= input(30);
output(2, 93) <= input(31);
output(2, 94) <= input(39);
output(2, 95) <= input(41);
output(2, 96) <= input(18);
output(2, 97) <= input(19);
output(2, 98) <= input(20);
output(2, 99) <= input(21);
output(2, 100) <= input(22);
output(2, 101) <= input(23);
output(2, 102) <= input(24);
output(2, 103) <= input(25);
output(2, 104) <= input(26);
output(2, 105) <= input(27);
output(2, 106) <= input(28);
output(2, 107) <= input(29);
output(2, 108) <= input(30);
output(2, 109) <= input(31);
output(2, 110) <= input(39);
output(2, 111) <= input(41);
output(2, 112) <= input(18);
output(2, 113) <= input(19);
output(2, 114) <= input(20);
output(2, 115) <= input(21);
output(2, 116) <= input(22);
output(2, 117) <= input(23);
output(2, 118) <= input(24);
output(2, 119) <= input(25);
output(2, 120) <= input(26);
output(2, 121) <= input(27);
output(2, 122) <= input(28);
output(2, 123) <= input(29);
output(2, 124) <= input(30);
output(2, 125) <= input(31);
output(2, 126) <= input(39);
output(2, 127) <= input(41);
output(2, 128) <= input(1);
output(2, 129) <= input(2);
output(2, 130) <= input(3);
output(2, 131) <= input(4);
output(2, 132) <= input(5);
output(2, 133) <= input(6);
output(2, 134) <= input(7);
output(2, 135) <= input(8);
output(2, 136) <= input(9);
output(2, 137) <= input(10);
output(2, 138) <= input(11);
output(2, 139) <= input(12);
output(2, 140) <= input(13);
output(2, 141) <= input(14);
output(2, 142) <= input(15);
output(2, 143) <= input(38);
output(2, 144) <= input(1);
output(2, 145) <= input(2);
output(2, 146) <= input(3);
output(2, 147) <= input(4);
output(2, 148) <= input(5);
output(2, 149) <= input(6);
output(2, 150) <= input(7);
output(2, 151) <= input(8);
output(2, 152) <= input(9);
output(2, 153) <= input(10);
output(2, 154) <= input(11);
output(2, 155) <= input(12);
output(2, 156) <= input(13);
output(2, 157) <= input(14);
output(2, 158) <= input(15);
output(2, 159) <= input(38);
output(2, 160) <= input(1);
output(2, 161) <= input(2);
output(2, 162) <= input(3);
output(2, 163) <= input(4);
output(2, 164) <= input(5);
output(2, 165) <= input(6);
output(2, 166) <= input(7);
output(2, 167) <= input(8);
output(2, 168) <= input(9);
output(2, 169) <= input(10);
output(2, 170) <= input(11);
output(2, 171) <= input(12);
output(2, 172) <= input(13);
output(2, 173) <= input(14);
output(2, 174) <= input(15);
output(2, 175) <= input(38);
output(2, 176) <= input(1);
output(2, 177) <= input(2);
output(2, 178) <= input(3);
output(2, 179) <= input(4);
output(2, 180) <= input(5);
output(2, 181) <= input(6);
output(2, 182) <= input(7);
output(2, 183) <= input(8);
output(2, 184) <= input(9);
output(2, 185) <= input(10);
output(2, 186) <= input(11);
output(2, 187) <= input(12);
output(2, 188) <= input(13);
output(2, 189) <= input(14);
output(2, 190) <= input(15);
output(2, 191) <= input(38);
output(2, 192) <= input(17);
output(2, 193) <= input(18);
output(2, 194) <= input(19);
output(2, 195) <= input(20);
output(2, 196) <= input(21);
output(2, 197) <= input(22);
output(2, 198) <= input(23);
output(2, 199) <= input(24);
output(2, 200) <= input(25);
output(2, 201) <= input(26);
output(2, 202) <= input(27);
output(2, 203) <= input(28);
output(2, 204) <= input(29);
output(2, 205) <= input(30);
output(2, 206) <= input(31);
output(2, 207) <= input(39);
output(2, 208) <= input(17);
output(2, 209) <= input(18);
output(2, 210) <= input(19);
output(2, 211) <= input(20);
output(2, 212) <= input(21);
output(2, 213) <= input(22);
output(2, 214) <= input(23);
output(2, 215) <= input(24);
output(2, 216) <= input(25);
output(2, 217) <= input(26);
output(2, 218) <= input(27);
output(2, 219) <= input(28);
output(2, 220) <= input(29);
output(2, 221) <= input(30);
output(2, 222) <= input(31);
output(2, 223) <= input(39);
output(2, 224) <= input(17);
output(2, 225) <= input(18);
output(2, 226) <= input(19);
output(2, 227) <= input(20);
output(2, 228) <= input(21);
output(2, 229) <= input(22);
output(2, 230) <= input(23);
output(2, 231) <= input(24);
output(2, 232) <= input(25);
output(2, 233) <= input(26);
output(2, 234) <= input(27);
output(2, 235) <= input(28);
output(2, 236) <= input(29);
output(2, 237) <= input(30);
output(2, 238) <= input(31);
output(2, 239) <= input(39);
output(2, 240) <= input(17);
output(2, 241) <= input(18);
output(2, 242) <= input(19);
output(2, 243) <= input(20);
output(2, 244) <= input(21);
output(2, 245) <= input(22);
output(2, 246) <= input(23);
output(2, 247) <= input(24);
output(2, 248) <= input(25);
output(2, 249) <= input(26);
output(2, 250) <= input(27);
output(2, 251) <= input(28);
output(2, 252) <= input(29);
output(2, 253) <= input(30);
output(2, 254) <= input(31);
output(2, 255) <= input(39);
when "1101" =>
output(0, 0) <= input(0);
output(0, 1) <= input(1);
output(0, 2) <= input(2);
output(0, 3) <= input(3);
output(0, 4) <= input(4);
output(0, 5) <= input(5);
output(0, 6) <= input(6);
output(0, 7) <= input(7);
output(0, 8) <= input(8);
output(0, 9) <= input(9);
output(0, 10) <= input(10);
output(0, 11) <= input(11);
output(0, 12) <= input(12);
output(0, 13) <= input(13);
output(0, 14) <= input(14);
output(0, 15) <= input(15);
output(0, 16) <= input(0);
output(0, 17) <= input(1);
output(0, 18) <= input(2);
output(0, 19) <= input(3);
output(0, 20) <= input(4);
output(0, 21) <= input(5);
output(0, 22) <= input(6);
output(0, 23) <= input(7);
output(0, 24) <= input(8);
output(0, 25) <= input(9);
output(0, 26) <= input(10);
output(0, 27) <= input(11);
output(0, 28) <= input(12);
output(0, 29) <= input(13);
output(0, 30) <= input(14);
output(0, 31) <= input(15);
output(0, 32) <= input(0);
output(0, 33) <= input(1);
output(0, 34) <= input(2);
output(0, 35) <= input(3);
output(0, 36) <= input(4);
output(0, 37) <= input(5);
output(0, 38) <= input(6);
output(0, 39) <= input(7);
output(0, 40) <= input(8);
output(0, 41) <= input(9);
output(0, 42) <= input(10);
output(0, 43) <= input(11);
output(0, 44) <= input(12);
output(0, 45) <= input(13);
output(0, 46) <= input(14);
output(0, 47) <= input(15);
output(0, 48) <= input(0);
output(0, 49) <= input(1);
output(0, 50) <= input(2);
output(0, 51) <= input(3);
output(0, 52) <= input(4);
output(0, 53) <= input(5);
output(0, 54) <= input(6);
output(0, 55) <= input(7);
output(0, 56) <= input(8);
output(0, 57) <= input(9);
output(0, 58) <= input(10);
output(0, 59) <= input(11);
output(0, 60) <= input(12);
output(0, 61) <= input(13);
output(0, 62) <= input(14);
output(0, 63) <= input(15);
output(0, 64) <= input(0);
output(0, 65) <= input(1);
output(0, 66) <= input(2);
output(0, 67) <= input(3);
output(0, 68) <= input(4);
output(0, 69) <= input(5);
output(0, 70) <= input(6);
output(0, 71) <= input(7);
output(0, 72) <= input(8);
output(0, 73) <= input(9);
output(0, 74) <= input(10);
output(0, 75) <= input(11);
output(0, 76) <= input(12);
output(0, 77) <= input(13);
output(0, 78) <= input(14);
output(0, 79) <= input(15);
output(0, 80) <= input(16);
output(0, 81) <= input(17);
output(0, 82) <= input(18);
output(0, 83) <= input(19);
output(0, 84) <= input(20);
output(0, 85) <= input(21);
output(0, 86) <= input(22);
output(0, 87) <= input(23);
output(0, 88) <= input(24);
output(0, 89) <= input(25);
output(0, 90) <= input(26);
output(0, 91) <= input(27);
output(0, 92) <= input(28);
output(0, 93) <= input(29);
output(0, 94) <= input(30);
output(0, 95) <= input(31);
output(0, 96) <= input(16);
output(0, 97) <= input(17);
output(0, 98) <= input(18);
output(0, 99) <= input(19);
output(0, 100) <= input(20);
output(0, 101) <= input(21);
output(0, 102) <= input(22);
output(0, 103) <= input(23);
output(0, 104) <= input(24);
output(0, 105) <= input(25);
output(0, 106) <= input(26);
output(0, 107) <= input(27);
output(0, 108) <= input(28);
output(0, 109) <= input(29);
output(0, 110) <= input(30);
output(0, 111) <= input(31);
output(0, 112) <= input(16);
output(0, 113) <= input(17);
output(0, 114) <= input(18);
output(0, 115) <= input(19);
output(0, 116) <= input(20);
output(0, 117) <= input(21);
output(0, 118) <= input(22);
output(0, 119) <= input(23);
output(0, 120) <= input(24);
output(0, 121) <= input(25);
output(0, 122) <= input(26);
output(0, 123) <= input(27);
output(0, 124) <= input(28);
output(0, 125) <= input(29);
output(0, 126) <= input(30);
output(0, 127) <= input(31);
output(0, 128) <= input(16);
output(0, 129) <= input(17);
output(0, 130) <= input(18);
output(0, 131) <= input(19);
output(0, 132) <= input(20);
output(0, 133) <= input(21);
output(0, 134) <= input(22);
output(0, 135) <= input(23);
output(0, 136) <= input(24);
output(0, 137) <= input(25);
output(0, 138) <= input(26);
output(0, 139) <= input(27);
output(0, 140) <= input(28);
output(0, 141) <= input(29);
output(0, 142) <= input(30);
output(0, 143) <= input(31);
output(0, 144) <= input(16);
output(0, 145) <= input(17);
output(0, 146) <= input(18);
output(0, 147) <= input(19);
output(0, 148) <= input(20);
output(0, 149) <= input(21);
output(0, 150) <= input(22);
output(0, 151) <= input(23);
output(0, 152) <= input(24);
output(0, 153) <= input(25);
output(0, 154) <= input(26);
output(0, 155) <= input(27);
output(0, 156) <= input(28);
output(0, 157) <= input(29);
output(0, 158) <= input(30);
output(0, 159) <= input(31);
output(0, 160) <= input(32);
output(0, 161) <= input(0);
output(0, 162) <= input(1);
output(0, 163) <= input(2);
output(0, 164) <= input(3);
output(0, 165) <= input(4);
output(0, 166) <= input(5);
output(0, 167) <= input(6);
output(0, 168) <= input(7);
output(0, 169) <= input(8);
output(0, 170) <= input(9);
output(0, 171) <= input(10);
output(0, 172) <= input(11);
output(0, 173) <= input(12);
output(0, 174) <= input(13);
output(0, 175) <= input(14);
output(0, 176) <= input(32);
output(0, 177) <= input(0);
output(0, 178) <= input(1);
output(0, 179) <= input(2);
output(0, 180) <= input(3);
output(0, 181) <= input(4);
output(0, 182) <= input(5);
output(0, 183) <= input(6);
output(0, 184) <= input(7);
output(0, 185) <= input(8);
output(0, 186) <= input(9);
output(0, 187) <= input(10);
output(0, 188) <= input(11);
output(0, 189) <= input(12);
output(0, 190) <= input(13);
output(0, 191) <= input(14);
output(0, 192) <= input(32);
output(0, 193) <= input(0);
output(0, 194) <= input(1);
output(0, 195) <= input(2);
output(0, 196) <= input(3);
output(0, 197) <= input(4);
output(0, 198) <= input(5);
output(0, 199) <= input(6);
output(0, 200) <= input(7);
output(0, 201) <= input(8);
output(0, 202) <= input(9);
output(0, 203) <= input(10);
output(0, 204) <= input(11);
output(0, 205) <= input(12);
output(0, 206) <= input(13);
output(0, 207) <= input(14);
output(0, 208) <= input(32);
output(0, 209) <= input(0);
output(0, 210) <= input(1);
output(0, 211) <= input(2);
output(0, 212) <= input(3);
output(0, 213) <= input(4);
output(0, 214) <= input(5);
output(0, 215) <= input(6);
output(0, 216) <= input(7);
output(0, 217) <= input(8);
output(0, 218) <= input(9);
output(0, 219) <= input(10);
output(0, 220) <= input(11);
output(0, 221) <= input(12);
output(0, 222) <= input(13);
output(0, 223) <= input(14);
output(0, 224) <= input(32);
output(0, 225) <= input(0);
output(0, 226) <= input(1);
output(0, 227) <= input(2);
output(0, 228) <= input(3);
output(0, 229) <= input(4);
output(0, 230) <= input(5);
output(0, 231) <= input(6);
output(0, 232) <= input(7);
output(0, 233) <= input(8);
output(0, 234) <= input(9);
output(0, 235) <= input(10);
output(0, 236) <= input(11);
output(0, 237) <= input(12);
output(0, 238) <= input(13);
output(0, 239) <= input(14);
output(0, 240) <= input(32);
output(0, 241) <= input(0);
output(0, 242) <= input(1);
output(0, 243) <= input(2);
output(0, 244) <= input(3);
output(0, 245) <= input(4);
output(0, 246) <= input(5);
output(0, 247) <= input(6);
output(0, 248) <= input(7);
output(0, 249) <= input(8);
output(0, 250) <= input(9);
output(0, 251) <= input(10);
output(0, 252) <= input(11);
output(0, 253) <= input(12);
output(0, 254) <= input(13);
output(0, 255) <= input(14);
output(1, 0) <= input(17);
output(1, 1) <= input(18);
output(1, 2) <= input(19);
output(1, 3) <= input(20);
output(1, 4) <= input(21);
output(1, 5) <= input(22);
output(1, 6) <= input(23);
output(1, 7) <= input(24);
output(1, 8) <= input(25);
output(1, 9) <= input(26);
output(1, 10) <= input(27);
output(1, 11) <= input(28);
output(1, 12) <= input(29);
output(1, 13) <= input(30);
output(1, 14) <= input(31);
output(1, 15) <= input(33);
output(1, 16) <= input(17);
output(1, 17) <= input(18);
output(1, 18) <= input(19);
output(1, 19) <= input(20);
output(1, 20) <= input(21);
output(1, 21) <= input(22);
output(1, 22) <= input(23);
output(1, 23) <= input(24);
output(1, 24) <= input(25);
output(1, 25) <= input(26);
output(1, 26) <= input(27);
output(1, 27) <= input(28);
output(1, 28) <= input(29);
output(1, 29) <= input(30);
output(1, 30) <= input(31);
output(1, 31) <= input(33);
output(1, 32) <= input(17);
output(1, 33) <= input(18);
output(1, 34) <= input(19);
output(1, 35) <= input(20);
output(1, 36) <= input(21);
output(1, 37) <= input(22);
output(1, 38) <= input(23);
output(1, 39) <= input(24);
output(1, 40) <= input(25);
output(1, 41) <= input(26);
output(1, 42) <= input(27);
output(1, 43) <= input(28);
output(1, 44) <= input(29);
output(1, 45) <= input(30);
output(1, 46) <= input(31);
output(1, 47) <= input(33);
output(1, 48) <= input(17);
output(1, 49) <= input(18);
output(1, 50) <= input(19);
output(1, 51) <= input(20);
output(1, 52) <= input(21);
output(1, 53) <= input(22);
output(1, 54) <= input(23);
output(1, 55) <= input(24);
output(1, 56) <= input(25);
output(1, 57) <= input(26);
output(1, 58) <= input(27);
output(1, 59) <= input(28);
output(1, 60) <= input(29);
output(1, 61) <= input(30);
output(1, 62) <= input(31);
output(1, 63) <= input(33);
output(1, 64) <= input(17);
output(1, 65) <= input(18);
output(1, 66) <= input(19);
output(1, 67) <= input(20);
output(1, 68) <= input(21);
output(1, 69) <= input(22);
output(1, 70) <= input(23);
output(1, 71) <= input(24);
output(1, 72) <= input(25);
output(1, 73) <= input(26);
output(1, 74) <= input(27);
output(1, 75) <= input(28);
output(1, 76) <= input(29);
output(1, 77) <= input(30);
output(1, 78) <= input(31);
output(1, 79) <= input(33);
output(1, 80) <= input(17);
output(1, 81) <= input(18);
output(1, 82) <= input(19);
output(1, 83) <= input(20);
output(1, 84) <= input(21);
output(1, 85) <= input(22);
output(1, 86) <= input(23);
output(1, 87) <= input(24);
output(1, 88) <= input(25);
output(1, 89) <= input(26);
output(1, 90) <= input(27);
output(1, 91) <= input(28);
output(1, 92) <= input(29);
output(1, 93) <= input(30);
output(1, 94) <= input(31);
output(1, 95) <= input(33);
output(1, 96) <= input(17);
output(1, 97) <= input(18);
output(1, 98) <= input(19);
output(1, 99) <= input(20);
output(1, 100) <= input(21);
output(1, 101) <= input(22);
output(1, 102) <= input(23);
output(1, 103) <= input(24);
output(1, 104) <= input(25);
output(1, 105) <= input(26);
output(1, 106) <= input(27);
output(1, 107) <= input(28);
output(1, 108) <= input(29);
output(1, 109) <= input(30);
output(1, 110) <= input(31);
output(1, 111) <= input(33);
output(1, 112) <= input(17);
output(1, 113) <= input(18);
output(1, 114) <= input(19);
output(1, 115) <= input(20);
output(1, 116) <= input(21);
output(1, 117) <= input(22);
output(1, 118) <= input(23);
output(1, 119) <= input(24);
output(1, 120) <= input(25);
output(1, 121) <= input(26);
output(1, 122) <= input(27);
output(1, 123) <= input(28);
output(1, 124) <= input(29);
output(1, 125) <= input(30);
output(1, 126) <= input(31);
output(1, 127) <= input(33);
output(1, 128) <= input(0);
output(1, 129) <= input(1);
output(1, 130) <= input(2);
output(1, 131) <= input(3);
output(1, 132) <= input(4);
output(1, 133) <= input(5);
output(1, 134) <= input(6);
output(1, 135) <= input(7);
output(1, 136) <= input(8);
output(1, 137) <= input(9);
output(1, 138) <= input(10);
output(1, 139) <= input(11);
output(1, 140) <= input(12);
output(1, 141) <= input(13);
output(1, 142) <= input(14);
output(1, 143) <= input(15);
output(1, 144) <= input(0);
output(1, 145) <= input(1);
output(1, 146) <= input(2);
output(1, 147) <= input(3);
output(1, 148) <= input(4);
output(1, 149) <= input(5);
output(1, 150) <= input(6);
output(1, 151) <= input(7);
output(1, 152) <= input(8);
output(1, 153) <= input(9);
output(1, 154) <= input(10);
output(1, 155) <= input(11);
output(1, 156) <= input(12);
output(1, 157) <= input(13);
output(1, 158) <= input(14);
output(1, 159) <= input(15);
output(1, 160) <= input(0);
output(1, 161) <= input(1);
output(1, 162) <= input(2);
output(1, 163) <= input(3);
output(1, 164) <= input(4);
output(1, 165) <= input(5);
output(1, 166) <= input(6);
output(1, 167) <= input(7);
output(1, 168) <= input(8);
output(1, 169) <= input(9);
output(1, 170) <= input(10);
output(1, 171) <= input(11);
output(1, 172) <= input(12);
output(1, 173) <= input(13);
output(1, 174) <= input(14);
output(1, 175) <= input(15);
output(1, 176) <= input(0);
output(1, 177) <= input(1);
output(1, 178) <= input(2);
output(1, 179) <= input(3);
output(1, 180) <= input(4);
output(1, 181) <= input(5);
output(1, 182) <= input(6);
output(1, 183) <= input(7);
output(1, 184) <= input(8);
output(1, 185) <= input(9);
output(1, 186) <= input(10);
output(1, 187) <= input(11);
output(1, 188) <= input(12);
output(1, 189) <= input(13);
output(1, 190) <= input(14);
output(1, 191) <= input(15);
output(1, 192) <= input(0);
output(1, 193) <= input(1);
output(1, 194) <= input(2);
output(1, 195) <= input(3);
output(1, 196) <= input(4);
output(1, 197) <= input(5);
output(1, 198) <= input(6);
output(1, 199) <= input(7);
output(1, 200) <= input(8);
output(1, 201) <= input(9);
output(1, 202) <= input(10);
output(1, 203) <= input(11);
output(1, 204) <= input(12);
output(1, 205) <= input(13);
output(1, 206) <= input(14);
output(1, 207) <= input(15);
output(1, 208) <= input(0);
output(1, 209) <= input(1);
output(1, 210) <= input(2);
output(1, 211) <= input(3);
output(1, 212) <= input(4);
output(1, 213) <= input(5);
output(1, 214) <= input(6);
output(1, 215) <= input(7);
output(1, 216) <= input(8);
output(1, 217) <= input(9);
output(1, 218) <= input(10);
output(1, 219) <= input(11);
output(1, 220) <= input(12);
output(1, 221) <= input(13);
output(1, 222) <= input(14);
output(1, 223) <= input(15);
output(1, 224) <= input(0);
output(1, 225) <= input(1);
output(1, 226) <= input(2);
output(1, 227) <= input(3);
output(1, 228) <= input(4);
output(1, 229) <= input(5);
output(1, 230) <= input(6);
output(1, 231) <= input(7);
output(1, 232) <= input(8);
output(1, 233) <= input(9);
output(1, 234) <= input(10);
output(1, 235) <= input(11);
output(1, 236) <= input(12);
output(1, 237) <= input(13);
output(1, 238) <= input(14);
output(1, 239) <= input(15);
output(1, 240) <= input(0);
output(1, 241) <= input(1);
output(1, 242) <= input(2);
output(1, 243) <= input(3);
output(1, 244) <= input(4);
output(1, 245) <= input(5);
output(1, 246) <= input(6);
output(1, 247) <= input(7);
output(1, 248) <= input(8);
output(1, 249) <= input(9);
output(1, 250) <= input(10);
output(1, 251) <= input(11);
output(1, 252) <= input(12);
output(1, 253) <= input(13);
output(1, 254) <= input(14);
output(1, 255) <= input(15);
output(2, 0) <= input(1);
output(2, 1) <= input(2);
output(2, 2) <= input(3);
output(2, 3) <= input(4);
output(2, 4) <= input(5);
output(2, 5) <= input(6);
output(2, 6) <= input(7);
output(2, 7) <= input(8);
output(2, 8) <= input(9);
output(2, 9) <= input(10);
output(2, 10) <= input(11);
output(2, 11) <= input(12);
output(2, 12) <= input(13);
output(2, 13) <= input(14);
output(2, 14) <= input(15);
output(2, 15) <= input(34);
output(2, 16) <= input(1);
output(2, 17) <= input(2);
output(2, 18) <= input(3);
output(2, 19) <= input(4);
output(2, 20) <= input(5);
output(2, 21) <= input(6);
output(2, 22) <= input(7);
output(2, 23) <= input(8);
output(2, 24) <= input(9);
output(2, 25) <= input(10);
output(2, 26) <= input(11);
output(2, 27) <= input(12);
output(2, 28) <= input(13);
output(2, 29) <= input(14);
output(2, 30) <= input(15);
output(2, 31) <= input(34);
output(2, 32) <= input(1);
output(2, 33) <= input(2);
output(2, 34) <= input(3);
output(2, 35) <= input(4);
output(2, 36) <= input(5);
output(2, 37) <= input(6);
output(2, 38) <= input(7);
output(2, 39) <= input(8);
output(2, 40) <= input(9);
output(2, 41) <= input(10);
output(2, 42) <= input(11);
output(2, 43) <= input(12);
output(2, 44) <= input(13);
output(2, 45) <= input(14);
output(2, 46) <= input(15);
output(2, 47) <= input(34);
output(2, 48) <= input(1);
output(2, 49) <= input(2);
output(2, 50) <= input(3);
output(2, 51) <= input(4);
output(2, 52) <= input(5);
output(2, 53) <= input(6);
output(2, 54) <= input(7);
output(2, 55) <= input(8);
output(2, 56) <= input(9);
output(2, 57) <= input(10);
output(2, 58) <= input(11);
output(2, 59) <= input(12);
output(2, 60) <= input(13);
output(2, 61) <= input(14);
output(2, 62) <= input(15);
output(2, 63) <= input(34);
output(2, 64) <= input(1);
output(2, 65) <= input(2);
output(2, 66) <= input(3);
output(2, 67) <= input(4);
output(2, 68) <= input(5);
output(2, 69) <= input(6);
output(2, 70) <= input(7);
output(2, 71) <= input(8);
output(2, 72) <= input(9);
output(2, 73) <= input(10);
output(2, 74) <= input(11);
output(2, 75) <= input(12);
output(2, 76) <= input(13);
output(2, 77) <= input(14);
output(2, 78) <= input(15);
output(2, 79) <= input(34);
output(2, 80) <= input(1);
output(2, 81) <= input(2);
output(2, 82) <= input(3);
output(2, 83) <= input(4);
output(2, 84) <= input(5);
output(2, 85) <= input(6);
output(2, 86) <= input(7);
output(2, 87) <= input(8);
output(2, 88) <= input(9);
output(2, 89) <= input(10);
output(2, 90) <= input(11);
output(2, 91) <= input(12);
output(2, 92) <= input(13);
output(2, 93) <= input(14);
output(2, 94) <= input(15);
output(2, 95) <= input(34);
output(2, 96) <= input(1);
output(2, 97) <= input(2);
output(2, 98) <= input(3);
output(2, 99) <= input(4);
output(2, 100) <= input(5);
output(2, 101) <= input(6);
output(2, 102) <= input(7);
output(2, 103) <= input(8);
output(2, 104) <= input(9);
output(2, 105) <= input(10);
output(2, 106) <= input(11);
output(2, 107) <= input(12);
output(2, 108) <= input(13);
output(2, 109) <= input(14);
output(2, 110) <= input(15);
output(2, 111) <= input(34);
output(2, 112) <= input(1);
output(2, 113) <= input(2);
output(2, 114) <= input(3);
output(2, 115) <= input(4);
output(2, 116) <= input(5);
output(2, 117) <= input(6);
output(2, 118) <= input(7);
output(2, 119) <= input(8);
output(2, 120) <= input(9);
output(2, 121) <= input(10);
output(2, 122) <= input(11);
output(2, 123) <= input(12);
output(2, 124) <= input(13);
output(2, 125) <= input(14);
output(2, 126) <= input(15);
output(2, 127) <= input(34);
output(2, 128) <= input(1);
output(2, 129) <= input(2);
output(2, 130) <= input(3);
output(2, 131) <= input(4);
output(2, 132) <= input(5);
output(2, 133) <= input(6);
output(2, 134) <= input(7);
output(2, 135) <= input(8);
output(2, 136) <= input(9);
output(2, 137) <= input(10);
output(2, 138) <= input(11);
output(2, 139) <= input(12);
output(2, 140) <= input(13);
output(2, 141) <= input(14);
output(2, 142) <= input(15);
output(2, 143) <= input(34);
output(2, 144) <= input(1);
output(2, 145) <= input(2);
output(2, 146) <= input(3);
output(2, 147) <= input(4);
output(2, 148) <= input(5);
output(2, 149) <= input(6);
output(2, 150) <= input(7);
output(2, 151) <= input(8);
output(2, 152) <= input(9);
output(2, 153) <= input(10);
output(2, 154) <= input(11);
output(2, 155) <= input(12);
output(2, 156) <= input(13);
output(2, 157) <= input(14);
output(2, 158) <= input(15);
output(2, 159) <= input(34);
output(2, 160) <= input(1);
output(2, 161) <= input(2);
output(2, 162) <= input(3);
output(2, 163) <= input(4);
output(2, 164) <= input(5);
output(2, 165) <= input(6);
output(2, 166) <= input(7);
output(2, 167) <= input(8);
output(2, 168) <= input(9);
output(2, 169) <= input(10);
output(2, 170) <= input(11);
output(2, 171) <= input(12);
output(2, 172) <= input(13);
output(2, 173) <= input(14);
output(2, 174) <= input(15);
output(2, 175) <= input(34);
output(2, 176) <= input(1);
output(2, 177) <= input(2);
output(2, 178) <= input(3);
output(2, 179) <= input(4);
output(2, 180) <= input(5);
output(2, 181) <= input(6);
output(2, 182) <= input(7);
output(2, 183) <= input(8);
output(2, 184) <= input(9);
output(2, 185) <= input(10);
output(2, 186) <= input(11);
output(2, 187) <= input(12);
output(2, 188) <= input(13);
output(2, 189) <= input(14);
output(2, 190) <= input(15);
output(2, 191) <= input(34);
output(2, 192) <= input(1);
output(2, 193) <= input(2);
output(2, 194) <= input(3);
output(2, 195) <= input(4);
output(2, 196) <= input(5);
output(2, 197) <= input(6);
output(2, 198) <= input(7);
output(2, 199) <= input(8);
output(2, 200) <= input(9);
output(2, 201) <= input(10);
output(2, 202) <= input(11);
output(2, 203) <= input(12);
output(2, 204) <= input(13);
output(2, 205) <= input(14);
output(2, 206) <= input(15);
output(2, 207) <= input(34);
output(2, 208) <= input(1);
output(2, 209) <= input(2);
output(2, 210) <= input(3);
output(2, 211) <= input(4);
output(2, 212) <= input(5);
output(2, 213) <= input(6);
output(2, 214) <= input(7);
output(2, 215) <= input(8);
output(2, 216) <= input(9);
output(2, 217) <= input(10);
output(2, 218) <= input(11);
output(2, 219) <= input(12);
output(2, 220) <= input(13);
output(2, 221) <= input(14);
output(2, 222) <= input(15);
output(2, 223) <= input(34);
output(2, 224) <= input(1);
output(2, 225) <= input(2);
output(2, 226) <= input(3);
output(2, 227) <= input(4);
output(2, 228) <= input(5);
output(2, 229) <= input(6);
output(2, 230) <= input(7);
output(2, 231) <= input(8);
output(2, 232) <= input(9);
output(2, 233) <= input(10);
output(2, 234) <= input(11);
output(2, 235) <= input(12);
output(2, 236) <= input(13);
output(2, 237) <= input(14);
output(2, 238) <= input(15);
output(2, 239) <= input(34);
output(2, 240) <= input(1);
output(2, 241) <= input(2);
output(2, 242) <= input(3);
output(2, 243) <= input(4);
output(2, 244) <= input(5);
output(2, 245) <= input(6);
output(2, 246) <= input(7);
output(2, 247) <= input(8);
output(2, 248) <= input(9);
output(2, 249) <= input(10);
output(2, 250) <= input(11);
output(2, 251) <= input(12);
output(2, 252) <= input(13);
output(2, 253) <= input(14);
output(2, 254) <= input(15);
output(2, 255) <= input(34);
output(3, 0) <= input(2);
output(3, 1) <= input(3);
output(3, 2) <= input(4);
output(3, 3) <= input(5);
output(3, 4) <= input(6);
output(3, 5) <= input(7);
output(3, 6) <= input(8);
output(3, 7) <= input(9);
output(3, 8) <= input(10);
output(3, 9) <= input(11);
output(3, 10) <= input(12);
output(3, 11) <= input(13);
output(3, 12) <= input(14);
output(3, 13) <= input(15);
output(3, 14) <= input(34);
output(3, 15) <= input(35);
output(3, 16) <= input(2);
output(3, 17) <= input(3);
output(3, 18) <= input(4);
output(3, 19) <= input(5);
output(3, 20) <= input(6);
output(3, 21) <= input(7);
output(3, 22) <= input(8);
output(3, 23) <= input(9);
output(3, 24) <= input(10);
output(3, 25) <= input(11);
output(3, 26) <= input(12);
output(3, 27) <= input(13);
output(3, 28) <= input(14);
output(3, 29) <= input(15);
output(3, 30) <= input(34);
output(3, 31) <= input(35);
output(3, 32) <= input(2);
output(3, 33) <= input(3);
output(3, 34) <= input(4);
output(3, 35) <= input(5);
output(3, 36) <= input(6);
output(3, 37) <= input(7);
output(3, 38) <= input(8);
output(3, 39) <= input(9);
output(3, 40) <= input(10);
output(3, 41) <= input(11);
output(3, 42) <= input(12);
output(3, 43) <= input(13);
output(3, 44) <= input(14);
output(3, 45) <= input(15);
output(3, 46) <= input(34);
output(3, 47) <= input(35);
output(3, 48) <= input(2);
output(3, 49) <= input(3);
output(3, 50) <= input(4);
output(3, 51) <= input(5);
output(3, 52) <= input(6);
output(3, 53) <= input(7);
output(3, 54) <= input(8);
output(3, 55) <= input(9);
output(3, 56) <= input(10);
output(3, 57) <= input(11);
output(3, 58) <= input(12);
output(3, 59) <= input(13);
output(3, 60) <= input(14);
output(3, 61) <= input(15);
output(3, 62) <= input(34);
output(3, 63) <= input(35);
output(3, 64) <= input(2);
output(3, 65) <= input(3);
output(3, 66) <= input(4);
output(3, 67) <= input(5);
output(3, 68) <= input(6);
output(3, 69) <= input(7);
output(3, 70) <= input(8);
output(3, 71) <= input(9);
output(3, 72) <= input(10);
output(3, 73) <= input(11);
output(3, 74) <= input(12);
output(3, 75) <= input(13);
output(3, 76) <= input(14);
output(3, 77) <= input(15);
output(3, 78) <= input(34);
output(3, 79) <= input(35);
output(3, 80) <= input(2);
output(3, 81) <= input(3);
output(3, 82) <= input(4);
output(3, 83) <= input(5);
output(3, 84) <= input(6);
output(3, 85) <= input(7);
output(3, 86) <= input(8);
output(3, 87) <= input(9);
output(3, 88) <= input(10);
output(3, 89) <= input(11);
output(3, 90) <= input(12);
output(3, 91) <= input(13);
output(3, 92) <= input(14);
output(3, 93) <= input(15);
output(3, 94) <= input(34);
output(3, 95) <= input(35);
output(3, 96) <= input(2);
output(3, 97) <= input(3);
output(3, 98) <= input(4);
output(3, 99) <= input(5);
output(3, 100) <= input(6);
output(3, 101) <= input(7);
output(3, 102) <= input(8);
output(3, 103) <= input(9);
output(3, 104) <= input(10);
output(3, 105) <= input(11);
output(3, 106) <= input(12);
output(3, 107) <= input(13);
output(3, 108) <= input(14);
output(3, 109) <= input(15);
output(3, 110) <= input(34);
output(3, 111) <= input(35);
output(3, 112) <= input(2);
output(3, 113) <= input(3);
output(3, 114) <= input(4);
output(3, 115) <= input(5);
output(3, 116) <= input(6);
output(3, 117) <= input(7);
output(3, 118) <= input(8);
output(3, 119) <= input(9);
output(3, 120) <= input(10);
output(3, 121) <= input(11);
output(3, 122) <= input(12);
output(3, 123) <= input(13);
output(3, 124) <= input(14);
output(3, 125) <= input(15);
output(3, 126) <= input(34);
output(3, 127) <= input(35);
output(3, 128) <= input(2);
output(3, 129) <= input(3);
output(3, 130) <= input(4);
output(3, 131) <= input(5);
output(3, 132) <= input(6);
output(3, 133) <= input(7);
output(3, 134) <= input(8);
output(3, 135) <= input(9);
output(3, 136) <= input(10);
output(3, 137) <= input(11);
output(3, 138) <= input(12);
output(3, 139) <= input(13);
output(3, 140) <= input(14);
output(3, 141) <= input(15);
output(3, 142) <= input(34);
output(3, 143) <= input(35);
output(3, 144) <= input(2);
output(3, 145) <= input(3);
output(3, 146) <= input(4);
output(3, 147) <= input(5);
output(3, 148) <= input(6);
output(3, 149) <= input(7);
output(3, 150) <= input(8);
output(3, 151) <= input(9);
output(3, 152) <= input(10);
output(3, 153) <= input(11);
output(3, 154) <= input(12);
output(3, 155) <= input(13);
output(3, 156) <= input(14);
output(3, 157) <= input(15);
output(3, 158) <= input(34);
output(3, 159) <= input(35);
output(3, 160) <= input(2);
output(3, 161) <= input(3);
output(3, 162) <= input(4);
output(3, 163) <= input(5);
output(3, 164) <= input(6);
output(3, 165) <= input(7);
output(3, 166) <= input(8);
output(3, 167) <= input(9);
output(3, 168) <= input(10);
output(3, 169) <= input(11);
output(3, 170) <= input(12);
output(3, 171) <= input(13);
output(3, 172) <= input(14);
output(3, 173) <= input(15);
output(3, 174) <= input(34);
output(3, 175) <= input(35);
output(3, 176) <= input(2);
output(3, 177) <= input(3);
output(3, 178) <= input(4);
output(3, 179) <= input(5);
output(3, 180) <= input(6);
output(3, 181) <= input(7);
output(3, 182) <= input(8);
output(3, 183) <= input(9);
output(3, 184) <= input(10);
output(3, 185) <= input(11);
output(3, 186) <= input(12);
output(3, 187) <= input(13);
output(3, 188) <= input(14);
output(3, 189) <= input(15);
output(3, 190) <= input(34);
output(3, 191) <= input(35);
output(3, 192) <= input(2);
output(3, 193) <= input(3);
output(3, 194) <= input(4);
output(3, 195) <= input(5);
output(3, 196) <= input(6);
output(3, 197) <= input(7);
output(3, 198) <= input(8);
output(3, 199) <= input(9);
output(3, 200) <= input(10);
output(3, 201) <= input(11);
output(3, 202) <= input(12);
output(3, 203) <= input(13);
output(3, 204) <= input(14);
output(3, 205) <= input(15);
output(3, 206) <= input(34);
output(3, 207) <= input(35);
output(3, 208) <= input(2);
output(3, 209) <= input(3);
output(3, 210) <= input(4);
output(3, 211) <= input(5);
output(3, 212) <= input(6);
output(3, 213) <= input(7);
output(3, 214) <= input(8);
output(3, 215) <= input(9);
output(3, 216) <= input(10);
output(3, 217) <= input(11);
output(3, 218) <= input(12);
output(3, 219) <= input(13);
output(3, 220) <= input(14);
output(3, 221) <= input(15);
output(3, 222) <= input(34);
output(3, 223) <= input(35);
output(3, 224) <= input(2);
output(3, 225) <= input(3);
output(3, 226) <= input(4);
output(3, 227) <= input(5);
output(3, 228) <= input(6);
output(3, 229) <= input(7);
output(3, 230) <= input(8);
output(3, 231) <= input(9);
output(3, 232) <= input(10);
output(3, 233) <= input(11);
output(3, 234) <= input(12);
output(3, 235) <= input(13);
output(3, 236) <= input(14);
output(3, 237) <= input(15);
output(3, 238) <= input(34);
output(3, 239) <= input(35);
output(3, 240) <= input(2);
output(3, 241) <= input(3);
output(3, 242) <= input(4);
output(3, 243) <= input(5);
output(3, 244) <= input(6);
output(3, 245) <= input(7);
output(3, 246) <= input(8);
output(3, 247) <= input(9);
output(3, 248) <= input(10);
output(3, 249) <= input(11);
output(3, 250) <= input(12);
output(3, 251) <= input(13);
output(3, 252) <= input(14);
output(3, 253) <= input(15);
output(3, 254) <= input(34);
output(3, 255) <= input(35);
output(4, 0) <= input(19);
output(4, 1) <= input(20);
output(4, 2) <= input(21);
output(4, 3) <= input(22);
output(4, 4) <= input(23);
output(4, 5) <= input(24);
output(4, 6) <= input(25);
output(4, 7) <= input(26);
output(4, 8) <= input(27);
output(4, 9) <= input(28);
output(4, 10) <= input(29);
output(4, 11) <= input(30);
output(4, 12) <= input(31);
output(4, 13) <= input(33);
output(4, 14) <= input(36);
output(4, 15) <= input(37);
output(4, 16) <= input(19);
output(4, 17) <= input(20);
output(4, 18) <= input(21);
output(4, 19) <= input(22);
output(4, 20) <= input(23);
output(4, 21) <= input(24);
output(4, 22) <= input(25);
output(4, 23) <= input(26);
output(4, 24) <= input(27);
output(4, 25) <= input(28);
output(4, 26) <= input(29);
output(4, 27) <= input(30);
output(4, 28) <= input(31);
output(4, 29) <= input(33);
output(4, 30) <= input(36);
output(4, 31) <= input(37);
output(4, 32) <= input(19);
output(4, 33) <= input(20);
output(4, 34) <= input(21);
output(4, 35) <= input(22);
output(4, 36) <= input(23);
output(4, 37) <= input(24);
output(4, 38) <= input(25);
output(4, 39) <= input(26);
output(4, 40) <= input(27);
output(4, 41) <= input(28);
output(4, 42) <= input(29);
output(4, 43) <= input(30);
output(4, 44) <= input(31);
output(4, 45) <= input(33);
output(4, 46) <= input(36);
output(4, 47) <= input(37);
output(4, 48) <= input(19);
output(4, 49) <= input(20);
output(4, 50) <= input(21);
output(4, 51) <= input(22);
output(4, 52) <= input(23);
output(4, 53) <= input(24);
output(4, 54) <= input(25);
output(4, 55) <= input(26);
output(4, 56) <= input(27);
output(4, 57) <= input(28);
output(4, 58) <= input(29);
output(4, 59) <= input(30);
output(4, 60) <= input(31);
output(4, 61) <= input(33);
output(4, 62) <= input(36);
output(4, 63) <= input(37);
output(4, 64) <= input(19);
output(4, 65) <= input(20);
output(4, 66) <= input(21);
output(4, 67) <= input(22);
output(4, 68) <= input(23);
output(4, 69) <= input(24);
output(4, 70) <= input(25);
output(4, 71) <= input(26);
output(4, 72) <= input(27);
output(4, 73) <= input(28);
output(4, 74) <= input(29);
output(4, 75) <= input(30);
output(4, 76) <= input(31);
output(4, 77) <= input(33);
output(4, 78) <= input(36);
output(4, 79) <= input(37);
output(4, 80) <= input(19);
output(4, 81) <= input(20);
output(4, 82) <= input(21);
output(4, 83) <= input(22);
output(4, 84) <= input(23);
output(4, 85) <= input(24);
output(4, 86) <= input(25);
output(4, 87) <= input(26);
output(4, 88) <= input(27);
output(4, 89) <= input(28);
output(4, 90) <= input(29);
output(4, 91) <= input(30);
output(4, 92) <= input(31);
output(4, 93) <= input(33);
output(4, 94) <= input(36);
output(4, 95) <= input(37);
output(4, 96) <= input(19);
output(4, 97) <= input(20);
output(4, 98) <= input(21);
output(4, 99) <= input(22);
output(4, 100) <= input(23);
output(4, 101) <= input(24);
output(4, 102) <= input(25);
output(4, 103) <= input(26);
output(4, 104) <= input(27);
output(4, 105) <= input(28);
output(4, 106) <= input(29);
output(4, 107) <= input(30);
output(4, 108) <= input(31);
output(4, 109) <= input(33);
output(4, 110) <= input(36);
output(4, 111) <= input(37);
output(4, 112) <= input(19);
output(4, 113) <= input(20);
output(4, 114) <= input(21);
output(4, 115) <= input(22);
output(4, 116) <= input(23);
output(4, 117) <= input(24);
output(4, 118) <= input(25);
output(4, 119) <= input(26);
output(4, 120) <= input(27);
output(4, 121) <= input(28);
output(4, 122) <= input(29);
output(4, 123) <= input(30);
output(4, 124) <= input(31);
output(4, 125) <= input(33);
output(4, 126) <= input(36);
output(4, 127) <= input(37);
output(4, 128) <= input(19);
output(4, 129) <= input(20);
output(4, 130) <= input(21);
output(4, 131) <= input(22);
output(4, 132) <= input(23);
output(4, 133) <= input(24);
output(4, 134) <= input(25);
output(4, 135) <= input(26);
output(4, 136) <= input(27);
output(4, 137) <= input(28);
output(4, 138) <= input(29);
output(4, 139) <= input(30);
output(4, 140) <= input(31);
output(4, 141) <= input(33);
output(4, 142) <= input(36);
output(4, 143) <= input(37);
output(4, 144) <= input(19);
output(4, 145) <= input(20);
output(4, 146) <= input(21);
output(4, 147) <= input(22);
output(4, 148) <= input(23);
output(4, 149) <= input(24);
output(4, 150) <= input(25);
output(4, 151) <= input(26);
output(4, 152) <= input(27);
output(4, 153) <= input(28);
output(4, 154) <= input(29);
output(4, 155) <= input(30);
output(4, 156) <= input(31);
output(4, 157) <= input(33);
output(4, 158) <= input(36);
output(4, 159) <= input(37);
output(4, 160) <= input(19);
output(4, 161) <= input(20);
output(4, 162) <= input(21);
output(4, 163) <= input(22);
output(4, 164) <= input(23);
output(4, 165) <= input(24);
output(4, 166) <= input(25);
output(4, 167) <= input(26);
output(4, 168) <= input(27);
output(4, 169) <= input(28);
output(4, 170) <= input(29);
output(4, 171) <= input(30);
output(4, 172) <= input(31);
output(4, 173) <= input(33);
output(4, 174) <= input(36);
output(4, 175) <= input(37);
output(4, 176) <= input(19);
output(4, 177) <= input(20);
output(4, 178) <= input(21);
output(4, 179) <= input(22);
output(4, 180) <= input(23);
output(4, 181) <= input(24);
output(4, 182) <= input(25);
output(4, 183) <= input(26);
output(4, 184) <= input(27);
output(4, 185) <= input(28);
output(4, 186) <= input(29);
output(4, 187) <= input(30);
output(4, 188) <= input(31);
output(4, 189) <= input(33);
output(4, 190) <= input(36);
output(4, 191) <= input(37);
output(4, 192) <= input(19);
output(4, 193) <= input(20);
output(4, 194) <= input(21);
output(4, 195) <= input(22);
output(4, 196) <= input(23);
output(4, 197) <= input(24);
output(4, 198) <= input(25);
output(4, 199) <= input(26);
output(4, 200) <= input(27);
output(4, 201) <= input(28);
output(4, 202) <= input(29);
output(4, 203) <= input(30);
output(4, 204) <= input(31);
output(4, 205) <= input(33);
output(4, 206) <= input(36);
output(4, 207) <= input(37);
output(4, 208) <= input(19);
output(4, 209) <= input(20);
output(4, 210) <= input(21);
output(4, 211) <= input(22);
output(4, 212) <= input(23);
output(4, 213) <= input(24);
output(4, 214) <= input(25);
output(4, 215) <= input(26);
output(4, 216) <= input(27);
output(4, 217) <= input(28);
output(4, 218) <= input(29);
output(4, 219) <= input(30);
output(4, 220) <= input(31);
output(4, 221) <= input(33);
output(4, 222) <= input(36);
output(4, 223) <= input(37);
output(4, 224) <= input(19);
output(4, 225) <= input(20);
output(4, 226) <= input(21);
output(4, 227) <= input(22);
output(4, 228) <= input(23);
output(4, 229) <= input(24);
output(4, 230) <= input(25);
output(4, 231) <= input(26);
output(4, 232) <= input(27);
output(4, 233) <= input(28);
output(4, 234) <= input(29);
output(4, 235) <= input(30);
output(4, 236) <= input(31);
output(4, 237) <= input(33);
output(4, 238) <= input(36);
output(4, 239) <= input(37);
output(4, 240) <= input(3);
output(4, 241) <= input(4);
output(4, 242) <= input(5);
output(4, 243) <= input(6);
output(4, 244) <= input(7);
output(4, 245) <= input(8);
output(4, 246) <= input(9);
output(4, 247) <= input(10);
output(4, 248) <= input(11);
output(4, 249) <= input(12);
output(4, 250) <= input(13);
output(4, 251) <= input(14);
output(4, 252) <= input(15);
output(4, 253) <= input(34);
output(4, 254) <= input(35);
output(4, 255) <= input(38);
output(5, 0) <= input(3);
output(5, 1) <= input(4);
output(5, 2) <= input(5);
output(5, 3) <= input(6);
output(5, 4) <= input(7);
output(5, 5) <= input(8);
output(5, 6) <= input(9);
output(5, 7) <= input(10);
output(5, 8) <= input(11);
output(5, 9) <= input(12);
output(5, 10) <= input(13);
output(5, 11) <= input(14);
output(5, 12) <= input(15);
output(5, 13) <= input(34);
output(5, 14) <= input(35);
output(5, 15) <= input(38);
output(5, 16) <= input(3);
output(5, 17) <= input(4);
output(5, 18) <= input(5);
output(5, 19) <= input(6);
output(5, 20) <= input(7);
output(5, 21) <= input(8);
output(5, 22) <= input(9);
output(5, 23) <= input(10);
output(5, 24) <= input(11);
output(5, 25) <= input(12);
output(5, 26) <= input(13);
output(5, 27) <= input(14);
output(5, 28) <= input(15);
output(5, 29) <= input(34);
output(5, 30) <= input(35);
output(5, 31) <= input(38);
output(5, 32) <= input(3);
output(5, 33) <= input(4);
output(5, 34) <= input(5);
output(5, 35) <= input(6);
output(5, 36) <= input(7);
output(5, 37) <= input(8);
output(5, 38) <= input(9);
output(5, 39) <= input(10);
output(5, 40) <= input(11);
output(5, 41) <= input(12);
output(5, 42) <= input(13);
output(5, 43) <= input(14);
output(5, 44) <= input(15);
output(5, 45) <= input(34);
output(5, 46) <= input(35);
output(5, 47) <= input(38);
output(5, 48) <= input(3);
output(5, 49) <= input(4);
output(5, 50) <= input(5);
output(5, 51) <= input(6);
output(5, 52) <= input(7);
output(5, 53) <= input(8);
output(5, 54) <= input(9);
output(5, 55) <= input(10);
output(5, 56) <= input(11);
output(5, 57) <= input(12);
output(5, 58) <= input(13);
output(5, 59) <= input(14);
output(5, 60) <= input(15);
output(5, 61) <= input(34);
output(5, 62) <= input(35);
output(5, 63) <= input(38);
output(5, 64) <= input(3);
output(5, 65) <= input(4);
output(5, 66) <= input(5);
output(5, 67) <= input(6);
output(5, 68) <= input(7);
output(5, 69) <= input(8);
output(5, 70) <= input(9);
output(5, 71) <= input(10);
output(5, 72) <= input(11);
output(5, 73) <= input(12);
output(5, 74) <= input(13);
output(5, 75) <= input(14);
output(5, 76) <= input(15);
output(5, 77) <= input(34);
output(5, 78) <= input(35);
output(5, 79) <= input(38);
output(5, 80) <= input(3);
output(5, 81) <= input(4);
output(5, 82) <= input(5);
output(5, 83) <= input(6);
output(5, 84) <= input(7);
output(5, 85) <= input(8);
output(5, 86) <= input(9);
output(5, 87) <= input(10);
output(5, 88) <= input(11);
output(5, 89) <= input(12);
output(5, 90) <= input(13);
output(5, 91) <= input(14);
output(5, 92) <= input(15);
output(5, 93) <= input(34);
output(5, 94) <= input(35);
output(5, 95) <= input(38);
output(5, 96) <= input(3);
output(5, 97) <= input(4);
output(5, 98) <= input(5);
output(5, 99) <= input(6);
output(5, 100) <= input(7);
output(5, 101) <= input(8);
output(5, 102) <= input(9);
output(5, 103) <= input(10);
output(5, 104) <= input(11);
output(5, 105) <= input(12);
output(5, 106) <= input(13);
output(5, 107) <= input(14);
output(5, 108) <= input(15);
output(5, 109) <= input(34);
output(5, 110) <= input(35);
output(5, 111) <= input(38);
output(5, 112) <= input(20);
output(5, 113) <= input(21);
output(5, 114) <= input(22);
output(5, 115) <= input(23);
output(5, 116) <= input(24);
output(5, 117) <= input(25);
output(5, 118) <= input(26);
output(5, 119) <= input(27);
output(5, 120) <= input(28);
output(5, 121) <= input(29);
output(5, 122) <= input(30);
output(5, 123) <= input(31);
output(5, 124) <= input(33);
output(5, 125) <= input(36);
output(5, 126) <= input(37);
output(5, 127) <= input(39);
output(5, 128) <= input(20);
output(5, 129) <= input(21);
output(5, 130) <= input(22);
output(5, 131) <= input(23);
output(5, 132) <= input(24);
output(5, 133) <= input(25);
output(5, 134) <= input(26);
output(5, 135) <= input(27);
output(5, 136) <= input(28);
output(5, 137) <= input(29);
output(5, 138) <= input(30);
output(5, 139) <= input(31);
output(5, 140) <= input(33);
output(5, 141) <= input(36);
output(5, 142) <= input(37);
output(5, 143) <= input(39);
output(5, 144) <= input(20);
output(5, 145) <= input(21);
output(5, 146) <= input(22);
output(5, 147) <= input(23);
output(5, 148) <= input(24);
output(5, 149) <= input(25);
output(5, 150) <= input(26);
output(5, 151) <= input(27);
output(5, 152) <= input(28);
output(5, 153) <= input(29);
output(5, 154) <= input(30);
output(5, 155) <= input(31);
output(5, 156) <= input(33);
output(5, 157) <= input(36);
output(5, 158) <= input(37);
output(5, 159) <= input(39);
output(5, 160) <= input(20);
output(5, 161) <= input(21);
output(5, 162) <= input(22);
output(5, 163) <= input(23);
output(5, 164) <= input(24);
output(5, 165) <= input(25);
output(5, 166) <= input(26);
output(5, 167) <= input(27);
output(5, 168) <= input(28);
output(5, 169) <= input(29);
output(5, 170) <= input(30);
output(5, 171) <= input(31);
output(5, 172) <= input(33);
output(5, 173) <= input(36);
output(5, 174) <= input(37);
output(5, 175) <= input(39);
output(5, 176) <= input(20);
output(5, 177) <= input(21);
output(5, 178) <= input(22);
output(5, 179) <= input(23);
output(5, 180) <= input(24);
output(5, 181) <= input(25);
output(5, 182) <= input(26);
output(5, 183) <= input(27);
output(5, 184) <= input(28);
output(5, 185) <= input(29);
output(5, 186) <= input(30);
output(5, 187) <= input(31);
output(5, 188) <= input(33);
output(5, 189) <= input(36);
output(5, 190) <= input(37);
output(5, 191) <= input(39);
output(5, 192) <= input(20);
output(5, 193) <= input(21);
output(5, 194) <= input(22);
output(5, 195) <= input(23);
output(5, 196) <= input(24);
output(5, 197) <= input(25);
output(5, 198) <= input(26);
output(5, 199) <= input(27);
output(5, 200) <= input(28);
output(5, 201) <= input(29);
output(5, 202) <= input(30);
output(5, 203) <= input(31);
output(5, 204) <= input(33);
output(5, 205) <= input(36);
output(5, 206) <= input(37);
output(5, 207) <= input(39);
output(5, 208) <= input(20);
output(5, 209) <= input(21);
output(5, 210) <= input(22);
output(5, 211) <= input(23);
output(5, 212) <= input(24);
output(5, 213) <= input(25);
output(5, 214) <= input(26);
output(5, 215) <= input(27);
output(5, 216) <= input(28);
output(5, 217) <= input(29);
output(5, 218) <= input(30);
output(5, 219) <= input(31);
output(5, 220) <= input(33);
output(5, 221) <= input(36);
output(5, 222) <= input(37);
output(5, 223) <= input(39);
output(5, 224) <= input(20);
output(5, 225) <= input(21);
output(5, 226) <= input(22);
output(5, 227) <= input(23);
output(5, 228) <= input(24);
output(5, 229) <= input(25);
output(5, 230) <= input(26);
output(5, 231) <= input(27);
output(5, 232) <= input(28);
output(5, 233) <= input(29);
output(5, 234) <= input(30);
output(5, 235) <= input(31);
output(5, 236) <= input(33);
output(5, 237) <= input(36);
output(5, 238) <= input(37);
output(5, 239) <= input(39);
output(5, 240) <= input(4);
output(5, 241) <= input(5);
output(5, 242) <= input(6);
output(5, 243) <= input(7);
output(5, 244) <= input(8);
output(5, 245) <= input(9);
output(5, 246) <= input(10);
output(5, 247) <= input(11);
output(5, 248) <= input(12);
output(5, 249) <= input(13);
output(5, 250) <= input(14);
output(5, 251) <= input(15);
output(5, 252) <= input(34);
output(5, 253) <= input(35);
output(5, 254) <= input(38);
output(5, 255) <= input(40);
output(6, 0) <= input(20);
output(6, 1) <= input(21);
output(6, 2) <= input(22);
output(6, 3) <= input(23);
output(6, 4) <= input(24);
output(6, 5) <= input(25);
output(6, 6) <= input(26);
output(6, 7) <= input(27);
output(6, 8) <= input(28);
output(6, 9) <= input(29);
output(6, 10) <= input(30);
output(6, 11) <= input(31);
output(6, 12) <= input(33);
output(6, 13) <= input(36);
output(6, 14) <= input(37);
output(6, 15) <= input(39);
output(6, 16) <= input(20);
output(6, 17) <= input(21);
output(6, 18) <= input(22);
output(6, 19) <= input(23);
output(6, 20) <= input(24);
output(6, 21) <= input(25);
output(6, 22) <= input(26);
output(6, 23) <= input(27);
output(6, 24) <= input(28);
output(6, 25) <= input(29);
output(6, 26) <= input(30);
output(6, 27) <= input(31);
output(6, 28) <= input(33);
output(6, 29) <= input(36);
output(6, 30) <= input(37);
output(6, 31) <= input(39);
output(6, 32) <= input(20);
output(6, 33) <= input(21);
output(6, 34) <= input(22);
output(6, 35) <= input(23);
output(6, 36) <= input(24);
output(6, 37) <= input(25);
output(6, 38) <= input(26);
output(6, 39) <= input(27);
output(6, 40) <= input(28);
output(6, 41) <= input(29);
output(6, 42) <= input(30);
output(6, 43) <= input(31);
output(6, 44) <= input(33);
output(6, 45) <= input(36);
output(6, 46) <= input(37);
output(6, 47) <= input(39);
output(6, 48) <= input(20);
output(6, 49) <= input(21);
output(6, 50) <= input(22);
output(6, 51) <= input(23);
output(6, 52) <= input(24);
output(6, 53) <= input(25);
output(6, 54) <= input(26);
output(6, 55) <= input(27);
output(6, 56) <= input(28);
output(6, 57) <= input(29);
output(6, 58) <= input(30);
output(6, 59) <= input(31);
output(6, 60) <= input(33);
output(6, 61) <= input(36);
output(6, 62) <= input(37);
output(6, 63) <= input(39);
output(6, 64) <= input(20);
output(6, 65) <= input(21);
output(6, 66) <= input(22);
output(6, 67) <= input(23);
output(6, 68) <= input(24);
output(6, 69) <= input(25);
output(6, 70) <= input(26);
output(6, 71) <= input(27);
output(6, 72) <= input(28);
output(6, 73) <= input(29);
output(6, 74) <= input(30);
output(6, 75) <= input(31);
output(6, 76) <= input(33);
output(6, 77) <= input(36);
output(6, 78) <= input(37);
output(6, 79) <= input(39);
output(6, 80) <= input(4);
output(6, 81) <= input(5);
output(6, 82) <= input(6);
output(6, 83) <= input(7);
output(6, 84) <= input(8);
output(6, 85) <= input(9);
output(6, 86) <= input(10);
output(6, 87) <= input(11);
output(6, 88) <= input(12);
output(6, 89) <= input(13);
output(6, 90) <= input(14);
output(6, 91) <= input(15);
output(6, 92) <= input(34);
output(6, 93) <= input(35);
output(6, 94) <= input(38);
output(6, 95) <= input(40);
output(6, 96) <= input(4);
output(6, 97) <= input(5);
output(6, 98) <= input(6);
output(6, 99) <= input(7);
output(6, 100) <= input(8);
output(6, 101) <= input(9);
output(6, 102) <= input(10);
output(6, 103) <= input(11);
output(6, 104) <= input(12);
output(6, 105) <= input(13);
output(6, 106) <= input(14);
output(6, 107) <= input(15);
output(6, 108) <= input(34);
output(6, 109) <= input(35);
output(6, 110) <= input(38);
output(6, 111) <= input(40);
output(6, 112) <= input(4);
output(6, 113) <= input(5);
output(6, 114) <= input(6);
output(6, 115) <= input(7);
output(6, 116) <= input(8);
output(6, 117) <= input(9);
output(6, 118) <= input(10);
output(6, 119) <= input(11);
output(6, 120) <= input(12);
output(6, 121) <= input(13);
output(6, 122) <= input(14);
output(6, 123) <= input(15);
output(6, 124) <= input(34);
output(6, 125) <= input(35);
output(6, 126) <= input(38);
output(6, 127) <= input(40);
output(6, 128) <= input(4);
output(6, 129) <= input(5);
output(6, 130) <= input(6);
output(6, 131) <= input(7);
output(6, 132) <= input(8);
output(6, 133) <= input(9);
output(6, 134) <= input(10);
output(6, 135) <= input(11);
output(6, 136) <= input(12);
output(6, 137) <= input(13);
output(6, 138) <= input(14);
output(6, 139) <= input(15);
output(6, 140) <= input(34);
output(6, 141) <= input(35);
output(6, 142) <= input(38);
output(6, 143) <= input(40);
output(6, 144) <= input(4);
output(6, 145) <= input(5);
output(6, 146) <= input(6);
output(6, 147) <= input(7);
output(6, 148) <= input(8);
output(6, 149) <= input(9);
output(6, 150) <= input(10);
output(6, 151) <= input(11);
output(6, 152) <= input(12);
output(6, 153) <= input(13);
output(6, 154) <= input(14);
output(6, 155) <= input(15);
output(6, 156) <= input(34);
output(6, 157) <= input(35);
output(6, 158) <= input(38);
output(6, 159) <= input(40);
output(6, 160) <= input(21);
output(6, 161) <= input(22);
output(6, 162) <= input(23);
output(6, 163) <= input(24);
output(6, 164) <= input(25);
output(6, 165) <= input(26);
output(6, 166) <= input(27);
output(6, 167) <= input(28);
output(6, 168) <= input(29);
output(6, 169) <= input(30);
output(6, 170) <= input(31);
output(6, 171) <= input(33);
output(6, 172) <= input(36);
output(6, 173) <= input(37);
output(6, 174) <= input(39);
output(6, 175) <= input(41);
output(6, 176) <= input(21);
output(6, 177) <= input(22);
output(6, 178) <= input(23);
output(6, 179) <= input(24);
output(6, 180) <= input(25);
output(6, 181) <= input(26);
output(6, 182) <= input(27);
output(6, 183) <= input(28);
output(6, 184) <= input(29);
output(6, 185) <= input(30);
output(6, 186) <= input(31);
output(6, 187) <= input(33);
output(6, 188) <= input(36);
output(6, 189) <= input(37);
output(6, 190) <= input(39);
output(6, 191) <= input(41);
output(6, 192) <= input(21);
output(6, 193) <= input(22);
output(6, 194) <= input(23);
output(6, 195) <= input(24);
output(6, 196) <= input(25);
output(6, 197) <= input(26);
output(6, 198) <= input(27);
output(6, 199) <= input(28);
output(6, 200) <= input(29);
output(6, 201) <= input(30);
output(6, 202) <= input(31);
output(6, 203) <= input(33);
output(6, 204) <= input(36);
output(6, 205) <= input(37);
output(6, 206) <= input(39);
output(6, 207) <= input(41);
output(6, 208) <= input(21);
output(6, 209) <= input(22);
output(6, 210) <= input(23);
output(6, 211) <= input(24);
output(6, 212) <= input(25);
output(6, 213) <= input(26);
output(6, 214) <= input(27);
output(6, 215) <= input(28);
output(6, 216) <= input(29);
output(6, 217) <= input(30);
output(6, 218) <= input(31);
output(6, 219) <= input(33);
output(6, 220) <= input(36);
output(6, 221) <= input(37);
output(6, 222) <= input(39);
output(6, 223) <= input(41);
output(6, 224) <= input(21);
output(6, 225) <= input(22);
output(6, 226) <= input(23);
output(6, 227) <= input(24);
output(6, 228) <= input(25);
output(6, 229) <= input(26);
output(6, 230) <= input(27);
output(6, 231) <= input(28);
output(6, 232) <= input(29);
output(6, 233) <= input(30);
output(6, 234) <= input(31);
output(6, 235) <= input(33);
output(6, 236) <= input(36);
output(6, 237) <= input(37);
output(6, 238) <= input(39);
output(6, 239) <= input(41);
output(6, 240) <= input(5);
output(6, 241) <= input(6);
output(6, 242) <= input(7);
output(6, 243) <= input(8);
output(6, 244) <= input(9);
output(6, 245) <= input(10);
output(6, 246) <= input(11);
output(6, 247) <= input(12);
output(6, 248) <= input(13);
output(6, 249) <= input(14);
output(6, 250) <= input(15);
output(6, 251) <= input(34);
output(6, 252) <= input(35);
output(6, 253) <= input(38);
output(6, 254) <= input(40);
output(6, 255) <= input(42);
output(7, 0) <= input(4);
output(7, 1) <= input(5);
output(7, 2) <= input(6);
output(7, 3) <= input(7);
output(7, 4) <= input(8);
output(7, 5) <= input(9);
output(7, 6) <= input(10);
output(7, 7) <= input(11);
output(7, 8) <= input(12);
output(7, 9) <= input(13);
output(7, 10) <= input(14);
output(7, 11) <= input(15);
output(7, 12) <= input(34);
output(7, 13) <= input(35);
output(7, 14) <= input(38);
output(7, 15) <= input(40);
output(7, 16) <= input(4);
output(7, 17) <= input(5);
output(7, 18) <= input(6);
output(7, 19) <= input(7);
output(7, 20) <= input(8);
output(7, 21) <= input(9);
output(7, 22) <= input(10);
output(7, 23) <= input(11);
output(7, 24) <= input(12);
output(7, 25) <= input(13);
output(7, 26) <= input(14);
output(7, 27) <= input(15);
output(7, 28) <= input(34);
output(7, 29) <= input(35);
output(7, 30) <= input(38);
output(7, 31) <= input(40);
output(7, 32) <= input(4);
output(7, 33) <= input(5);
output(7, 34) <= input(6);
output(7, 35) <= input(7);
output(7, 36) <= input(8);
output(7, 37) <= input(9);
output(7, 38) <= input(10);
output(7, 39) <= input(11);
output(7, 40) <= input(12);
output(7, 41) <= input(13);
output(7, 42) <= input(14);
output(7, 43) <= input(15);
output(7, 44) <= input(34);
output(7, 45) <= input(35);
output(7, 46) <= input(38);
output(7, 47) <= input(40);
output(7, 48) <= input(21);
output(7, 49) <= input(22);
output(7, 50) <= input(23);
output(7, 51) <= input(24);
output(7, 52) <= input(25);
output(7, 53) <= input(26);
output(7, 54) <= input(27);
output(7, 55) <= input(28);
output(7, 56) <= input(29);
output(7, 57) <= input(30);
output(7, 58) <= input(31);
output(7, 59) <= input(33);
output(7, 60) <= input(36);
output(7, 61) <= input(37);
output(7, 62) <= input(39);
output(7, 63) <= input(41);
output(7, 64) <= input(21);
output(7, 65) <= input(22);
output(7, 66) <= input(23);
output(7, 67) <= input(24);
output(7, 68) <= input(25);
output(7, 69) <= input(26);
output(7, 70) <= input(27);
output(7, 71) <= input(28);
output(7, 72) <= input(29);
output(7, 73) <= input(30);
output(7, 74) <= input(31);
output(7, 75) <= input(33);
output(7, 76) <= input(36);
output(7, 77) <= input(37);
output(7, 78) <= input(39);
output(7, 79) <= input(41);
output(7, 80) <= input(21);
output(7, 81) <= input(22);
output(7, 82) <= input(23);
output(7, 83) <= input(24);
output(7, 84) <= input(25);
output(7, 85) <= input(26);
output(7, 86) <= input(27);
output(7, 87) <= input(28);
output(7, 88) <= input(29);
output(7, 89) <= input(30);
output(7, 90) <= input(31);
output(7, 91) <= input(33);
output(7, 92) <= input(36);
output(7, 93) <= input(37);
output(7, 94) <= input(39);
output(7, 95) <= input(41);
output(7, 96) <= input(21);
output(7, 97) <= input(22);
output(7, 98) <= input(23);
output(7, 99) <= input(24);
output(7, 100) <= input(25);
output(7, 101) <= input(26);
output(7, 102) <= input(27);
output(7, 103) <= input(28);
output(7, 104) <= input(29);
output(7, 105) <= input(30);
output(7, 106) <= input(31);
output(7, 107) <= input(33);
output(7, 108) <= input(36);
output(7, 109) <= input(37);
output(7, 110) <= input(39);
output(7, 111) <= input(41);
output(7, 112) <= input(5);
output(7, 113) <= input(6);
output(7, 114) <= input(7);
output(7, 115) <= input(8);
output(7, 116) <= input(9);
output(7, 117) <= input(10);
output(7, 118) <= input(11);
output(7, 119) <= input(12);
output(7, 120) <= input(13);
output(7, 121) <= input(14);
output(7, 122) <= input(15);
output(7, 123) <= input(34);
output(7, 124) <= input(35);
output(7, 125) <= input(38);
output(7, 126) <= input(40);
output(7, 127) <= input(42);
output(7, 128) <= input(5);
output(7, 129) <= input(6);
output(7, 130) <= input(7);
output(7, 131) <= input(8);
output(7, 132) <= input(9);
output(7, 133) <= input(10);
output(7, 134) <= input(11);
output(7, 135) <= input(12);
output(7, 136) <= input(13);
output(7, 137) <= input(14);
output(7, 138) <= input(15);
output(7, 139) <= input(34);
output(7, 140) <= input(35);
output(7, 141) <= input(38);
output(7, 142) <= input(40);
output(7, 143) <= input(42);
output(7, 144) <= input(5);
output(7, 145) <= input(6);
output(7, 146) <= input(7);
output(7, 147) <= input(8);
output(7, 148) <= input(9);
output(7, 149) <= input(10);
output(7, 150) <= input(11);
output(7, 151) <= input(12);
output(7, 152) <= input(13);
output(7, 153) <= input(14);
output(7, 154) <= input(15);
output(7, 155) <= input(34);
output(7, 156) <= input(35);
output(7, 157) <= input(38);
output(7, 158) <= input(40);
output(7, 159) <= input(42);
output(7, 160) <= input(5);
output(7, 161) <= input(6);
output(7, 162) <= input(7);
output(7, 163) <= input(8);
output(7, 164) <= input(9);
output(7, 165) <= input(10);
output(7, 166) <= input(11);
output(7, 167) <= input(12);
output(7, 168) <= input(13);
output(7, 169) <= input(14);
output(7, 170) <= input(15);
output(7, 171) <= input(34);
output(7, 172) <= input(35);
output(7, 173) <= input(38);
output(7, 174) <= input(40);
output(7, 175) <= input(42);
output(7, 176) <= input(22);
output(7, 177) <= input(23);
output(7, 178) <= input(24);
output(7, 179) <= input(25);
output(7, 180) <= input(26);
output(7, 181) <= input(27);
output(7, 182) <= input(28);
output(7, 183) <= input(29);
output(7, 184) <= input(30);
output(7, 185) <= input(31);
output(7, 186) <= input(33);
output(7, 187) <= input(36);
output(7, 188) <= input(37);
output(7, 189) <= input(39);
output(7, 190) <= input(41);
output(7, 191) <= input(43);
output(7, 192) <= input(22);
output(7, 193) <= input(23);
output(7, 194) <= input(24);
output(7, 195) <= input(25);
output(7, 196) <= input(26);
output(7, 197) <= input(27);
output(7, 198) <= input(28);
output(7, 199) <= input(29);
output(7, 200) <= input(30);
output(7, 201) <= input(31);
output(7, 202) <= input(33);
output(7, 203) <= input(36);
output(7, 204) <= input(37);
output(7, 205) <= input(39);
output(7, 206) <= input(41);
output(7, 207) <= input(43);
output(7, 208) <= input(22);
output(7, 209) <= input(23);
output(7, 210) <= input(24);
output(7, 211) <= input(25);
output(7, 212) <= input(26);
output(7, 213) <= input(27);
output(7, 214) <= input(28);
output(7, 215) <= input(29);
output(7, 216) <= input(30);
output(7, 217) <= input(31);
output(7, 218) <= input(33);
output(7, 219) <= input(36);
output(7, 220) <= input(37);
output(7, 221) <= input(39);
output(7, 222) <= input(41);
output(7, 223) <= input(43);
output(7, 224) <= input(22);
output(7, 225) <= input(23);
output(7, 226) <= input(24);
output(7, 227) <= input(25);
output(7, 228) <= input(26);
output(7, 229) <= input(27);
output(7, 230) <= input(28);
output(7, 231) <= input(29);
output(7, 232) <= input(30);
output(7, 233) <= input(31);
output(7, 234) <= input(33);
output(7, 235) <= input(36);
output(7, 236) <= input(37);
output(7, 237) <= input(39);
output(7, 238) <= input(41);
output(7, 239) <= input(43);
output(7, 240) <= input(6);
output(7, 241) <= input(7);
output(7, 242) <= input(8);
output(7, 243) <= input(9);
output(7, 244) <= input(10);
output(7, 245) <= input(11);
output(7, 246) <= input(12);
output(7, 247) <= input(13);
output(7, 248) <= input(14);
output(7, 249) <= input(15);
output(7, 250) <= input(34);
output(7, 251) <= input(35);
output(7, 252) <= input(38);
output(7, 253) <= input(40);
output(7, 254) <= input(42);
output(7, 255) <= input(44);
when "1110" =>
output(0, 0) <= input(0);
output(0, 1) <= input(1);
output(0, 2) <= input(2);
output(0, 3) <= input(3);
output(0, 4) <= input(4);
output(0, 5) <= input(5);
output(0, 6) <= input(6);
output(0, 7) <= input(7);
output(0, 8) <= input(8);
output(0, 9) <= input(9);
output(0, 10) <= input(10);
output(0, 11) <= input(11);
output(0, 12) <= input(12);
output(0, 13) <= input(13);
output(0, 14) <= input(14);
output(0, 15) <= input(15);
output(0, 16) <= input(0);
output(0, 17) <= input(1);
output(0, 18) <= input(2);
output(0, 19) <= input(3);
output(0, 20) <= input(4);
output(0, 21) <= input(5);
output(0, 22) <= input(6);
output(0, 23) <= input(7);
output(0, 24) <= input(8);
output(0, 25) <= input(9);
output(0, 26) <= input(10);
output(0, 27) <= input(11);
output(0, 28) <= input(12);
output(0, 29) <= input(13);
output(0, 30) <= input(14);
output(0, 31) <= input(15);
output(0, 32) <= input(16);
output(0, 33) <= input(17);
output(0, 34) <= input(18);
output(0, 35) <= input(19);
output(0, 36) <= input(20);
output(0, 37) <= input(21);
output(0, 38) <= input(22);
output(0, 39) <= input(23);
output(0, 40) <= input(24);
output(0, 41) <= input(25);
output(0, 42) <= input(26);
output(0, 43) <= input(27);
output(0, 44) <= input(28);
output(0, 45) <= input(29);
output(0, 46) <= input(30);
output(0, 47) <= input(31);
output(0, 48) <= input(16);
output(0, 49) <= input(17);
output(0, 50) <= input(18);
output(0, 51) <= input(19);
output(0, 52) <= input(20);
output(0, 53) <= input(21);
output(0, 54) <= input(22);
output(0, 55) <= input(23);
output(0, 56) <= input(24);
output(0, 57) <= input(25);
output(0, 58) <= input(26);
output(0, 59) <= input(27);
output(0, 60) <= input(28);
output(0, 61) <= input(29);
output(0, 62) <= input(30);
output(0, 63) <= input(31);
output(0, 64) <= input(16);
output(0, 65) <= input(17);
output(0, 66) <= input(18);
output(0, 67) <= input(19);
output(0, 68) <= input(20);
output(0, 69) <= input(21);
output(0, 70) <= input(22);
output(0, 71) <= input(23);
output(0, 72) <= input(24);
output(0, 73) <= input(25);
output(0, 74) <= input(26);
output(0, 75) <= input(27);
output(0, 76) <= input(28);
output(0, 77) <= input(29);
output(0, 78) <= input(30);
output(0, 79) <= input(31);
output(0, 80) <= input(1);
output(0, 81) <= input(2);
output(0, 82) <= input(3);
output(0, 83) <= input(4);
output(0, 84) <= input(5);
output(0, 85) <= input(6);
output(0, 86) <= input(7);
output(0, 87) <= input(8);
output(0, 88) <= input(9);
output(0, 89) <= input(10);
output(0, 90) <= input(11);
output(0, 91) <= input(12);
output(0, 92) <= input(13);
output(0, 93) <= input(14);
output(0, 94) <= input(15);
output(0, 95) <= input(32);
output(0, 96) <= input(1);
output(0, 97) <= input(2);
output(0, 98) <= input(3);
output(0, 99) <= input(4);
output(0, 100) <= input(5);
output(0, 101) <= input(6);
output(0, 102) <= input(7);
output(0, 103) <= input(8);
output(0, 104) <= input(9);
output(0, 105) <= input(10);
output(0, 106) <= input(11);
output(0, 107) <= input(12);
output(0, 108) <= input(13);
output(0, 109) <= input(14);
output(0, 110) <= input(15);
output(0, 111) <= input(32);
output(0, 112) <= input(17);
output(0, 113) <= input(18);
output(0, 114) <= input(19);
output(0, 115) <= input(20);
output(0, 116) <= input(21);
output(0, 117) <= input(22);
output(0, 118) <= input(23);
output(0, 119) <= input(24);
output(0, 120) <= input(25);
output(0, 121) <= input(26);
output(0, 122) <= input(27);
output(0, 123) <= input(28);
output(0, 124) <= input(29);
output(0, 125) <= input(30);
output(0, 126) <= input(31);
output(0, 127) <= input(33);
output(0, 128) <= input(17);
output(0, 129) <= input(18);
output(0, 130) <= input(19);
output(0, 131) <= input(20);
output(0, 132) <= input(21);
output(0, 133) <= input(22);
output(0, 134) <= input(23);
output(0, 135) <= input(24);
output(0, 136) <= input(25);
output(0, 137) <= input(26);
output(0, 138) <= input(27);
output(0, 139) <= input(28);
output(0, 140) <= input(29);
output(0, 141) <= input(30);
output(0, 142) <= input(31);
output(0, 143) <= input(33);
output(0, 144) <= input(17);
output(0, 145) <= input(18);
output(0, 146) <= input(19);
output(0, 147) <= input(20);
output(0, 148) <= input(21);
output(0, 149) <= input(22);
output(0, 150) <= input(23);
output(0, 151) <= input(24);
output(0, 152) <= input(25);
output(0, 153) <= input(26);
output(0, 154) <= input(27);
output(0, 155) <= input(28);
output(0, 156) <= input(29);
output(0, 157) <= input(30);
output(0, 158) <= input(31);
output(0, 159) <= input(33);
output(0, 160) <= input(2);
output(0, 161) <= input(3);
output(0, 162) <= input(4);
output(0, 163) <= input(5);
output(0, 164) <= input(6);
output(0, 165) <= input(7);
output(0, 166) <= input(8);
output(0, 167) <= input(9);
output(0, 168) <= input(10);
output(0, 169) <= input(11);
output(0, 170) <= input(12);
output(0, 171) <= input(13);
output(0, 172) <= input(14);
output(0, 173) <= input(15);
output(0, 174) <= input(32);
output(0, 175) <= input(34);
output(0, 176) <= input(2);
output(0, 177) <= input(3);
output(0, 178) <= input(4);
output(0, 179) <= input(5);
output(0, 180) <= input(6);
output(0, 181) <= input(7);
output(0, 182) <= input(8);
output(0, 183) <= input(9);
output(0, 184) <= input(10);
output(0, 185) <= input(11);
output(0, 186) <= input(12);
output(0, 187) <= input(13);
output(0, 188) <= input(14);
output(0, 189) <= input(15);
output(0, 190) <= input(32);
output(0, 191) <= input(34);
output(0, 192) <= input(2);
output(0, 193) <= input(3);
output(0, 194) <= input(4);
output(0, 195) <= input(5);
output(0, 196) <= input(6);
output(0, 197) <= input(7);
output(0, 198) <= input(8);
output(0, 199) <= input(9);
output(0, 200) <= input(10);
output(0, 201) <= input(11);
output(0, 202) <= input(12);
output(0, 203) <= input(13);
output(0, 204) <= input(14);
output(0, 205) <= input(15);
output(0, 206) <= input(32);
output(0, 207) <= input(34);
output(0, 208) <= input(18);
output(0, 209) <= input(19);
output(0, 210) <= input(20);
output(0, 211) <= input(21);
output(0, 212) <= input(22);
output(0, 213) <= input(23);
output(0, 214) <= input(24);
output(0, 215) <= input(25);
output(0, 216) <= input(26);
output(0, 217) <= input(27);
output(0, 218) <= input(28);
output(0, 219) <= input(29);
output(0, 220) <= input(30);
output(0, 221) <= input(31);
output(0, 222) <= input(33);
output(0, 223) <= input(35);
output(0, 224) <= input(18);
output(0, 225) <= input(19);
output(0, 226) <= input(20);
output(0, 227) <= input(21);
output(0, 228) <= input(22);
output(0, 229) <= input(23);
output(0, 230) <= input(24);
output(0, 231) <= input(25);
output(0, 232) <= input(26);
output(0, 233) <= input(27);
output(0, 234) <= input(28);
output(0, 235) <= input(29);
output(0, 236) <= input(30);
output(0, 237) <= input(31);
output(0, 238) <= input(33);
output(0, 239) <= input(35);
output(0, 240) <= input(3);
output(0, 241) <= input(4);
output(0, 242) <= input(5);
output(0, 243) <= input(6);
output(0, 244) <= input(7);
output(0, 245) <= input(8);
output(0, 246) <= input(9);
output(0, 247) <= input(10);
output(0, 248) <= input(11);
output(0, 249) <= input(12);
output(0, 250) <= input(13);
output(0, 251) <= input(14);
output(0, 252) <= input(15);
output(0, 253) <= input(32);
output(0, 254) <= input(34);
output(0, 255) <= input(36);
output(1, 0) <= input(1);
output(1, 1) <= input(2);
output(1, 2) <= input(3);
output(1, 3) <= input(4);
output(1, 4) <= input(5);
output(1, 5) <= input(6);
output(1, 6) <= input(7);
output(1, 7) <= input(8);
output(1, 8) <= input(9);
output(1, 9) <= input(10);
output(1, 10) <= input(11);
output(1, 11) <= input(12);
output(1, 12) <= input(13);
output(1, 13) <= input(14);
output(1, 14) <= input(15);
output(1, 15) <= input(32);
output(1, 16) <= input(17);
output(1, 17) <= input(18);
output(1, 18) <= input(19);
output(1, 19) <= input(20);
output(1, 20) <= input(21);
output(1, 21) <= input(22);
output(1, 22) <= input(23);
output(1, 23) <= input(24);
output(1, 24) <= input(25);
output(1, 25) <= input(26);
output(1, 26) <= input(27);
output(1, 27) <= input(28);
output(1, 28) <= input(29);
output(1, 29) <= input(30);
output(1, 30) <= input(31);
output(1, 31) <= input(33);
output(1, 32) <= input(17);
output(1, 33) <= input(18);
output(1, 34) <= input(19);
output(1, 35) <= input(20);
output(1, 36) <= input(21);
output(1, 37) <= input(22);
output(1, 38) <= input(23);
output(1, 39) <= input(24);
output(1, 40) <= input(25);
output(1, 41) <= input(26);
output(1, 42) <= input(27);
output(1, 43) <= input(28);
output(1, 44) <= input(29);
output(1, 45) <= input(30);
output(1, 46) <= input(31);
output(1, 47) <= input(33);
output(1, 48) <= input(2);
output(1, 49) <= input(3);
output(1, 50) <= input(4);
output(1, 51) <= input(5);
output(1, 52) <= input(6);
output(1, 53) <= input(7);
output(1, 54) <= input(8);
output(1, 55) <= input(9);
output(1, 56) <= input(10);
output(1, 57) <= input(11);
output(1, 58) <= input(12);
output(1, 59) <= input(13);
output(1, 60) <= input(14);
output(1, 61) <= input(15);
output(1, 62) <= input(32);
output(1, 63) <= input(34);
output(1, 64) <= input(2);
output(1, 65) <= input(3);
output(1, 66) <= input(4);
output(1, 67) <= input(5);
output(1, 68) <= input(6);
output(1, 69) <= input(7);
output(1, 70) <= input(8);
output(1, 71) <= input(9);
output(1, 72) <= input(10);
output(1, 73) <= input(11);
output(1, 74) <= input(12);
output(1, 75) <= input(13);
output(1, 76) <= input(14);
output(1, 77) <= input(15);
output(1, 78) <= input(32);
output(1, 79) <= input(34);
output(1, 80) <= input(18);
output(1, 81) <= input(19);
output(1, 82) <= input(20);
output(1, 83) <= input(21);
output(1, 84) <= input(22);
output(1, 85) <= input(23);
output(1, 86) <= input(24);
output(1, 87) <= input(25);
output(1, 88) <= input(26);
output(1, 89) <= input(27);
output(1, 90) <= input(28);
output(1, 91) <= input(29);
output(1, 92) <= input(30);
output(1, 93) <= input(31);
output(1, 94) <= input(33);
output(1, 95) <= input(35);
output(1, 96) <= input(18);
output(1, 97) <= input(19);
output(1, 98) <= input(20);
output(1, 99) <= input(21);
output(1, 100) <= input(22);
output(1, 101) <= input(23);
output(1, 102) <= input(24);
output(1, 103) <= input(25);
output(1, 104) <= input(26);
output(1, 105) <= input(27);
output(1, 106) <= input(28);
output(1, 107) <= input(29);
output(1, 108) <= input(30);
output(1, 109) <= input(31);
output(1, 110) <= input(33);
output(1, 111) <= input(35);
output(1, 112) <= input(3);
output(1, 113) <= input(4);
output(1, 114) <= input(5);
output(1, 115) <= input(6);
output(1, 116) <= input(7);
output(1, 117) <= input(8);
output(1, 118) <= input(9);
output(1, 119) <= input(10);
output(1, 120) <= input(11);
output(1, 121) <= input(12);
output(1, 122) <= input(13);
output(1, 123) <= input(14);
output(1, 124) <= input(15);
output(1, 125) <= input(32);
output(1, 126) <= input(34);
output(1, 127) <= input(36);
output(1, 128) <= input(3);
output(1, 129) <= input(4);
output(1, 130) <= input(5);
output(1, 131) <= input(6);
output(1, 132) <= input(7);
output(1, 133) <= input(8);
output(1, 134) <= input(9);
output(1, 135) <= input(10);
output(1, 136) <= input(11);
output(1, 137) <= input(12);
output(1, 138) <= input(13);
output(1, 139) <= input(14);
output(1, 140) <= input(15);
output(1, 141) <= input(32);
output(1, 142) <= input(34);
output(1, 143) <= input(36);
output(1, 144) <= input(19);
output(1, 145) <= input(20);
output(1, 146) <= input(21);
output(1, 147) <= input(22);
output(1, 148) <= input(23);
output(1, 149) <= input(24);
output(1, 150) <= input(25);
output(1, 151) <= input(26);
output(1, 152) <= input(27);
output(1, 153) <= input(28);
output(1, 154) <= input(29);
output(1, 155) <= input(30);
output(1, 156) <= input(31);
output(1, 157) <= input(33);
output(1, 158) <= input(35);
output(1, 159) <= input(37);
output(1, 160) <= input(19);
output(1, 161) <= input(20);
output(1, 162) <= input(21);
output(1, 163) <= input(22);
output(1, 164) <= input(23);
output(1, 165) <= input(24);
output(1, 166) <= input(25);
output(1, 167) <= input(26);
output(1, 168) <= input(27);
output(1, 169) <= input(28);
output(1, 170) <= input(29);
output(1, 171) <= input(30);
output(1, 172) <= input(31);
output(1, 173) <= input(33);
output(1, 174) <= input(35);
output(1, 175) <= input(37);
output(1, 176) <= input(4);
output(1, 177) <= input(5);
output(1, 178) <= input(6);
output(1, 179) <= input(7);
output(1, 180) <= input(8);
output(1, 181) <= input(9);
output(1, 182) <= input(10);
output(1, 183) <= input(11);
output(1, 184) <= input(12);
output(1, 185) <= input(13);
output(1, 186) <= input(14);
output(1, 187) <= input(15);
output(1, 188) <= input(32);
output(1, 189) <= input(34);
output(1, 190) <= input(36);
output(1, 191) <= input(38);
output(1, 192) <= input(4);
output(1, 193) <= input(5);
output(1, 194) <= input(6);
output(1, 195) <= input(7);
output(1, 196) <= input(8);
output(1, 197) <= input(9);
output(1, 198) <= input(10);
output(1, 199) <= input(11);
output(1, 200) <= input(12);
output(1, 201) <= input(13);
output(1, 202) <= input(14);
output(1, 203) <= input(15);
output(1, 204) <= input(32);
output(1, 205) <= input(34);
output(1, 206) <= input(36);
output(1, 207) <= input(38);
output(1, 208) <= input(20);
output(1, 209) <= input(21);
output(1, 210) <= input(22);
output(1, 211) <= input(23);
output(1, 212) <= input(24);
output(1, 213) <= input(25);
output(1, 214) <= input(26);
output(1, 215) <= input(27);
output(1, 216) <= input(28);
output(1, 217) <= input(29);
output(1, 218) <= input(30);
output(1, 219) <= input(31);
output(1, 220) <= input(33);
output(1, 221) <= input(35);
output(1, 222) <= input(37);
output(1, 223) <= input(39);
output(1, 224) <= input(20);
output(1, 225) <= input(21);
output(1, 226) <= input(22);
output(1, 227) <= input(23);
output(1, 228) <= input(24);
output(1, 229) <= input(25);
output(1, 230) <= input(26);
output(1, 231) <= input(27);
output(1, 232) <= input(28);
output(1, 233) <= input(29);
output(1, 234) <= input(30);
output(1, 235) <= input(31);
output(1, 236) <= input(33);
output(1, 237) <= input(35);
output(1, 238) <= input(37);
output(1, 239) <= input(39);
output(1, 240) <= input(5);
output(1, 241) <= input(6);
output(1, 242) <= input(7);
output(1, 243) <= input(8);
output(1, 244) <= input(9);
output(1, 245) <= input(10);
output(1, 246) <= input(11);
output(1, 247) <= input(12);
output(1, 248) <= input(13);
output(1, 249) <= input(14);
output(1, 250) <= input(15);
output(1, 251) <= input(32);
output(1, 252) <= input(34);
output(1, 253) <= input(36);
output(1, 254) <= input(38);
output(1, 255) <= input(40);
output(2, 0) <= input(2);
output(2, 1) <= input(3);
output(2, 2) <= input(4);
output(2, 3) <= input(5);
output(2, 4) <= input(6);
output(2, 5) <= input(7);
output(2, 6) <= input(8);
output(2, 7) <= input(9);
output(2, 8) <= input(10);
output(2, 9) <= input(11);
output(2, 10) <= input(12);
output(2, 11) <= input(13);
output(2, 12) <= input(14);
output(2, 13) <= input(15);
output(2, 14) <= input(32);
output(2, 15) <= input(34);
output(2, 16) <= input(18);
output(2, 17) <= input(19);
output(2, 18) <= input(20);
output(2, 19) <= input(21);
output(2, 20) <= input(22);
output(2, 21) <= input(23);
output(2, 22) <= input(24);
output(2, 23) <= input(25);
output(2, 24) <= input(26);
output(2, 25) <= input(27);
output(2, 26) <= input(28);
output(2, 27) <= input(29);
output(2, 28) <= input(30);
output(2, 29) <= input(31);
output(2, 30) <= input(33);
output(2, 31) <= input(35);
output(2, 32) <= input(18);
output(2, 33) <= input(19);
output(2, 34) <= input(20);
output(2, 35) <= input(21);
output(2, 36) <= input(22);
output(2, 37) <= input(23);
output(2, 38) <= input(24);
output(2, 39) <= input(25);
output(2, 40) <= input(26);
output(2, 41) <= input(27);
output(2, 42) <= input(28);
output(2, 43) <= input(29);
output(2, 44) <= input(30);
output(2, 45) <= input(31);
output(2, 46) <= input(33);
output(2, 47) <= input(35);
output(2, 48) <= input(3);
output(2, 49) <= input(4);
output(2, 50) <= input(5);
output(2, 51) <= input(6);
output(2, 52) <= input(7);
output(2, 53) <= input(8);
output(2, 54) <= input(9);
output(2, 55) <= input(10);
output(2, 56) <= input(11);
output(2, 57) <= input(12);
output(2, 58) <= input(13);
output(2, 59) <= input(14);
output(2, 60) <= input(15);
output(2, 61) <= input(32);
output(2, 62) <= input(34);
output(2, 63) <= input(36);
output(2, 64) <= input(19);
output(2, 65) <= input(20);
output(2, 66) <= input(21);
output(2, 67) <= input(22);
output(2, 68) <= input(23);
output(2, 69) <= input(24);
output(2, 70) <= input(25);
output(2, 71) <= input(26);
output(2, 72) <= input(27);
output(2, 73) <= input(28);
output(2, 74) <= input(29);
output(2, 75) <= input(30);
output(2, 76) <= input(31);
output(2, 77) <= input(33);
output(2, 78) <= input(35);
output(2, 79) <= input(37);
output(2, 80) <= input(19);
output(2, 81) <= input(20);
output(2, 82) <= input(21);
output(2, 83) <= input(22);
output(2, 84) <= input(23);
output(2, 85) <= input(24);
output(2, 86) <= input(25);
output(2, 87) <= input(26);
output(2, 88) <= input(27);
output(2, 89) <= input(28);
output(2, 90) <= input(29);
output(2, 91) <= input(30);
output(2, 92) <= input(31);
output(2, 93) <= input(33);
output(2, 94) <= input(35);
output(2, 95) <= input(37);
output(2, 96) <= input(4);
output(2, 97) <= input(5);
output(2, 98) <= input(6);
output(2, 99) <= input(7);
output(2, 100) <= input(8);
output(2, 101) <= input(9);
output(2, 102) <= input(10);
output(2, 103) <= input(11);
output(2, 104) <= input(12);
output(2, 105) <= input(13);
output(2, 106) <= input(14);
output(2, 107) <= input(15);
output(2, 108) <= input(32);
output(2, 109) <= input(34);
output(2, 110) <= input(36);
output(2, 111) <= input(38);
output(2, 112) <= input(20);
output(2, 113) <= input(21);
output(2, 114) <= input(22);
output(2, 115) <= input(23);
output(2, 116) <= input(24);
output(2, 117) <= input(25);
output(2, 118) <= input(26);
output(2, 119) <= input(27);
output(2, 120) <= input(28);
output(2, 121) <= input(29);
output(2, 122) <= input(30);
output(2, 123) <= input(31);
output(2, 124) <= input(33);
output(2, 125) <= input(35);
output(2, 126) <= input(37);
output(2, 127) <= input(39);
output(2, 128) <= input(20);
output(2, 129) <= input(21);
output(2, 130) <= input(22);
output(2, 131) <= input(23);
output(2, 132) <= input(24);
output(2, 133) <= input(25);
output(2, 134) <= input(26);
output(2, 135) <= input(27);
output(2, 136) <= input(28);
output(2, 137) <= input(29);
output(2, 138) <= input(30);
output(2, 139) <= input(31);
output(2, 140) <= input(33);
output(2, 141) <= input(35);
output(2, 142) <= input(37);
output(2, 143) <= input(39);
output(2, 144) <= input(5);
output(2, 145) <= input(6);
output(2, 146) <= input(7);
output(2, 147) <= input(8);
output(2, 148) <= input(9);
output(2, 149) <= input(10);
output(2, 150) <= input(11);
output(2, 151) <= input(12);
output(2, 152) <= input(13);
output(2, 153) <= input(14);
output(2, 154) <= input(15);
output(2, 155) <= input(32);
output(2, 156) <= input(34);
output(2, 157) <= input(36);
output(2, 158) <= input(38);
output(2, 159) <= input(40);
output(2, 160) <= input(5);
output(2, 161) <= input(6);
output(2, 162) <= input(7);
output(2, 163) <= input(8);
output(2, 164) <= input(9);
output(2, 165) <= input(10);
output(2, 166) <= input(11);
output(2, 167) <= input(12);
output(2, 168) <= input(13);
output(2, 169) <= input(14);
output(2, 170) <= input(15);
output(2, 171) <= input(32);
output(2, 172) <= input(34);
output(2, 173) <= input(36);
output(2, 174) <= input(38);
output(2, 175) <= input(40);
output(2, 176) <= input(21);
output(2, 177) <= input(22);
output(2, 178) <= input(23);
output(2, 179) <= input(24);
output(2, 180) <= input(25);
output(2, 181) <= input(26);
output(2, 182) <= input(27);
output(2, 183) <= input(28);
output(2, 184) <= input(29);
output(2, 185) <= input(30);
output(2, 186) <= input(31);
output(2, 187) <= input(33);
output(2, 188) <= input(35);
output(2, 189) <= input(37);
output(2, 190) <= input(39);
output(2, 191) <= input(41);
output(2, 192) <= input(6);
output(2, 193) <= input(7);
output(2, 194) <= input(8);
output(2, 195) <= input(9);
output(2, 196) <= input(10);
output(2, 197) <= input(11);
output(2, 198) <= input(12);
output(2, 199) <= input(13);
output(2, 200) <= input(14);
output(2, 201) <= input(15);
output(2, 202) <= input(32);
output(2, 203) <= input(34);
output(2, 204) <= input(36);
output(2, 205) <= input(38);
output(2, 206) <= input(40);
output(2, 207) <= input(42);
output(2, 208) <= input(6);
output(2, 209) <= input(7);
output(2, 210) <= input(8);
output(2, 211) <= input(9);
output(2, 212) <= input(10);
output(2, 213) <= input(11);
output(2, 214) <= input(12);
output(2, 215) <= input(13);
output(2, 216) <= input(14);
output(2, 217) <= input(15);
output(2, 218) <= input(32);
output(2, 219) <= input(34);
output(2, 220) <= input(36);
output(2, 221) <= input(38);
output(2, 222) <= input(40);
output(2, 223) <= input(42);
output(2, 224) <= input(22);
output(2, 225) <= input(23);
output(2, 226) <= input(24);
output(2, 227) <= input(25);
output(2, 228) <= input(26);
output(2, 229) <= input(27);
output(2, 230) <= input(28);
output(2, 231) <= input(29);
output(2, 232) <= input(30);
output(2, 233) <= input(31);
output(2, 234) <= input(33);
output(2, 235) <= input(35);
output(2, 236) <= input(37);
output(2, 237) <= input(39);
output(2, 238) <= input(41);
output(2, 239) <= input(43);
output(2, 240) <= input(7);
output(2, 241) <= input(8);
output(2, 242) <= input(9);
output(2, 243) <= input(10);
output(2, 244) <= input(11);
output(2, 245) <= input(12);
output(2, 246) <= input(13);
output(2, 247) <= input(14);
output(2, 248) <= input(15);
output(2, 249) <= input(32);
output(2, 250) <= input(34);
output(2, 251) <= input(36);
output(2, 252) <= input(38);
output(2, 253) <= input(40);
output(2, 254) <= input(42);
output(2, 255) <= input(44);
output(3, 0) <= input(3);
output(3, 1) <= input(4);
output(3, 2) <= input(5);
output(3, 3) <= input(6);
output(3, 4) <= input(7);
output(3, 5) <= input(8);
output(3, 6) <= input(9);
output(3, 7) <= input(10);
output(3, 8) <= input(11);
output(3, 9) <= input(12);
output(3, 10) <= input(13);
output(3, 11) <= input(14);
output(3, 12) <= input(15);
output(3, 13) <= input(32);
output(3, 14) <= input(34);
output(3, 15) <= input(36);
output(3, 16) <= input(19);
output(3, 17) <= input(20);
output(3, 18) <= input(21);
output(3, 19) <= input(22);
output(3, 20) <= input(23);
output(3, 21) <= input(24);
output(3, 22) <= input(25);
output(3, 23) <= input(26);
output(3, 24) <= input(27);
output(3, 25) <= input(28);
output(3, 26) <= input(29);
output(3, 27) <= input(30);
output(3, 28) <= input(31);
output(3, 29) <= input(33);
output(3, 30) <= input(35);
output(3, 31) <= input(37);
output(3, 32) <= input(4);
output(3, 33) <= input(5);
output(3, 34) <= input(6);
output(3, 35) <= input(7);
output(3, 36) <= input(8);
output(3, 37) <= input(9);
output(3, 38) <= input(10);
output(3, 39) <= input(11);
output(3, 40) <= input(12);
output(3, 41) <= input(13);
output(3, 42) <= input(14);
output(3, 43) <= input(15);
output(3, 44) <= input(32);
output(3, 45) <= input(34);
output(3, 46) <= input(36);
output(3, 47) <= input(38);
output(3, 48) <= input(20);
output(3, 49) <= input(21);
output(3, 50) <= input(22);
output(3, 51) <= input(23);
output(3, 52) <= input(24);
output(3, 53) <= input(25);
output(3, 54) <= input(26);
output(3, 55) <= input(27);
output(3, 56) <= input(28);
output(3, 57) <= input(29);
output(3, 58) <= input(30);
output(3, 59) <= input(31);
output(3, 60) <= input(33);
output(3, 61) <= input(35);
output(3, 62) <= input(37);
output(3, 63) <= input(39);
output(3, 64) <= input(20);
output(3, 65) <= input(21);
output(3, 66) <= input(22);
output(3, 67) <= input(23);
output(3, 68) <= input(24);
output(3, 69) <= input(25);
output(3, 70) <= input(26);
output(3, 71) <= input(27);
output(3, 72) <= input(28);
output(3, 73) <= input(29);
output(3, 74) <= input(30);
output(3, 75) <= input(31);
output(3, 76) <= input(33);
output(3, 77) <= input(35);
output(3, 78) <= input(37);
output(3, 79) <= input(39);
output(3, 80) <= input(5);
output(3, 81) <= input(6);
output(3, 82) <= input(7);
output(3, 83) <= input(8);
output(3, 84) <= input(9);
output(3, 85) <= input(10);
output(3, 86) <= input(11);
output(3, 87) <= input(12);
output(3, 88) <= input(13);
output(3, 89) <= input(14);
output(3, 90) <= input(15);
output(3, 91) <= input(32);
output(3, 92) <= input(34);
output(3, 93) <= input(36);
output(3, 94) <= input(38);
output(3, 95) <= input(40);
output(3, 96) <= input(21);
output(3, 97) <= input(22);
output(3, 98) <= input(23);
output(3, 99) <= input(24);
output(3, 100) <= input(25);
output(3, 101) <= input(26);
output(3, 102) <= input(27);
output(3, 103) <= input(28);
output(3, 104) <= input(29);
output(3, 105) <= input(30);
output(3, 106) <= input(31);
output(3, 107) <= input(33);
output(3, 108) <= input(35);
output(3, 109) <= input(37);
output(3, 110) <= input(39);
output(3, 111) <= input(41);
output(3, 112) <= input(6);
output(3, 113) <= input(7);
output(3, 114) <= input(8);
output(3, 115) <= input(9);
output(3, 116) <= input(10);
output(3, 117) <= input(11);
output(3, 118) <= input(12);
output(3, 119) <= input(13);
output(3, 120) <= input(14);
output(3, 121) <= input(15);
output(3, 122) <= input(32);
output(3, 123) <= input(34);
output(3, 124) <= input(36);
output(3, 125) <= input(38);
output(3, 126) <= input(40);
output(3, 127) <= input(42);
output(3, 128) <= input(6);
output(3, 129) <= input(7);
output(3, 130) <= input(8);
output(3, 131) <= input(9);
output(3, 132) <= input(10);
output(3, 133) <= input(11);
output(3, 134) <= input(12);
output(3, 135) <= input(13);
output(3, 136) <= input(14);
output(3, 137) <= input(15);
output(3, 138) <= input(32);
output(3, 139) <= input(34);
output(3, 140) <= input(36);
output(3, 141) <= input(38);
output(3, 142) <= input(40);
output(3, 143) <= input(42);
output(3, 144) <= input(22);
output(3, 145) <= input(23);
output(3, 146) <= input(24);
output(3, 147) <= input(25);
output(3, 148) <= input(26);
output(3, 149) <= input(27);
output(3, 150) <= input(28);
output(3, 151) <= input(29);
output(3, 152) <= input(30);
output(3, 153) <= input(31);
output(3, 154) <= input(33);
output(3, 155) <= input(35);
output(3, 156) <= input(37);
output(3, 157) <= input(39);
output(3, 158) <= input(41);
output(3, 159) <= input(43);
output(3, 160) <= input(7);
output(3, 161) <= input(8);
output(3, 162) <= input(9);
output(3, 163) <= input(10);
output(3, 164) <= input(11);
output(3, 165) <= input(12);
output(3, 166) <= input(13);
output(3, 167) <= input(14);
output(3, 168) <= input(15);
output(3, 169) <= input(32);
output(3, 170) <= input(34);
output(3, 171) <= input(36);
output(3, 172) <= input(38);
output(3, 173) <= input(40);
output(3, 174) <= input(42);
output(3, 175) <= input(44);
output(3, 176) <= input(23);
output(3, 177) <= input(24);
output(3, 178) <= input(25);
output(3, 179) <= input(26);
output(3, 180) <= input(27);
output(3, 181) <= input(28);
output(3, 182) <= input(29);
output(3, 183) <= input(30);
output(3, 184) <= input(31);
output(3, 185) <= input(33);
output(3, 186) <= input(35);
output(3, 187) <= input(37);
output(3, 188) <= input(39);
output(3, 189) <= input(41);
output(3, 190) <= input(43);
output(3, 191) <= input(45);
output(3, 192) <= input(23);
output(3, 193) <= input(24);
output(3, 194) <= input(25);
output(3, 195) <= input(26);
output(3, 196) <= input(27);
output(3, 197) <= input(28);
output(3, 198) <= input(29);
output(3, 199) <= input(30);
output(3, 200) <= input(31);
output(3, 201) <= input(33);
output(3, 202) <= input(35);
output(3, 203) <= input(37);
output(3, 204) <= input(39);
output(3, 205) <= input(41);
output(3, 206) <= input(43);
output(3, 207) <= input(45);
output(3, 208) <= input(8);
output(3, 209) <= input(9);
output(3, 210) <= input(10);
output(3, 211) <= input(11);
output(3, 212) <= input(12);
output(3, 213) <= input(13);
output(3, 214) <= input(14);
output(3, 215) <= input(15);
output(3, 216) <= input(32);
output(3, 217) <= input(34);
output(3, 218) <= input(36);
output(3, 219) <= input(38);
output(3, 220) <= input(40);
output(3, 221) <= input(42);
output(3, 222) <= input(44);
output(3, 223) <= input(46);
output(3, 224) <= input(24);
output(3, 225) <= input(25);
output(3, 226) <= input(26);
output(3, 227) <= input(27);
output(3, 228) <= input(28);
output(3, 229) <= input(29);
output(3, 230) <= input(30);
output(3, 231) <= input(31);
output(3, 232) <= input(33);
output(3, 233) <= input(35);
output(3, 234) <= input(37);
output(3, 235) <= input(39);
output(3, 236) <= input(41);
output(3, 237) <= input(43);
output(3, 238) <= input(45);
output(3, 239) <= input(47);
output(3, 240) <= input(9);
output(3, 241) <= input(10);
output(3, 242) <= input(11);
output(3, 243) <= input(12);
output(3, 244) <= input(13);
output(3, 245) <= input(14);
output(3, 246) <= input(15);
output(3, 247) <= input(32);
output(3, 248) <= input(34);
output(3, 249) <= input(36);
output(3, 250) <= input(38);
output(3, 251) <= input(40);
output(3, 252) <= input(42);
output(3, 253) <= input(44);
output(3, 254) <= input(46);
output(3, 255) <= input(48);
output(4, 0) <= input(4);
output(4, 1) <= input(5);
output(4, 2) <= input(6);
output(4, 3) <= input(7);
output(4, 4) <= input(8);
output(4, 5) <= input(9);
output(4, 6) <= input(10);
output(4, 7) <= input(11);
output(4, 8) <= input(12);
output(4, 9) <= input(13);
output(4, 10) <= input(14);
output(4, 11) <= input(15);
output(4, 12) <= input(32);
output(4, 13) <= input(34);
output(4, 14) <= input(36);
output(4, 15) <= input(38);
output(4, 16) <= input(20);
output(4, 17) <= input(21);
output(4, 18) <= input(22);
output(4, 19) <= input(23);
output(4, 20) <= input(24);
output(4, 21) <= input(25);
output(4, 22) <= input(26);
output(4, 23) <= input(27);
output(4, 24) <= input(28);
output(4, 25) <= input(29);
output(4, 26) <= input(30);
output(4, 27) <= input(31);
output(4, 28) <= input(33);
output(4, 29) <= input(35);
output(4, 30) <= input(37);
output(4, 31) <= input(39);
output(4, 32) <= input(5);
output(4, 33) <= input(6);
output(4, 34) <= input(7);
output(4, 35) <= input(8);
output(4, 36) <= input(9);
output(4, 37) <= input(10);
output(4, 38) <= input(11);
output(4, 39) <= input(12);
output(4, 40) <= input(13);
output(4, 41) <= input(14);
output(4, 42) <= input(15);
output(4, 43) <= input(32);
output(4, 44) <= input(34);
output(4, 45) <= input(36);
output(4, 46) <= input(38);
output(4, 47) <= input(40);
output(4, 48) <= input(21);
output(4, 49) <= input(22);
output(4, 50) <= input(23);
output(4, 51) <= input(24);
output(4, 52) <= input(25);
output(4, 53) <= input(26);
output(4, 54) <= input(27);
output(4, 55) <= input(28);
output(4, 56) <= input(29);
output(4, 57) <= input(30);
output(4, 58) <= input(31);
output(4, 59) <= input(33);
output(4, 60) <= input(35);
output(4, 61) <= input(37);
output(4, 62) <= input(39);
output(4, 63) <= input(41);
output(4, 64) <= input(6);
output(4, 65) <= input(7);
output(4, 66) <= input(8);
output(4, 67) <= input(9);
output(4, 68) <= input(10);
output(4, 69) <= input(11);
output(4, 70) <= input(12);
output(4, 71) <= input(13);
output(4, 72) <= input(14);
output(4, 73) <= input(15);
output(4, 74) <= input(32);
output(4, 75) <= input(34);
output(4, 76) <= input(36);
output(4, 77) <= input(38);
output(4, 78) <= input(40);
output(4, 79) <= input(42);
output(4, 80) <= input(22);
output(4, 81) <= input(23);
output(4, 82) <= input(24);
output(4, 83) <= input(25);
output(4, 84) <= input(26);
output(4, 85) <= input(27);
output(4, 86) <= input(28);
output(4, 87) <= input(29);
output(4, 88) <= input(30);
output(4, 89) <= input(31);
output(4, 90) <= input(33);
output(4, 91) <= input(35);
output(4, 92) <= input(37);
output(4, 93) <= input(39);
output(4, 94) <= input(41);
output(4, 95) <= input(43);
output(4, 96) <= input(7);
output(4, 97) <= input(8);
output(4, 98) <= input(9);
output(4, 99) <= input(10);
output(4, 100) <= input(11);
output(4, 101) <= input(12);
output(4, 102) <= input(13);
output(4, 103) <= input(14);
output(4, 104) <= input(15);
output(4, 105) <= input(32);
output(4, 106) <= input(34);
output(4, 107) <= input(36);
output(4, 108) <= input(38);
output(4, 109) <= input(40);
output(4, 110) <= input(42);
output(4, 111) <= input(44);
output(4, 112) <= input(23);
output(4, 113) <= input(24);
output(4, 114) <= input(25);
output(4, 115) <= input(26);
output(4, 116) <= input(27);
output(4, 117) <= input(28);
output(4, 118) <= input(29);
output(4, 119) <= input(30);
output(4, 120) <= input(31);
output(4, 121) <= input(33);
output(4, 122) <= input(35);
output(4, 123) <= input(37);
output(4, 124) <= input(39);
output(4, 125) <= input(41);
output(4, 126) <= input(43);
output(4, 127) <= input(45);
output(4, 128) <= input(23);
output(4, 129) <= input(24);
output(4, 130) <= input(25);
output(4, 131) <= input(26);
output(4, 132) <= input(27);
output(4, 133) <= input(28);
output(4, 134) <= input(29);
output(4, 135) <= input(30);
output(4, 136) <= input(31);
output(4, 137) <= input(33);
output(4, 138) <= input(35);
output(4, 139) <= input(37);
output(4, 140) <= input(39);
output(4, 141) <= input(41);
output(4, 142) <= input(43);
output(4, 143) <= input(45);
output(4, 144) <= input(8);
output(4, 145) <= input(9);
output(4, 146) <= input(10);
output(4, 147) <= input(11);
output(4, 148) <= input(12);
output(4, 149) <= input(13);
output(4, 150) <= input(14);
output(4, 151) <= input(15);
output(4, 152) <= input(32);
output(4, 153) <= input(34);
output(4, 154) <= input(36);
output(4, 155) <= input(38);
output(4, 156) <= input(40);
output(4, 157) <= input(42);
output(4, 158) <= input(44);
output(4, 159) <= input(46);
output(4, 160) <= input(24);
output(4, 161) <= input(25);
output(4, 162) <= input(26);
output(4, 163) <= input(27);
output(4, 164) <= input(28);
output(4, 165) <= input(29);
output(4, 166) <= input(30);
output(4, 167) <= input(31);
output(4, 168) <= input(33);
output(4, 169) <= input(35);
output(4, 170) <= input(37);
output(4, 171) <= input(39);
output(4, 172) <= input(41);
output(4, 173) <= input(43);
output(4, 174) <= input(45);
output(4, 175) <= input(47);
output(4, 176) <= input(9);
output(4, 177) <= input(10);
output(4, 178) <= input(11);
output(4, 179) <= input(12);
output(4, 180) <= input(13);
output(4, 181) <= input(14);
output(4, 182) <= input(15);
output(4, 183) <= input(32);
output(4, 184) <= input(34);
output(4, 185) <= input(36);
output(4, 186) <= input(38);
output(4, 187) <= input(40);
output(4, 188) <= input(42);
output(4, 189) <= input(44);
output(4, 190) <= input(46);
output(4, 191) <= input(48);
output(4, 192) <= input(25);
output(4, 193) <= input(26);
output(4, 194) <= input(27);
output(4, 195) <= input(28);
output(4, 196) <= input(29);
output(4, 197) <= input(30);
output(4, 198) <= input(31);
output(4, 199) <= input(33);
output(4, 200) <= input(35);
output(4, 201) <= input(37);
output(4, 202) <= input(39);
output(4, 203) <= input(41);
output(4, 204) <= input(43);
output(4, 205) <= input(45);
output(4, 206) <= input(47);
output(4, 207) <= input(49);
output(4, 208) <= input(10);
output(4, 209) <= input(11);
output(4, 210) <= input(12);
output(4, 211) <= input(13);
output(4, 212) <= input(14);
output(4, 213) <= input(15);
output(4, 214) <= input(32);
output(4, 215) <= input(34);
output(4, 216) <= input(36);
output(4, 217) <= input(38);
output(4, 218) <= input(40);
output(4, 219) <= input(42);
output(4, 220) <= input(44);
output(4, 221) <= input(46);
output(4, 222) <= input(48);
output(4, 223) <= input(50);
output(4, 224) <= input(26);
output(4, 225) <= input(27);
output(4, 226) <= input(28);
output(4, 227) <= input(29);
output(4, 228) <= input(30);
output(4, 229) <= input(31);
output(4, 230) <= input(33);
output(4, 231) <= input(35);
output(4, 232) <= input(37);
output(4, 233) <= input(39);
output(4, 234) <= input(41);
output(4, 235) <= input(43);
output(4, 236) <= input(45);
output(4, 237) <= input(47);
output(4, 238) <= input(49);
output(4, 239) <= input(51);
output(4, 240) <= input(11);
output(4, 241) <= input(12);
output(4, 242) <= input(13);
output(4, 243) <= input(14);
output(4, 244) <= input(15);
output(4, 245) <= input(32);
output(4, 246) <= input(34);
output(4, 247) <= input(36);
output(4, 248) <= input(38);
output(4, 249) <= input(40);
output(4, 250) <= input(42);
output(4, 251) <= input(44);
output(4, 252) <= input(46);
output(4, 253) <= input(48);
output(4, 254) <= input(50);
output(4, 255) <= input(52);
output(5, 0) <= input(21);
output(5, 1) <= input(22);
output(5, 2) <= input(23);
output(5, 3) <= input(24);
output(5, 4) <= input(25);
output(5, 5) <= input(26);
output(5, 6) <= input(27);
output(5, 7) <= input(28);
output(5, 8) <= input(29);
output(5, 9) <= input(30);
output(5, 10) <= input(31);
output(5, 11) <= input(33);
output(5, 12) <= input(35);
output(5, 13) <= input(37);
output(5, 14) <= input(39);
output(5, 15) <= input(41);
output(5, 16) <= input(6);
output(5, 17) <= input(7);
output(5, 18) <= input(8);
output(5, 19) <= input(9);
output(5, 20) <= input(10);
output(5, 21) <= input(11);
output(5, 22) <= input(12);
output(5, 23) <= input(13);
output(5, 24) <= input(14);
output(5, 25) <= input(15);
output(5, 26) <= input(32);
output(5, 27) <= input(34);
output(5, 28) <= input(36);
output(5, 29) <= input(38);
output(5, 30) <= input(40);
output(5, 31) <= input(42);
output(5, 32) <= input(22);
output(5, 33) <= input(23);
output(5, 34) <= input(24);
output(5, 35) <= input(25);
output(5, 36) <= input(26);
output(5, 37) <= input(27);
output(5, 38) <= input(28);
output(5, 39) <= input(29);
output(5, 40) <= input(30);
output(5, 41) <= input(31);
output(5, 42) <= input(33);
output(5, 43) <= input(35);
output(5, 44) <= input(37);
output(5, 45) <= input(39);
output(5, 46) <= input(41);
output(5, 47) <= input(43);
output(5, 48) <= input(7);
output(5, 49) <= input(8);
output(5, 50) <= input(9);
output(5, 51) <= input(10);
output(5, 52) <= input(11);
output(5, 53) <= input(12);
output(5, 54) <= input(13);
output(5, 55) <= input(14);
output(5, 56) <= input(15);
output(5, 57) <= input(32);
output(5, 58) <= input(34);
output(5, 59) <= input(36);
output(5, 60) <= input(38);
output(5, 61) <= input(40);
output(5, 62) <= input(42);
output(5, 63) <= input(44);
output(5, 64) <= input(23);
output(5, 65) <= input(24);
output(5, 66) <= input(25);
output(5, 67) <= input(26);
output(5, 68) <= input(27);
output(5, 69) <= input(28);
output(5, 70) <= input(29);
output(5, 71) <= input(30);
output(5, 72) <= input(31);
output(5, 73) <= input(33);
output(5, 74) <= input(35);
output(5, 75) <= input(37);
output(5, 76) <= input(39);
output(5, 77) <= input(41);
output(5, 78) <= input(43);
output(5, 79) <= input(45);
output(5, 80) <= input(8);
output(5, 81) <= input(9);
output(5, 82) <= input(10);
output(5, 83) <= input(11);
output(5, 84) <= input(12);
output(5, 85) <= input(13);
output(5, 86) <= input(14);
output(5, 87) <= input(15);
output(5, 88) <= input(32);
output(5, 89) <= input(34);
output(5, 90) <= input(36);
output(5, 91) <= input(38);
output(5, 92) <= input(40);
output(5, 93) <= input(42);
output(5, 94) <= input(44);
output(5, 95) <= input(46);
output(5, 96) <= input(24);
output(5, 97) <= input(25);
output(5, 98) <= input(26);
output(5, 99) <= input(27);
output(5, 100) <= input(28);
output(5, 101) <= input(29);
output(5, 102) <= input(30);
output(5, 103) <= input(31);
output(5, 104) <= input(33);
output(5, 105) <= input(35);
output(5, 106) <= input(37);
output(5, 107) <= input(39);
output(5, 108) <= input(41);
output(5, 109) <= input(43);
output(5, 110) <= input(45);
output(5, 111) <= input(47);
output(5, 112) <= input(9);
output(5, 113) <= input(10);
output(5, 114) <= input(11);
output(5, 115) <= input(12);
output(5, 116) <= input(13);
output(5, 117) <= input(14);
output(5, 118) <= input(15);
output(5, 119) <= input(32);
output(5, 120) <= input(34);
output(5, 121) <= input(36);
output(5, 122) <= input(38);
output(5, 123) <= input(40);
output(5, 124) <= input(42);
output(5, 125) <= input(44);
output(5, 126) <= input(46);
output(5, 127) <= input(48);
output(5, 128) <= input(25);
output(5, 129) <= input(26);
output(5, 130) <= input(27);
output(5, 131) <= input(28);
output(5, 132) <= input(29);
output(5, 133) <= input(30);
output(5, 134) <= input(31);
output(5, 135) <= input(33);
output(5, 136) <= input(35);
output(5, 137) <= input(37);
output(5, 138) <= input(39);
output(5, 139) <= input(41);
output(5, 140) <= input(43);
output(5, 141) <= input(45);
output(5, 142) <= input(47);
output(5, 143) <= input(49);
output(5, 144) <= input(10);
output(5, 145) <= input(11);
output(5, 146) <= input(12);
output(5, 147) <= input(13);
output(5, 148) <= input(14);
output(5, 149) <= input(15);
output(5, 150) <= input(32);
output(5, 151) <= input(34);
output(5, 152) <= input(36);
output(5, 153) <= input(38);
output(5, 154) <= input(40);
output(5, 155) <= input(42);
output(5, 156) <= input(44);
output(5, 157) <= input(46);
output(5, 158) <= input(48);
output(5, 159) <= input(50);
output(5, 160) <= input(26);
output(5, 161) <= input(27);
output(5, 162) <= input(28);
output(5, 163) <= input(29);
output(5, 164) <= input(30);
output(5, 165) <= input(31);
output(5, 166) <= input(33);
output(5, 167) <= input(35);
output(5, 168) <= input(37);
output(5, 169) <= input(39);
output(5, 170) <= input(41);
output(5, 171) <= input(43);
output(5, 172) <= input(45);
output(5, 173) <= input(47);
output(5, 174) <= input(49);
output(5, 175) <= input(51);
output(5, 176) <= input(11);
output(5, 177) <= input(12);
output(5, 178) <= input(13);
output(5, 179) <= input(14);
output(5, 180) <= input(15);
output(5, 181) <= input(32);
output(5, 182) <= input(34);
output(5, 183) <= input(36);
output(5, 184) <= input(38);
output(5, 185) <= input(40);
output(5, 186) <= input(42);
output(5, 187) <= input(44);
output(5, 188) <= input(46);
output(5, 189) <= input(48);
output(5, 190) <= input(50);
output(5, 191) <= input(52);
output(5, 192) <= input(27);
output(5, 193) <= input(28);
output(5, 194) <= input(29);
output(5, 195) <= input(30);
output(5, 196) <= input(31);
output(5, 197) <= input(33);
output(5, 198) <= input(35);
output(5, 199) <= input(37);
output(5, 200) <= input(39);
output(5, 201) <= input(41);
output(5, 202) <= input(43);
output(5, 203) <= input(45);
output(5, 204) <= input(47);
output(5, 205) <= input(49);
output(5, 206) <= input(51);
output(5, 207) <= input(53);
output(5, 208) <= input(12);
output(5, 209) <= input(13);
output(5, 210) <= input(14);
output(5, 211) <= input(15);
output(5, 212) <= input(32);
output(5, 213) <= input(34);
output(5, 214) <= input(36);
output(5, 215) <= input(38);
output(5, 216) <= input(40);
output(5, 217) <= input(42);
output(5, 218) <= input(44);
output(5, 219) <= input(46);
output(5, 220) <= input(48);
output(5, 221) <= input(50);
output(5, 222) <= input(52);
output(5, 223) <= input(54);
output(5, 224) <= input(28);
output(5, 225) <= input(29);
output(5, 226) <= input(30);
output(5, 227) <= input(31);
output(5, 228) <= input(33);
output(5, 229) <= input(35);
output(5, 230) <= input(37);
output(5, 231) <= input(39);
output(5, 232) <= input(41);
output(5, 233) <= input(43);
output(5, 234) <= input(45);
output(5, 235) <= input(47);
output(5, 236) <= input(49);
output(5, 237) <= input(51);
output(5, 238) <= input(53);
output(5, 239) <= input(55);
output(5, 240) <= input(13);
output(5, 241) <= input(14);
output(5, 242) <= input(15);
output(5, 243) <= input(32);
output(5, 244) <= input(34);
output(5, 245) <= input(36);
output(5, 246) <= input(38);
output(5, 247) <= input(40);
output(5, 248) <= input(42);
output(5, 249) <= input(44);
output(5, 250) <= input(46);
output(5, 251) <= input(48);
output(5, 252) <= input(50);
output(5, 253) <= input(52);
output(5, 254) <= input(54);
output(5, 255) <= input(56);
when "1111" =>
output(0, 0) <= input(0);
output(0, 1) <= input(1);
output(0, 2) <= input(2);
output(0, 3) <= input(3);
output(0, 4) <= input(4);
output(0, 5) <= input(5);
output(0, 6) <= input(6);
output(0, 7) <= input(7);
output(0, 8) <= input(8);
output(0, 9) <= input(9);
output(0, 10) <= input(10);
output(0, 11) <= input(11);
output(0, 12) <= input(12);
output(0, 13) <= input(13);
output(0, 14) <= input(14);
output(0, 15) <= input(15);
output(0, 16) <= input(16);
output(0, 17) <= input(17);
output(0, 18) <= input(18);
output(0, 19) <= input(19);
output(0, 20) <= input(20);
output(0, 21) <= input(21);
output(0, 22) <= input(22);
output(0, 23) <= input(23);
output(0, 24) <= input(24);
output(0, 25) <= input(25);
output(0, 26) <= input(26);
output(0, 27) <= input(27);
output(0, 28) <= input(28);
output(0, 29) <= input(29);
output(0, 30) <= input(30);
output(0, 31) <= input(31);
output(0, 32) <= input(1);
output(0, 33) <= input(2);
output(0, 34) <= input(3);
output(0, 35) <= input(4);
output(0, 36) <= input(5);
output(0, 37) <= input(6);
output(0, 38) <= input(7);
output(0, 39) <= input(8);
output(0, 40) <= input(9);
output(0, 41) <= input(10);
output(0, 42) <= input(11);
output(0, 43) <= input(12);
output(0, 44) <= input(13);
output(0, 45) <= input(14);
output(0, 46) <= input(15);
output(0, 47) <= input(32);
output(0, 48) <= input(17);
output(0, 49) <= input(18);
output(0, 50) <= input(19);
output(0, 51) <= input(20);
output(0, 52) <= input(21);
output(0, 53) <= input(22);
output(0, 54) <= input(23);
output(0, 55) <= input(24);
output(0, 56) <= input(25);
output(0, 57) <= input(26);
output(0, 58) <= input(27);
output(0, 59) <= input(28);
output(0, 60) <= input(29);
output(0, 61) <= input(30);
output(0, 62) <= input(31);
output(0, 63) <= input(33);
output(0, 64) <= input(2);
output(0, 65) <= input(3);
output(0, 66) <= input(4);
output(0, 67) <= input(5);
output(0, 68) <= input(6);
output(0, 69) <= input(7);
output(0, 70) <= input(8);
output(0, 71) <= input(9);
output(0, 72) <= input(10);
output(0, 73) <= input(11);
output(0, 74) <= input(12);
output(0, 75) <= input(13);
output(0, 76) <= input(14);
output(0, 77) <= input(15);
output(0, 78) <= input(32);
output(0, 79) <= input(34);
output(0, 80) <= input(18);
output(0, 81) <= input(19);
output(0, 82) <= input(20);
output(0, 83) <= input(21);
output(0, 84) <= input(22);
output(0, 85) <= input(23);
output(0, 86) <= input(24);
output(0, 87) <= input(25);
output(0, 88) <= input(26);
output(0, 89) <= input(27);
output(0, 90) <= input(28);
output(0, 91) <= input(29);
output(0, 92) <= input(30);
output(0, 93) <= input(31);
output(0, 94) <= input(33);
output(0, 95) <= input(35);
output(0, 96) <= input(3);
output(0, 97) <= input(4);
output(0, 98) <= input(5);
output(0, 99) <= input(6);
output(0, 100) <= input(7);
output(0, 101) <= input(8);
output(0, 102) <= input(9);
output(0, 103) <= input(10);
output(0, 104) <= input(11);
output(0, 105) <= input(12);
output(0, 106) <= input(13);
output(0, 107) <= input(14);
output(0, 108) <= input(15);
output(0, 109) <= input(32);
output(0, 110) <= input(34);
output(0, 111) <= input(36);
output(0, 112) <= input(4);
output(0, 113) <= input(5);
output(0, 114) <= input(6);
output(0, 115) <= input(7);
output(0, 116) <= input(8);
output(0, 117) <= input(9);
output(0, 118) <= input(10);
output(0, 119) <= input(11);
output(0, 120) <= input(12);
output(0, 121) <= input(13);
output(0, 122) <= input(14);
output(0, 123) <= input(15);
output(0, 124) <= input(32);
output(0, 125) <= input(34);
output(0, 126) <= input(36);
output(0, 127) <= input(37);
output(0, 128) <= input(20);
output(0, 129) <= input(21);
output(0, 130) <= input(22);
output(0, 131) <= input(23);
output(0, 132) <= input(24);
output(0, 133) <= input(25);
output(0, 134) <= input(26);
output(0, 135) <= input(27);
output(0, 136) <= input(28);
output(0, 137) <= input(29);
output(0, 138) <= input(30);
output(0, 139) <= input(31);
output(0, 140) <= input(33);
output(0, 141) <= input(35);
output(0, 142) <= input(38);
output(0, 143) <= input(39);
output(0, 144) <= input(5);
output(0, 145) <= input(6);
output(0, 146) <= input(7);
output(0, 147) <= input(8);
output(0, 148) <= input(9);
output(0, 149) <= input(10);
output(0, 150) <= input(11);
output(0, 151) <= input(12);
output(0, 152) <= input(13);
output(0, 153) <= input(14);
output(0, 154) <= input(15);
output(0, 155) <= input(32);
output(0, 156) <= input(34);
output(0, 157) <= input(36);
output(0, 158) <= input(37);
output(0, 159) <= input(40);
output(0, 160) <= input(21);
output(0, 161) <= input(22);
output(0, 162) <= input(23);
output(0, 163) <= input(24);
output(0, 164) <= input(25);
output(0, 165) <= input(26);
output(0, 166) <= input(27);
output(0, 167) <= input(28);
output(0, 168) <= input(29);
output(0, 169) <= input(30);
output(0, 170) <= input(31);
output(0, 171) <= input(33);
output(0, 172) <= input(35);
output(0, 173) <= input(38);
output(0, 174) <= input(39);
output(0, 175) <= input(41);
output(0, 176) <= input(6);
output(0, 177) <= input(7);
output(0, 178) <= input(8);
output(0, 179) <= input(9);
output(0, 180) <= input(10);
output(0, 181) <= input(11);
output(0, 182) <= input(12);
output(0, 183) <= input(13);
output(0, 184) <= input(14);
output(0, 185) <= input(15);
output(0, 186) <= input(32);
output(0, 187) <= input(34);
output(0, 188) <= input(36);
output(0, 189) <= input(37);
output(0, 190) <= input(40);
output(0, 191) <= input(42);
output(0, 192) <= input(22);
output(0, 193) <= input(23);
output(0, 194) <= input(24);
output(0, 195) <= input(25);
output(0, 196) <= input(26);
output(0, 197) <= input(27);
output(0, 198) <= input(28);
output(0, 199) <= input(29);
output(0, 200) <= input(30);
output(0, 201) <= input(31);
output(0, 202) <= input(33);
output(0, 203) <= input(35);
output(0, 204) <= input(38);
output(0, 205) <= input(39);
output(0, 206) <= input(41);
output(0, 207) <= input(43);
output(0, 208) <= input(7);
output(0, 209) <= input(8);
output(0, 210) <= input(9);
output(0, 211) <= input(10);
output(0, 212) <= input(11);
output(0, 213) <= input(12);
output(0, 214) <= input(13);
output(0, 215) <= input(14);
output(0, 216) <= input(15);
output(0, 217) <= input(32);
output(0, 218) <= input(34);
output(0, 219) <= input(36);
output(0, 220) <= input(37);
output(0, 221) <= input(40);
output(0, 222) <= input(42);
output(0, 223) <= input(44);
output(0, 224) <= input(23);
output(0, 225) <= input(24);
output(0, 226) <= input(25);
output(0, 227) <= input(26);
output(0, 228) <= input(27);
output(0, 229) <= input(28);
output(0, 230) <= input(29);
output(0, 231) <= input(30);
output(0, 232) <= input(31);
output(0, 233) <= input(33);
output(0, 234) <= input(35);
output(0, 235) <= input(38);
output(0, 236) <= input(39);
output(0, 237) <= input(41);
output(0, 238) <= input(43);
output(0, 239) <= input(45);
output(0, 240) <= input(24);
output(0, 241) <= input(25);
output(0, 242) <= input(26);
output(0, 243) <= input(27);
output(0, 244) <= input(28);
output(0, 245) <= input(29);
output(0, 246) <= input(30);
output(0, 247) <= input(31);
output(0, 248) <= input(33);
output(0, 249) <= input(35);
output(0, 250) <= input(38);
output(0, 251) <= input(39);
output(0, 252) <= input(41);
output(0, 253) <= input(43);
output(0, 254) <= input(45);
output(0, 255) <= input(46);
output(1, 0) <= input(1);
output(1, 1) <= input(2);
output(1, 2) <= input(3);
output(1, 3) <= input(4);
output(1, 4) <= input(5);
output(1, 5) <= input(6);
output(1, 6) <= input(7);
output(1, 7) <= input(8);
output(1, 8) <= input(9);
output(1, 9) <= input(10);
output(1, 10) <= input(11);
output(1, 11) <= input(12);
output(1, 12) <= input(13);
output(1, 13) <= input(14);
output(1, 14) <= input(15);
output(1, 15) <= input(32);
output(1, 16) <= input(17);
output(1, 17) <= input(18);
output(1, 18) <= input(19);
output(1, 19) <= input(20);
output(1, 20) <= input(21);
output(1, 21) <= input(22);
output(1, 22) <= input(23);
output(1, 23) <= input(24);
output(1, 24) <= input(25);
output(1, 25) <= input(26);
output(1, 26) <= input(27);
output(1, 27) <= input(28);
output(1, 28) <= input(29);
output(1, 29) <= input(30);
output(1, 30) <= input(31);
output(1, 31) <= input(33);
output(1, 32) <= input(2);
output(1, 33) <= input(3);
output(1, 34) <= input(4);
output(1, 35) <= input(5);
output(1, 36) <= input(6);
output(1, 37) <= input(7);
output(1, 38) <= input(8);
output(1, 39) <= input(9);
output(1, 40) <= input(10);
output(1, 41) <= input(11);
output(1, 42) <= input(12);
output(1, 43) <= input(13);
output(1, 44) <= input(14);
output(1, 45) <= input(15);
output(1, 46) <= input(32);
output(1, 47) <= input(34);
output(1, 48) <= input(3);
output(1, 49) <= input(4);
output(1, 50) <= input(5);
output(1, 51) <= input(6);
output(1, 52) <= input(7);
output(1, 53) <= input(8);
output(1, 54) <= input(9);
output(1, 55) <= input(10);
output(1, 56) <= input(11);
output(1, 57) <= input(12);
output(1, 58) <= input(13);
output(1, 59) <= input(14);
output(1, 60) <= input(15);
output(1, 61) <= input(32);
output(1, 62) <= input(34);
output(1, 63) <= input(36);
output(1, 64) <= input(19);
output(1, 65) <= input(20);
output(1, 66) <= input(21);
output(1, 67) <= input(22);
output(1, 68) <= input(23);
output(1, 69) <= input(24);
output(1, 70) <= input(25);
output(1, 71) <= input(26);
output(1, 72) <= input(27);
output(1, 73) <= input(28);
output(1, 74) <= input(29);
output(1, 75) <= input(30);
output(1, 76) <= input(31);
output(1, 77) <= input(33);
output(1, 78) <= input(35);
output(1, 79) <= input(38);
output(1, 80) <= input(4);
output(1, 81) <= input(5);
output(1, 82) <= input(6);
output(1, 83) <= input(7);
output(1, 84) <= input(8);
output(1, 85) <= input(9);
output(1, 86) <= input(10);
output(1, 87) <= input(11);
output(1, 88) <= input(12);
output(1, 89) <= input(13);
output(1, 90) <= input(14);
output(1, 91) <= input(15);
output(1, 92) <= input(32);
output(1, 93) <= input(34);
output(1, 94) <= input(36);
output(1, 95) <= input(37);
output(1, 96) <= input(20);
output(1, 97) <= input(21);
output(1, 98) <= input(22);
output(1, 99) <= input(23);
output(1, 100) <= input(24);
output(1, 101) <= input(25);
output(1, 102) <= input(26);
output(1, 103) <= input(27);
output(1, 104) <= input(28);
output(1, 105) <= input(29);
output(1, 106) <= input(30);
output(1, 107) <= input(31);
output(1, 108) <= input(33);
output(1, 109) <= input(35);
output(1, 110) <= input(38);
output(1, 111) <= input(39);
output(1, 112) <= input(21);
output(1, 113) <= input(22);
output(1, 114) <= input(23);
output(1, 115) <= input(24);
output(1, 116) <= input(25);
output(1, 117) <= input(26);
output(1, 118) <= input(27);
output(1, 119) <= input(28);
output(1, 120) <= input(29);
output(1, 121) <= input(30);
output(1, 122) <= input(31);
output(1, 123) <= input(33);
output(1, 124) <= input(35);
output(1, 125) <= input(38);
output(1, 126) <= input(39);
output(1, 127) <= input(41);
output(1, 128) <= input(6);
output(1, 129) <= input(7);
output(1, 130) <= input(8);
output(1, 131) <= input(9);
output(1, 132) <= input(10);
output(1, 133) <= input(11);
output(1, 134) <= input(12);
output(1, 135) <= input(13);
output(1, 136) <= input(14);
output(1, 137) <= input(15);
output(1, 138) <= input(32);
output(1, 139) <= input(34);
output(1, 140) <= input(36);
output(1, 141) <= input(37);
output(1, 142) <= input(40);
output(1, 143) <= input(42);
output(1, 144) <= input(22);
output(1, 145) <= input(23);
output(1, 146) <= input(24);
output(1, 147) <= input(25);
output(1, 148) <= input(26);
output(1, 149) <= input(27);
output(1, 150) <= input(28);
output(1, 151) <= input(29);
output(1, 152) <= input(30);
output(1, 153) <= input(31);
output(1, 154) <= input(33);
output(1, 155) <= input(35);
output(1, 156) <= input(38);
output(1, 157) <= input(39);
output(1, 158) <= input(41);
output(1, 159) <= input(43);
output(1, 160) <= input(7);
output(1, 161) <= input(8);
output(1, 162) <= input(9);
output(1, 163) <= input(10);
output(1, 164) <= input(11);
output(1, 165) <= input(12);
output(1, 166) <= input(13);
output(1, 167) <= input(14);
output(1, 168) <= input(15);
output(1, 169) <= input(32);
output(1, 170) <= input(34);
output(1, 171) <= input(36);
output(1, 172) <= input(37);
output(1, 173) <= input(40);
output(1, 174) <= input(42);
output(1, 175) <= input(44);
output(1, 176) <= input(8);
output(1, 177) <= input(9);
output(1, 178) <= input(10);
output(1, 179) <= input(11);
output(1, 180) <= input(12);
output(1, 181) <= input(13);
output(1, 182) <= input(14);
output(1, 183) <= input(15);
output(1, 184) <= input(32);
output(1, 185) <= input(34);
output(1, 186) <= input(36);
output(1, 187) <= input(37);
output(1, 188) <= input(40);
output(1, 189) <= input(42);
output(1, 190) <= input(44);
output(1, 191) <= input(47);
output(1, 192) <= input(24);
output(1, 193) <= input(25);
output(1, 194) <= input(26);
output(1, 195) <= input(27);
output(1, 196) <= input(28);
output(1, 197) <= input(29);
output(1, 198) <= input(30);
output(1, 199) <= input(31);
output(1, 200) <= input(33);
output(1, 201) <= input(35);
output(1, 202) <= input(38);
output(1, 203) <= input(39);
output(1, 204) <= input(41);
output(1, 205) <= input(43);
output(1, 206) <= input(45);
output(1, 207) <= input(46);
output(1, 208) <= input(9);
output(1, 209) <= input(10);
output(1, 210) <= input(11);
output(1, 211) <= input(12);
output(1, 212) <= input(13);
output(1, 213) <= input(14);
output(1, 214) <= input(15);
output(1, 215) <= input(32);
output(1, 216) <= input(34);
output(1, 217) <= input(36);
output(1, 218) <= input(37);
output(1, 219) <= input(40);
output(1, 220) <= input(42);
output(1, 221) <= input(44);
output(1, 222) <= input(47);
output(1, 223) <= input(48);
output(1, 224) <= input(25);
output(1, 225) <= input(26);
output(1, 226) <= input(27);
output(1, 227) <= input(28);
output(1, 228) <= input(29);
output(1, 229) <= input(30);
output(1, 230) <= input(31);
output(1, 231) <= input(33);
output(1, 232) <= input(35);
output(1, 233) <= input(38);
output(1, 234) <= input(39);
output(1, 235) <= input(41);
output(1, 236) <= input(43);
output(1, 237) <= input(45);
output(1, 238) <= input(46);
output(1, 239) <= input(49);
output(1, 240) <= input(26);
output(1, 241) <= input(27);
output(1, 242) <= input(28);
output(1, 243) <= input(29);
output(1, 244) <= input(30);
output(1, 245) <= input(31);
output(1, 246) <= input(33);
output(1, 247) <= input(35);
output(1, 248) <= input(38);
output(1, 249) <= input(39);
output(1, 250) <= input(41);
output(1, 251) <= input(43);
output(1, 252) <= input(45);
output(1, 253) <= input(46);
output(1, 254) <= input(49);
output(1, 255) <= input(50);
output(2, 0) <= input(18);
output(2, 1) <= input(19);
output(2, 2) <= input(20);
output(2, 3) <= input(21);
output(2, 4) <= input(22);
output(2, 5) <= input(23);
output(2, 6) <= input(24);
output(2, 7) <= input(25);
output(2, 8) <= input(26);
output(2, 9) <= input(27);
output(2, 10) <= input(28);
output(2, 11) <= input(29);
output(2, 12) <= input(30);
output(2, 13) <= input(31);
output(2, 14) <= input(33);
output(2, 15) <= input(35);
output(2, 16) <= input(3);
output(2, 17) <= input(4);
output(2, 18) <= input(5);
output(2, 19) <= input(6);
output(2, 20) <= input(7);
output(2, 21) <= input(8);
output(2, 22) <= input(9);
output(2, 23) <= input(10);
output(2, 24) <= input(11);
output(2, 25) <= input(12);
output(2, 26) <= input(13);
output(2, 27) <= input(14);
output(2, 28) <= input(15);
output(2, 29) <= input(32);
output(2, 30) <= input(34);
output(2, 31) <= input(36);
output(2, 32) <= input(4);
output(2, 33) <= input(5);
output(2, 34) <= input(6);
output(2, 35) <= input(7);
output(2, 36) <= input(8);
output(2, 37) <= input(9);
output(2, 38) <= input(10);
output(2, 39) <= input(11);
output(2, 40) <= input(12);
output(2, 41) <= input(13);
output(2, 42) <= input(14);
output(2, 43) <= input(15);
output(2, 44) <= input(32);
output(2, 45) <= input(34);
output(2, 46) <= input(36);
output(2, 47) <= input(37);
output(2, 48) <= input(20);
output(2, 49) <= input(21);
output(2, 50) <= input(22);
output(2, 51) <= input(23);
output(2, 52) <= input(24);
output(2, 53) <= input(25);
output(2, 54) <= input(26);
output(2, 55) <= input(27);
output(2, 56) <= input(28);
output(2, 57) <= input(29);
output(2, 58) <= input(30);
output(2, 59) <= input(31);
output(2, 60) <= input(33);
output(2, 61) <= input(35);
output(2, 62) <= input(38);
output(2, 63) <= input(39);
output(2, 64) <= input(21);
output(2, 65) <= input(22);
output(2, 66) <= input(23);
output(2, 67) <= input(24);
output(2, 68) <= input(25);
output(2, 69) <= input(26);
output(2, 70) <= input(27);
output(2, 71) <= input(28);
output(2, 72) <= input(29);
output(2, 73) <= input(30);
output(2, 74) <= input(31);
output(2, 75) <= input(33);
output(2, 76) <= input(35);
output(2, 77) <= input(38);
output(2, 78) <= input(39);
output(2, 79) <= input(41);
output(2, 80) <= input(6);
output(2, 81) <= input(7);
output(2, 82) <= input(8);
output(2, 83) <= input(9);
output(2, 84) <= input(10);
output(2, 85) <= input(11);
output(2, 86) <= input(12);
output(2, 87) <= input(13);
output(2, 88) <= input(14);
output(2, 89) <= input(15);
output(2, 90) <= input(32);
output(2, 91) <= input(34);
output(2, 92) <= input(36);
output(2, 93) <= input(37);
output(2, 94) <= input(40);
output(2, 95) <= input(42);
output(2, 96) <= input(7);
output(2, 97) <= input(8);
output(2, 98) <= input(9);
output(2, 99) <= input(10);
output(2, 100) <= input(11);
output(2, 101) <= input(12);
output(2, 102) <= input(13);
output(2, 103) <= input(14);
output(2, 104) <= input(15);
output(2, 105) <= input(32);
output(2, 106) <= input(34);
output(2, 107) <= input(36);
output(2, 108) <= input(37);
output(2, 109) <= input(40);
output(2, 110) <= input(42);
output(2, 111) <= input(44);
output(2, 112) <= input(23);
output(2, 113) <= input(24);
output(2, 114) <= input(25);
output(2, 115) <= input(26);
output(2, 116) <= input(27);
output(2, 117) <= input(28);
output(2, 118) <= input(29);
output(2, 119) <= input(30);
output(2, 120) <= input(31);
output(2, 121) <= input(33);
output(2, 122) <= input(35);
output(2, 123) <= input(38);
output(2, 124) <= input(39);
output(2, 125) <= input(41);
output(2, 126) <= input(43);
output(2, 127) <= input(45);
output(2, 128) <= input(8);
output(2, 129) <= input(9);
output(2, 130) <= input(10);
output(2, 131) <= input(11);
output(2, 132) <= input(12);
output(2, 133) <= input(13);
output(2, 134) <= input(14);
output(2, 135) <= input(15);
output(2, 136) <= input(32);
output(2, 137) <= input(34);
output(2, 138) <= input(36);
output(2, 139) <= input(37);
output(2, 140) <= input(40);
output(2, 141) <= input(42);
output(2, 142) <= input(44);
output(2, 143) <= input(47);
output(2, 144) <= input(9);
output(2, 145) <= input(10);
output(2, 146) <= input(11);
output(2, 147) <= input(12);
output(2, 148) <= input(13);
output(2, 149) <= input(14);
output(2, 150) <= input(15);
output(2, 151) <= input(32);
output(2, 152) <= input(34);
output(2, 153) <= input(36);
output(2, 154) <= input(37);
output(2, 155) <= input(40);
output(2, 156) <= input(42);
output(2, 157) <= input(44);
output(2, 158) <= input(47);
output(2, 159) <= input(48);
output(2, 160) <= input(25);
output(2, 161) <= input(26);
output(2, 162) <= input(27);
output(2, 163) <= input(28);
output(2, 164) <= input(29);
output(2, 165) <= input(30);
output(2, 166) <= input(31);
output(2, 167) <= input(33);
output(2, 168) <= input(35);
output(2, 169) <= input(38);
output(2, 170) <= input(39);
output(2, 171) <= input(41);
output(2, 172) <= input(43);
output(2, 173) <= input(45);
output(2, 174) <= input(46);
output(2, 175) <= input(49);
output(2, 176) <= input(26);
output(2, 177) <= input(27);
output(2, 178) <= input(28);
output(2, 179) <= input(29);
output(2, 180) <= input(30);
output(2, 181) <= input(31);
output(2, 182) <= input(33);
output(2, 183) <= input(35);
output(2, 184) <= input(38);
output(2, 185) <= input(39);
output(2, 186) <= input(41);
output(2, 187) <= input(43);
output(2, 188) <= input(45);
output(2, 189) <= input(46);
output(2, 190) <= input(49);
output(2, 191) <= input(50);
output(2, 192) <= input(11);
output(2, 193) <= input(12);
output(2, 194) <= input(13);
output(2, 195) <= input(14);
output(2, 196) <= input(15);
output(2, 197) <= input(32);
output(2, 198) <= input(34);
output(2, 199) <= input(36);
output(2, 200) <= input(37);
output(2, 201) <= input(40);
output(2, 202) <= input(42);
output(2, 203) <= input(44);
output(2, 204) <= input(47);
output(2, 205) <= input(48);
output(2, 206) <= input(51);
output(2, 207) <= input(52);
output(2, 208) <= input(12);
output(2, 209) <= input(13);
output(2, 210) <= input(14);
output(2, 211) <= input(15);
output(2, 212) <= input(32);
output(2, 213) <= input(34);
output(2, 214) <= input(36);
output(2, 215) <= input(37);
output(2, 216) <= input(40);
output(2, 217) <= input(42);
output(2, 218) <= input(44);
output(2, 219) <= input(47);
output(2, 220) <= input(48);
output(2, 221) <= input(51);
output(2, 222) <= input(52);
output(2, 223) <= input(53);
output(2, 224) <= input(28);
output(2, 225) <= input(29);
output(2, 226) <= input(30);
output(2, 227) <= input(31);
output(2, 228) <= input(33);
output(2, 229) <= input(35);
output(2, 230) <= input(38);
output(2, 231) <= input(39);
output(2, 232) <= input(41);
output(2, 233) <= input(43);
output(2, 234) <= input(45);
output(2, 235) <= input(46);
output(2, 236) <= input(49);
output(2, 237) <= input(50);
output(2, 238) <= input(54);
output(2, 239) <= input(55);
output(2, 240) <= input(29);
output(2, 241) <= input(30);
output(2, 242) <= input(31);
output(2, 243) <= input(33);
output(2, 244) <= input(35);
output(2, 245) <= input(38);
output(2, 246) <= input(39);
output(2, 247) <= input(41);
output(2, 248) <= input(43);
output(2, 249) <= input(45);
output(2, 250) <= input(46);
output(2, 251) <= input(49);
output(2, 252) <= input(50);
output(2, 253) <= input(54);
output(2, 254) <= input(55);
output(2, 255) <= input(56);
output(3, 0) <= input(4);
output(3, 1) <= input(5);
output(3, 2) <= input(6);
output(3, 3) <= input(7);
output(3, 4) <= input(8);
output(3, 5) <= input(9);
output(3, 6) <= input(10);
output(3, 7) <= input(11);
output(3, 8) <= input(12);
output(3, 9) <= input(13);
output(3, 10) <= input(14);
output(3, 11) <= input(15);
output(3, 12) <= input(32);
output(3, 13) <= input(34);
output(3, 14) <= input(36);
output(3, 15) <= input(37);
output(3, 16) <= input(5);
output(3, 17) <= input(6);
output(3, 18) <= input(7);
output(3, 19) <= input(8);
output(3, 20) <= input(9);
output(3, 21) <= input(10);
output(3, 22) <= input(11);
output(3, 23) <= input(12);
output(3, 24) <= input(13);
output(3, 25) <= input(14);
output(3, 26) <= input(15);
output(3, 27) <= input(32);
output(3, 28) <= input(34);
output(3, 29) <= input(36);
output(3, 30) <= input(37);
output(3, 31) <= input(40);
output(3, 32) <= input(21);
output(3, 33) <= input(22);
output(3, 34) <= input(23);
output(3, 35) <= input(24);
output(3, 36) <= input(25);
output(3, 37) <= input(26);
output(3, 38) <= input(27);
output(3, 39) <= input(28);
output(3, 40) <= input(29);
output(3, 41) <= input(30);
output(3, 42) <= input(31);
output(3, 43) <= input(33);
output(3, 44) <= input(35);
output(3, 45) <= input(38);
output(3, 46) <= input(39);
output(3, 47) <= input(41);
output(3, 48) <= input(22);
output(3, 49) <= input(23);
output(3, 50) <= input(24);
output(3, 51) <= input(25);
output(3, 52) <= input(26);
output(3, 53) <= input(27);
output(3, 54) <= input(28);
output(3, 55) <= input(29);
output(3, 56) <= input(30);
output(3, 57) <= input(31);
output(3, 58) <= input(33);
output(3, 59) <= input(35);
output(3, 60) <= input(38);
output(3, 61) <= input(39);
output(3, 62) <= input(41);
output(3, 63) <= input(43);
output(3, 64) <= input(23);
output(3, 65) <= input(24);
output(3, 66) <= input(25);
output(3, 67) <= input(26);
output(3, 68) <= input(27);
output(3, 69) <= input(28);
output(3, 70) <= input(29);
output(3, 71) <= input(30);
output(3, 72) <= input(31);
output(3, 73) <= input(33);
output(3, 74) <= input(35);
output(3, 75) <= input(38);
output(3, 76) <= input(39);
output(3, 77) <= input(41);
output(3, 78) <= input(43);
output(3, 79) <= input(45);
output(3, 80) <= input(8);
output(3, 81) <= input(9);
output(3, 82) <= input(10);
output(3, 83) <= input(11);
output(3, 84) <= input(12);
output(3, 85) <= input(13);
output(3, 86) <= input(14);
output(3, 87) <= input(15);
output(3, 88) <= input(32);
output(3, 89) <= input(34);
output(3, 90) <= input(36);
output(3, 91) <= input(37);
output(3, 92) <= input(40);
output(3, 93) <= input(42);
output(3, 94) <= input(44);
output(3, 95) <= input(47);
output(3, 96) <= input(9);
output(3, 97) <= input(10);
output(3, 98) <= input(11);
output(3, 99) <= input(12);
output(3, 100) <= input(13);
output(3, 101) <= input(14);
output(3, 102) <= input(15);
output(3, 103) <= input(32);
output(3, 104) <= input(34);
output(3, 105) <= input(36);
output(3, 106) <= input(37);
output(3, 107) <= input(40);
output(3, 108) <= input(42);
output(3, 109) <= input(44);
output(3, 110) <= input(47);
output(3, 111) <= input(48);
output(3, 112) <= input(10);
output(3, 113) <= input(11);
output(3, 114) <= input(12);
output(3, 115) <= input(13);
output(3, 116) <= input(14);
output(3, 117) <= input(15);
output(3, 118) <= input(32);
output(3, 119) <= input(34);
output(3, 120) <= input(36);
output(3, 121) <= input(37);
output(3, 122) <= input(40);
output(3, 123) <= input(42);
output(3, 124) <= input(44);
output(3, 125) <= input(47);
output(3, 126) <= input(48);
output(3, 127) <= input(51);
output(3, 128) <= input(26);
output(3, 129) <= input(27);
output(3, 130) <= input(28);
output(3, 131) <= input(29);
output(3, 132) <= input(30);
output(3, 133) <= input(31);
output(3, 134) <= input(33);
output(3, 135) <= input(35);
output(3, 136) <= input(38);
output(3, 137) <= input(39);
output(3, 138) <= input(41);
output(3, 139) <= input(43);
output(3, 140) <= input(45);
output(3, 141) <= input(46);
output(3, 142) <= input(49);
output(3, 143) <= input(50);
output(3, 144) <= input(27);
output(3, 145) <= input(28);
output(3, 146) <= input(29);
output(3, 147) <= input(30);
output(3, 148) <= input(31);
output(3, 149) <= input(33);
output(3, 150) <= input(35);
output(3, 151) <= input(38);
output(3, 152) <= input(39);
output(3, 153) <= input(41);
output(3, 154) <= input(43);
output(3, 155) <= input(45);
output(3, 156) <= input(46);
output(3, 157) <= input(49);
output(3, 158) <= input(50);
output(3, 159) <= input(54);
output(3, 160) <= input(12);
output(3, 161) <= input(13);
output(3, 162) <= input(14);
output(3, 163) <= input(15);
output(3, 164) <= input(32);
output(3, 165) <= input(34);
output(3, 166) <= input(36);
output(3, 167) <= input(37);
output(3, 168) <= input(40);
output(3, 169) <= input(42);
output(3, 170) <= input(44);
output(3, 171) <= input(47);
output(3, 172) <= input(48);
output(3, 173) <= input(51);
output(3, 174) <= input(52);
output(3, 175) <= input(53);
output(3, 176) <= input(13);
output(3, 177) <= input(14);
output(3, 178) <= input(15);
output(3, 179) <= input(32);
output(3, 180) <= input(34);
output(3, 181) <= input(36);
output(3, 182) <= input(37);
output(3, 183) <= input(40);
output(3, 184) <= input(42);
output(3, 185) <= input(44);
output(3, 186) <= input(47);
output(3, 187) <= input(48);
output(3, 188) <= input(51);
output(3, 189) <= input(52);
output(3, 190) <= input(53);
output(3, 191) <= input(57);
output(3, 192) <= input(14);
output(3, 193) <= input(15);
output(3, 194) <= input(32);
output(3, 195) <= input(34);
output(3, 196) <= input(36);
output(3, 197) <= input(37);
output(3, 198) <= input(40);
output(3, 199) <= input(42);
output(3, 200) <= input(44);
output(3, 201) <= input(47);
output(3, 202) <= input(48);
output(3, 203) <= input(51);
output(3, 204) <= input(52);
output(3, 205) <= input(53);
output(3, 206) <= input(57);
output(3, 207) <= input(58);
output(3, 208) <= input(30);
output(3, 209) <= input(31);
output(3, 210) <= input(33);
output(3, 211) <= input(35);
output(3, 212) <= input(38);
output(3, 213) <= input(39);
output(3, 214) <= input(41);
output(3, 215) <= input(43);
output(3, 216) <= input(45);
output(3, 217) <= input(46);
output(3, 218) <= input(49);
output(3, 219) <= input(50);
output(3, 220) <= input(54);
output(3, 221) <= input(55);
output(3, 222) <= input(56);
output(3, 223) <= input(59);
output(3, 224) <= input(31);
output(3, 225) <= input(33);
output(3, 226) <= input(35);
output(3, 227) <= input(38);
output(3, 228) <= input(39);
output(3, 229) <= input(41);
output(3, 230) <= input(43);
output(3, 231) <= input(45);
output(3, 232) <= input(46);
output(3, 233) <= input(49);
output(3, 234) <= input(50);
output(3, 235) <= input(54);
output(3, 236) <= input(55);
output(3, 237) <= input(56);
output(3, 238) <= input(59);
output(3, 239) <= input(60);
output(3, 240) <= input(33);
output(3, 241) <= input(35);
output(3, 242) <= input(38);
output(3, 243) <= input(39);
output(3, 244) <= input(41);
output(3, 245) <= input(43);
output(3, 246) <= input(45);
output(3, 247) <= input(46);
output(3, 248) <= input(49);
output(3, 249) <= input(50);
output(3, 250) <= input(54);
output(3, 251) <= input(55);
output(3, 252) <= input(56);
output(3, 253) <= input(59);
output(3, 254) <= input(60);
output(3, 255) <= input(61);
output(4, 0) <= input(21);
output(4, 1) <= input(22);
output(4, 2) <= input(23);
output(4, 3) <= input(24);
output(4, 4) <= input(25);
output(4, 5) <= input(26);
output(4, 6) <= input(27);
output(4, 7) <= input(28);
output(4, 8) <= input(29);
output(4, 9) <= input(30);
output(4, 10) <= input(31);
output(4, 11) <= input(33);
output(4, 12) <= input(35);
output(4, 13) <= input(38);
output(4, 14) <= input(39);
output(4, 15) <= input(41);
output(4, 16) <= input(22);
output(4, 17) <= input(23);
output(4, 18) <= input(24);
output(4, 19) <= input(25);
output(4, 20) <= input(26);
output(4, 21) <= input(27);
output(4, 22) <= input(28);
output(4, 23) <= input(29);
output(4, 24) <= input(30);
output(4, 25) <= input(31);
output(4, 26) <= input(33);
output(4, 27) <= input(35);
output(4, 28) <= input(38);
output(4, 29) <= input(39);
output(4, 30) <= input(41);
output(4, 31) <= input(43);
output(4, 32) <= input(23);
output(4, 33) <= input(24);
output(4, 34) <= input(25);
output(4, 35) <= input(26);
output(4, 36) <= input(27);
output(4, 37) <= input(28);
output(4, 38) <= input(29);
output(4, 39) <= input(30);
output(4, 40) <= input(31);
output(4, 41) <= input(33);
output(4, 42) <= input(35);
output(4, 43) <= input(38);
output(4, 44) <= input(39);
output(4, 45) <= input(41);
output(4, 46) <= input(43);
output(4, 47) <= input(45);
output(4, 48) <= input(24);
output(4, 49) <= input(25);
output(4, 50) <= input(26);
output(4, 51) <= input(27);
output(4, 52) <= input(28);
output(4, 53) <= input(29);
output(4, 54) <= input(30);
output(4, 55) <= input(31);
output(4, 56) <= input(33);
output(4, 57) <= input(35);
output(4, 58) <= input(38);
output(4, 59) <= input(39);
output(4, 60) <= input(41);
output(4, 61) <= input(43);
output(4, 62) <= input(45);
output(4, 63) <= input(46);
output(4, 64) <= input(25);
output(4, 65) <= input(26);
output(4, 66) <= input(27);
output(4, 67) <= input(28);
output(4, 68) <= input(29);
output(4, 69) <= input(30);
output(4, 70) <= input(31);
output(4, 71) <= input(33);
output(4, 72) <= input(35);
output(4, 73) <= input(38);
output(4, 74) <= input(39);
output(4, 75) <= input(41);
output(4, 76) <= input(43);
output(4, 77) <= input(45);
output(4, 78) <= input(46);
output(4, 79) <= input(49);
output(4, 80) <= input(10);
output(4, 81) <= input(11);
output(4, 82) <= input(12);
output(4, 83) <= input(13);
output(4, 84) <= input(14);
output(4, 85) <= input(15);
output(4, 86) <= input(32);
output(4, 87) <= input(34);
output(4, 88) <= input(36);
output(4, 89) <= input(37);
output(4, 90) <= input(40);
output(4, 91) <= input(42);
output(4, 92) <= input(44);
output(4, 93) <= input(47);
output(4, 94) <= input(48);
output(4, 95) <= input(51);
output(4, 96) <= input(11);
output(4, 97) <= input(12);
output(4, 98) <= input(13);
output(4, 99) <= input(14);
output(4, 100) <= input(15);
output(4, 101) <= input(32);
output(4, 102) <= input(34);
output(4, 103) <= input(36);
output(4, 104) <= input(37);
output(4, 105) <= input(40);
output(4, 106) <= input(42);
output(4, 107) <= input(44);
output(4, 108) <= input(47);
output(4, 109) <= input(48);
output(4, 110) <= input(51);
output(4, 111) <= input(52);
output(4, 112) <= input(12);
output(4, 113) <= input(13);
output(4, 114) <= input(14);
output(4, 115) <= input(15);
output(4, 116) <= input(32);
output(4, 117) <= input(34);
output(4, 118) <= input(36);
output(4, 119) <= input(37);
output(4, 120) <= input(40);
output(4, 121) <= input(42);
output(4, 122) <= input(44);
output(4, 123) <= input(47);
output(4, 124) <= input(48);
output(4, 125) <= input(51);
output(4, 126) <= input(52);
output(4, 127) <= input(53);
output(4, 128) <= input(13);
output(4, 129) <= input(14);
output(4, 130) <= input(15);
output(4, 131) <= input(32);
output(4, 132) <= input(34);
output(4, 133) <= input(36);
output(4, 134) <= input(37);
output(4, 135) <= input(40);
output(4, 136) <= input(42);
output(4, 137) <= input(44);
output(4, 138) <= input(47);
output(4, 139) <= input(48);
output(4, 140) <= input(51);
output(4, 141) <= input(52);
output(4, 142) <= input(53);
output(4, 143) <= input(57);
output(4, 144) <= input(14);
output(4, 145) <= input(15);
output(4, 146) <= input(32);
output(4, 147) <= input(34);
output(4, 148) <= input(36);
output(4, 149) <= input(37);
output(4, 150) <= input(40);
output(4, 151) <= input(42);
output(4, 152) <= input(44);
output(4, 153) <= input(47);
output(4, 154) <= input(48);
output(4, 155) <= input(51);
output(4, 156) <= input(52);
output(4, 157) <= input(53);
output(4, 158) <= input(57);
output(4, 159) <= input(58);
output(4, 160) <= input(30);
output(4, 161) <= input(31);
output(4, 162) <= input(33);
output(4, 163) <= input(35);
output(4, 164) <= input(38);
output(4, 165) <= input(39);
output(4, 166) <= input(41);
output(4, 167) <= input(43);
output(4, 168) <= input(45);
output(4, 169) <= input(46);
output(4, 170) <= input(49);
output(4, 171) <= input(50);
output(4, 172) <= input(54);
output(4, 173) <= input(55);
output(4, 174) <= input(56);
output(4, 175) <= input(59);
output(4, 176) <= input(31);
output(4, 177) <= input(33);
output(4, 178) <= input(35);
output(4, 179) <= input(38);
output(4, 180) <= input(39);
output(4, 181) <= input(41);
output(4, 182) <= input(43);
output(4, 183) <= input(45);
output(4, 184) <= input(46);
output(4, 185) <= input(49);
output(4, 186) <= input(50);
output(4, 187) <= input(54);
output(4, 188) <= input(55);
output(4, 189) <= input(56);
output(4, 190) <= input(59);
output(4, 191) <= input(60);
output(4, 192) <= input(33);
output(4, 193) <= input(35);
output(4, 194) <= input(38);
output(4, 195) <= input(39);
output(4, 196) <= input(41);
output(4, 197) <= input(43);
output(4, 198) <= input(45);
output(4, 199) <= input(46);
output(4, 200) <= input(49);
output(4, 201) <= input(50);
output(4, 202) <= input(54);
output(4, 203) <= input(55);
output(4, 204) <= input(56);
output(4, 205) <= input(59);
output(4, 206) <= input(60);
output(4, 207) <= input(61);
output(4, 208) <= input(35);
output(4, 209) <= input(38);
output(4, 210) <= input(39);
output(4, 211) <= input(41);
output(4, 212) <= input(43);
output(4, 213) <= input(45);
output(4, 214) <= input(46);
output(4, 215) <= input(49);
output(4, 216) <= input(50);
output(4, 217) <= input(54);
output(4, 218) <= input(55);
output(4, 219) <= input(56);
output(4, 220) <= input(59);
output(4, 221) <= input(60);
output(4, 222) <= input(61);
output(4, 223) <= input(62);
output(4, 224) <= input(38);
output(4, 225) <= input(39);
output(4, 226) <= input(41);
output(4, 227) <= input(43);
output(4, 228) <= input(45);
output(4, 229) <= input(46);
output(4, 230) <= input(49);
output(4, 231) <= input(50);
output(4, 232) <= input(54);
output(4, 233) <= input(55);
output(4, 234) <= input(56);
output(4, 235) <= input(59);
output(4, 236) <= input(60);
output(4, 237) <= input(61);
output(4, 238) <= input(62);
output(4, 239) <= input(63);
output(4, 240) <= input(39);
output(4, 241) <= input(41);
output(4, 242) <= input(43);
output(4, 243) <= input(45);
output(4, 244) <= input(46);
output(4, 245) <= input(49);
output(4, 246) <= input(50);
output(4, 247) <= input(54);
output(4, 248) <= input(55);
output(4, 249) <= input(56);
output(4, 250) <= input(59);
output(4, 251) <= input(60);
output(4, 252) <= input(61);
output(4, 253) <= input(62);
output(4, 254) <= input(63);
output(4, 255) <= input(64);
output(5, 0) <= input(23);
output(5, 1) <= input(24);
output(5, 2) <= input(25);
output(5, 3) <= input(26);
output(5, 4) <= input(27);
output(5, 5) <= input(28);
output(5, 6) <= input(29);
output(5, 7) <= input(30);
output(5, 8) <= input(31);
output(5, 9) <= input(33);
output(5, 10) <= input(35);
output(5, 11) <= input(38);
output(5, 12) <= input(39);
output(5, 13) <= input(41);
output(5, 14) <= input(43);
output(5, 15) <= input(45);
output(5, 16) <= input(24);
output(5, 17) <= input(25);
output(5, 18) <= input(26);
output(5, 19) <= input(27);
output(5, 20) <= input(28);
output(5, 21) <= input(29);
output(5, 22) <= input(30);
output(5, 23) <= input(31);
output(5, 24) <= input(33);
output(5, 25) <= input(35);
output(5, 26) <= input(38);
output(5, 27) <= input(39);
output(5, 28) <= input(41);
output(5, 29) <= input(43);
output(5, 30) <= input(45);
output(5, 31) <= input(46);
output(5, 32) <= input(25);
output(5, 33) <= input(26);
output(5, 34) <= input(27);
output(5, 35) <= input(28);
output(5, 36) <= input(29);
output(5, 37) <= input(30);
output(5, 38) <= input(31);
output(5, 39) <= input(33);
output(5, 40) <= input(35);
output(5, 41) <= input(38);
output(5, 42) <= input(39);
output(5, 43) <= input(41);
output(5, 44) <= input(43);
output(5, 45) <= input(45);
output(5, 46) <= input(46);
output(5, 47) <= input(49);
output(5, 48) <= input(26);
output(5, 49) <= input(27);
output(5, 50) <= input(28);
output(5, 51) <= input(29);
output(5, 52) <= input(30);
output(5, 53) <= input(31);
output(5, 54) <= input(33);
output(5, 55) <= input(35);
output(5, 56) <= input(38);
output(5, 57) <= input(39);
output(5, 58) <= input(41);
output(5, 59) <= input(43);
output(5, 60) <= input(45);
output(5, 61) <= input(46);
output(5, 62) <= input(49);
output(5, 63) <= input(50);
output(5, 64) <= input(27);
output(5, 65) <= input(28);
output(5, 66) <= input(29);
output(5, 67) <= input(30);
output(5, 68) <= input(31);
output(5, 69) <= input(33);
output(5, 70) <= input(35);
output(5, 71) <= input(38);
output(5, 72) <= input(39);
output(5, 73) <= input(41);
output(5, 74) <= input(43);
output(5, 75) <= input(45);
output(5, 76) <= input(46);
output(5, 77) <= input(49);
output(5, 78) <= input(50);
output(5, 79) <= input(54);
output(5, 80) <= input(28);
output(5, 81) <= input(29);
output(5, 82) <= input(30);
output(5, 83) <= input(31);
output(5, 84) <= input(33);
output(5, 85) <= input(35);
output(5, 86) <= input(38);
output(5, 87) <= input(39);
output(5, 88) <= input(41);
output(5, 89) <= input(43);
output(5, 90) <= input(45);
output(5, 91) <= input(46);
output(5, 92) <= input(49);
output(5, 93) <= input(50);
output(5, 94) <= input(54);
output(5, 95) <= input(55);
output(5, 96) <= input(29);
output(5, 97) <= input(30);
output(5, 98) <= input(31);
output(5, 99) <= input(33);
output(5, 100) <= input(35);
output(5, 101) <= input(38);
output(5, 102) <= input(39);
output(5, 103) <= input(41);
output(5, 104) <= input(43);
output(5, 105) <= input(45);
output(5, 106) <= input(46);
output(5, 107) <= input(49);
output(5, 108) <= input(50);
output(5, 109) <= input(54);
output(5, 110) <= input(55);
output(5, 111) <= input(56);
output(5, 112) <= input(30);
output(5, 113) <= input(31);
output(5, 114) <= input(33);
output(5, 115) <= input(35);
output(5, 116) <= input(38);
output(5, 117) <= input(39);
output(5, 118) <= input(41);
output(5, 119) <= input(43);
output(5, 120) <= input(45);
output(5, 121) <= input(46);
output(5, 122) <= input(49);
output(5, 123) <= input(50);
output(5, 124) <= input(54);
output(5, 125) <= input(55);
output(5, 126) <= input(56);
output(5, 127) <= input(59);
output(5, 128) <= input(31);
output(5, 129) <= input(33);
output(5, 130) <= input(35);
output(5, 131) <= input(38);
output(5, 132) <= input(39);
output(5, 133) <= input(41);
output(5, 134) <= input(43);
output(5, 135) <= input(45);
output(5, 136) <= input(46);
output(5, 137) <= input(49);
output(5, 138) <= input(50);
output(5, 139) <= input(54);
output(5, 140) <= input(55);
output(5, 141) <= input(56);
output(5, 142) <= input(59);
output(5, 143) <= input(60);
output(5, 144) <= input(33);
output(5, 145) <= input(35);
output(5, 146) <= input(38);
output(5, 147) <= input(39);
output(5, 148) <= input(41);
output(5, 149) <= input(43);
output(5, 150) <= input(45);
output(5, 151) <= input(46);
output(5, 152) <= input(49);
output(5, 153) <= input(50);
output(5, 154) <= input(54);
output(5, 155) <= input(55);
output(5, 156) <= input(56);
output(5, 157) <= input(59);
output(5, 158) <= input(60);
output(5, 159) <= input(61);
output(5, 160) <= input(35);
output(5, 161) <= input(38);
output(5, 162) <= input(39);
output(5, 163) <= input(41);
output(5, 164) <= input(43);
output(5, 165) <= input(45);
output(5, 166) <= input(46);
output(5, 167) <= input(49);
output(5, 168) <= input(50);
output(5, 169) <= input(54);
output(5, 170) <= input(55);
output(5, 171) <= input(56);
output(5, 172) <= input(59);
output(5, 173) <= input(60);
output(5, 174) <= input(61);
output(5, 175) <= input(62);
output(5, 176) <= input(38);
output(5, 177) <= input(39);
output(5, 178) <= input(41);
output(5, 179) <= input(43);
output(5, 180) <= input(45);
output(5, 181) <= input(46);
output(5, 182) <= input(49);
output(5, 183) <= input(50);
output(5, 184) <= input(54);
output(5, 185) <= input(55);
output(5, 186) <= input(56);
output(5, 187) <= input(59);
output(5, 188) <= input(60);
output(5, 189) <= input(61);
output(5, 190) <= input(62);
output(5, 191) <= input(63);
output(5, 192) <= input(39);
output(5, 193) <= input(41);
output(5, 194) <= input(43);
output(5, 195) <= input(45);
output(5, 196) <= input(46);
output(5, 197) <= input(49);
output(5, 198) <= input(50);
output(5, 199) <= input(54);
output(5, 200) <= input(55);
output(5, 201) <= input(56);
output(5, 202) <= input(59);
output(5, 203) <= input(60);
output(5, 204) <= input(61);
output(5, 205) <= input(62);
output(5, 206) <= input(63);
output(5, 207) <= input(64);
output(5, 208) <= input(41);
output(5, 209) <= input(43);
output(5, 210) <= input(45);
output(5, 211) <= input(46);
output(5, 212) <= input(49);
output(5, 213) <= input(50);
output(5, 214) <= input(54);
output(5, 215) <= input(55);
output(5, 216) <= input(56);
output(5, 217) <= input(59);
output(5, 218) <= input(60);
output(5, 219) <= input(61);
output(5, 220) <= input(62);
output(5, 221) <= input(63);
output(5, 222) <= input(64);
output(5, 223) <= input(65);
output(5, 224) <= input(43);
output(5, 225) <= input(45);
output(5, 226) <= input(46);
output(5, 227) <= input(49);
output(5, 228) <= input(50);
output(5, 229) <= input(54);
output(5, 230) <= input(55);
output(5, 231) <= input(56);
output(5, 232) <= input(59);
output(5, 233) <= input(60);
output(5, 234) <= input(61);
output(5, 235) <= input(62);
output(5, 236) <= input(63);
output(5, 237) <= input(64);
output(5, 238) <= input(65);
output(5, 239) <= input(66);
output(5, 240) <= input(45);
output(5, 241) <= input(46);
output(5, 242) <= input(49);
output(5, 243) <= input(50);
output(5, 244) <= input(54);
output(5, 245) <= input(55);
output(5, 246) <= input(56);
output(5, 247) <= input(59);
output(5, 248) <= input(60);
output(5, 249) <= input(61);
output(5, 250) <= input(62);
output(5, 251) <= input(63);
output(5, 252) <= input(64);
output(5, 253) <= input(65);
output(5, 254) <= input(66);
output(5, 255) <= input(67);
when others => for i in 0 to 7 loop for j in 0 to 255 loop output(i,j) <= "00000000"; end loop; end loop;
end case;
elsif control = "110" then 
case iteration_control is
when "0000" =>
output(0, 0) <= input(0);
output(0, 1) <= input(1);
output(0, 2) <= input(2);
output(0, 3) <= input(3);
output(0, 4) <= input(4);
output(0, 5) <= input(5);
output(0, 6) <= input(6);
output(0, 7) <= input(7);
output(0, 8) <= input(8);
output(0, 9) <= input(9);
output(0, 10) <= input(10);
output(0, 11) <= input(11);
output(0, 12) <= input(12);
output(0, 13) <= input(13);
output(0, 14) <= input(14);
output(0, 15) <= input(15);
output(0, 16) <= input(1);
output(0, 17) <= input(2);
output(0, 18) <= input(3);
output(0, 19) <= input(4);
output(0, 20) <= input(5);
output(0, 21) <= input(6);
output(0, 22) <= input(7);
output(0, 23) <= input(8);
output(0, 24) <= input(9);
output(0, 25) <= input(10);
output(0, 26) <= input(11);
output(0, 27) <= input(12);
output(0, 28) <= input(13);
output(0, 29) <= input(14);
output(0, 30) <= input(15);
output(0, 31) <= input(16);
output(0, 32) <= input(2);
output(0, 33) <= input(3);
output(0, 34) <= input(4);
output(0, 35) <= input(5);
output(0, 36) <= input(6);
output(0, 37) <= input(7);
output(0, 38) <= input(8);
output(0, 39) <= input(9);
output(0, 40) <= input(10);
output(0, 41) <= input(11);
output(0, 42) <= input(12);
output(0, 43) <= input(13);
output(0, 44) <= input(14);
output(0, 45) <= input(15);
output(0, 46) <= input(16);
output(0, 47) <= input(17);
output(0, 48) <= input(3);
output(0, 49) <= input(4);
output(0, 50) <= input(5);
output(0, 51) <= input(6);
output(0, 52) <= input(7);
output(0, 53) <= input(8);
output(0, 54) <= input(9);
output(0, 55) <= input(10);
output(0, 56) <= input(11);
output(0, 57) <= input(12);
output(0, 58) <= input(13);
output(0, 59) <= input(14);
output(0, 60) <= input(15);
output(0, 61) <= input(16);
output(0, 62) <= input(17);
output(0, 63) <= input(18);
output(0, 64) <= input(4);
output(0, 65) <= input(5);
output(0, 66) <= input(6);
output(0, 67) <= input(7);
output(0, 68) <= input(8);
output(0, 69) <= input(9);
output(0, 70) <= input(10);
output(0, 71) <= input(11);
output(0, 72) <= input(12);
output(0, 73) <= input(13);
output(0, 74) <= input(14);
output(0, 75) <= input(15);
output(0, 76) <= input(16);
output(0, 77) <= input(17);
output(0, 78) <= input(18);
output(0, 79) <= input(19);
output(0, 80) <= input(5);
output(0, 81) <= input(6);
output(0, 82) <= input(7);
output(0, 83) <= input(8);
output(0, 84) <= input(9);
output(0, 85) <= input(10);
output(0, 86) <= input(11);
output(0, 87) <= input(12);
output(0, 88) <= input(13);
output(0, 89) <= input(14);
output(0, 90) <= input(15);
output(0, 91) <= input(16);
output(0, 92) <= input(17);
output(0, 93) <= input(18);
output(0, 94) <= input(19);
output(0, 95) <= input(20);
output(0, 96) <= input(6);
output(0, 97) <= input(7);
output(0, 98) <= input(8);
output(0, 99) <= input(9);
output(0, 100) <= input(10);
output(0, 101) <= input(11);
output(0, 102) <= input(12);
output(0, 103) <= input(13);
output(0, 104) <= input(14);
output(0, 105) <= input(15);
output(0, 106) <= input(16);
output(0, 107) <= input(17);
output(0, 108) <= input(18);
output(0, 109) <= input(19);
output(0, 110) <= input(20);
output(0, 111) <= input(21);
output(0, 112) <= input(7);
output(0, 113) <= input(8);
output(0, 114) <= input(9);
output(0, 115) <= input(10);
output(0, 116) <= input(11);
output(0, 117) <= input(12);
output(0, 118) <= input(13);
output(0, 119) <= input(14);
output(0, 120) <= input(15);
output(0, 121) <= input(16);
output(0, 122) <= input(17);
output(0, 123) <= input(18);
output(0, 124) <= input(19);
output(0, 125) <= input(20);
output(0, 126) <= input(21);
output(0, 127) <= input(22);
output(0, 128) <= input(8);
output(0, 129) <= input(9);
output(0, 130) <= input(10);
output(0, 131) <= input(11);
output(0, 132) <= input(12);
output(0, 133) <= input(13);
output(0, 134) <= input(14);
output(0, 135) <= input(15);
output(0, 136) <= input(16);
output(0, 137) <= input(17);
output(0, 138) <= input(18);
output(0, 139) <= input(19);
output(0, 140) <= input(20);
output(0, 141) <= input(21);
output(0, 142) <= input(22);
output(0, 143) <= input(23);
output(0, 144) <= input(9);
output(0, 145) <= input(10);
output(0, 146) <= input(11);
output(0, 147) <= input(12);
output(0, 148) <= input(13);
output(0, 149) <= input(14);
output(0, 150) <= input(15);
output(0, 151) <= input(16);
output(0, 152) <= input(17);
output(0, 153) <= input(18);
output(0, 154) <= input(19);
output(0, 155) <= input(20);
output(0, 156) <= input(21);
output(0, 157) <= input(22);
output(0, 158) <= input(23);
output(0, 159) <= input(24);
output(0, 160) <= input(10);
output(0, 161) <= input(11);
output(0, 162) <= input(12);
output(0, 163) <= input(13);
output(0, 164) <= input(14);
output(0, 165) <= input(15);
output(0, 166) <= input(16);
output(0, 167) <= input(17);
output(0, 168) <= input(18);
output(0, 169) <= input(19);
output(0, 170) <= input(20);
output(0, 171) <= input(21);
output(0, 172) <= input(22);
output(0, 173) <= input(23);
output(0, 174) <= input(24);
output(0, 175) <= input(25);
output(0, 176) <= input(11);
output(0, 177) <= input(12);
output(0, 178) <= input(13);
output(0, 179) <= input(14);
output(0, 180) <= input(15);
output(0, 181) <= input(16);
output(0, 182) <= input(17);
output(0, 183) <= input(18);
output(0, 184) <= input(19);
output(0, 185) <= input(20);
output(0, 186) <= input(21);
output(0, 187) <= input(22);
output(0, 188) <= input(23);
output(0, 189) <= input(24);
output(0, 190) <= input(25);
output(0, 191) <= input(26);
output(0, 192) <= input(12);
output(0, 193) <= input(13);
output(0, 194) <= input(14);
output(0, 195) <= input(15);
output(0, 196) <= input(16);
output(0, 197) <= input(17);
output(0, 198) <= input(18);
output(0, 199) <= input(19);
output(0, 200) <= input(20);
output(0, 201) <= input(21);
output(0, 202) <= input(22);
output(0, 203) <= input(23);
output(0, 204) <= input(24);
output(0, 205) <= input(25);
output(0, 206) <= input(26);
output(0, 207) <= input(27);
output(0, 208) <= input(13);
output(0, 209) <= input(14);
output(0, 210) <= input(15);
output(0, 211) <= input(16);
output(0, 212) <= input(17);
output(0, 213) <= input(18);
output(0, 214) <= input(19);
output(0, 215) <= input(20);
output(0, 216) <= input(21);
output(0, 217) <= input(22);
output(0, 218) <= input(23);
output(0, 219) <= input(24);
output(0, 220) <= input(25);
output(0, 221) <= input(26);
output(0, 222) <= input(27);
output(0, 223) <= input(28);
output(0, 224) <= input(14);
output(0, 225) <= input(15);
output(0, 226) <= input(16);
output(0, 227) <= input(17);
output(0, 228) <= input(18);
output(0, 229) <= input(19);
output(0, 230) <= input(20);
output(0, 231) <= input(21);
output(0, 232) <= input(22);
output(0, 233) <= input(23);
output(0, 234) <= input(24);
output(0, 235) <= input(25);
output(0, 236) <= input(26);
output(0, 237) <= input(27);
output(0, 238) <= input(28);
output(0, 239) <= input(29);
output(0, 240) <= input(15);
output(0, 241) <= input(16);
output(0, 242) <= input(17);
output(0, 243) <= input(18);
output(0, 244) <= input(19);
output(0, 245) <= input(20);
output(0, 246) <= input(21);
output(0, 247) <= input(22);
output(0, 248) <= input(23);
output(0, 249) <= input(24);
output(0, 250) <= input(25);
output(0, 251) <= input(26);
output(0, 252) <= input(27);
output(0, 253) <= input(28);
output(0, 254) <= input(29);
output(0, 255) <= input(30);
output(1, 0) <= input(31);
output(1, 1) <= input(32);
output(1, 2) <= input(0);
output(1, 3) <= input(1);
output(1, 4) <= input(2);
output(1, 5) <= input(3);
output(1, 6) <= input(4);
output(1, 7) <= input(5);
output(1, 8) <= input(6);
output(1, 9) <= input(7);
output(1, 10) <= input(8);
output(1, 11) <= input(9);
output(1, 12) <= input(10);
output(1, 13) <= input(11);
output(1, 14) <= input(12);
output(1, 15) <= input(13);
output(1, 16) <= input(32);
output(1, 17) <= input(0);
output(1, 18) <= input(1);
output(1, 19) <= input(2);
output(1, 20) <= input(3);
output(1, 21) <= input(4);
output(1, 22) <= input(5);
output(1, 23) <= input(6);
output(1, 24) <= input(7);
output(1, 25) <= input(8);
output(1, 26) <= input(9);
output(1, 27) <= input(10);
output(1, 28) <= input(11);
output(1, 29) <= input(12);
output(1, 30) <= input(13);
output(1, 31) <= input(14);
output(1, 32) <= input(0);
output(1, 33) <= input(1);
output(1, 34) <= input(2);
output(1, 35) <= input(3);
output(1, 36) <= input(4);
output(1, 37) <= input(5);
output(1, 38) <= input(6);
output(1, 39) <= input(7);
output(1, 40) <= input(8);
output(1, 41) <= input(9);
output(1, 42) <= input(10);
output(1, 43) <= input(11);
output(1, 44) <= input(12);
output(1, 45) <= input(13);
output(1, 46) <= input(14);
output(1, 47) <= input(15);
output(1, 48) <= input(1);
output(1, 49) <= input(2);
output(1, 50) <= input(3);
output(1, 51) <= input(4);
output(1, 52) <= input(5);
output(1, 53) <= input(6);
output(1, 54) <= input(7);
output(1, 55) <= input(8);
output(1, 56) <= input(9);
output(1, 57) <= input(10);
output(1, 58) <= input(11);
output(1, 59) <= input(12);
output(1, 60) <= input(13);
output(1, 61) <= input(14);
output(1, 62) <= input(15);
output(1, 63) <= input(16);
output(1, 64) <= input(2);
output(1, 65) <= input(3);
output(1, 66) <= input(4);
output(1, 67) <= input(5);
output(1, 68) <= input(6);
output(1, 69) <= input(7);
output(1, 70) <= input(8);
output(1, 71) <= input(9);
output(1, 72) <= input(10);
output(1, 73) <= input(11);
output(1, 74) <= input(12);
output(1, 75) <= input(13);
output(1, 76) <= input(14);
output(1, 77) <= input(15);
output(1, 78) <= input(16);
output(1, 79) <= input(17);
output(1, 80) <= input(33);
output(1, 81) <= input(34);
output(1, 82) <= input(35);
output(1, 83) <= input(36);
output(1, 84) <= input(37);
output(1, 85) <= input(38);
output(1, 86) <= input(39);
output(1, 87) <= input(40);
output(1, 88) <= input(41);
output(1, 89) <= input(42);
output(1, 90) <= input(43);
output(1, 91) <= input(44);
output(1, 92) <= input(45);
output(1, 93) <= input(46);
output(1, 94) <= input(47);
output(1, 95) <= input(48);
output(1, 96) <= input(34);
output(1, 97) <= input(35);
output(1, 98) <= input(36);
output(1, 99) <= input(37);
output(1, 100) <= input(38);
output(1, 101) <= input(39);
output(1, 102) <= input(40);
output(1, 103) <= input(41);
output(1, 104) <= input(42);
output(1, 105) <= input(43);
output(1, 106) <= input(44);
output(1, 107) <= input(45);
output(1, 108) <= input(46);
output(1, 109) <= input(47);
output(1, 110) <= input(48);
output(1, 111) <= input(49);
output(1, 112) <= input(35);
output(1, 113) <= input(36);
output(1, 114) <= input(37);
output(1, 115) <= input(38);
output(1, 116) <= input(39);
output(1, 117) <= input(40);
output(1, 118) <= input(41);
output(1, 119) <= input(42);
output(1, 120) <= input(43);
output(1, 121) <= input(44);
output(1, 122) <= input(45);
output(1, 123) <= input(46);
output(1, 124) <= input(47);
output(1, 125) <= input(48);
output(1, 126) <= input(49);
output(1, 127) <= input(50);
output(1, 128) <= input(36);
output(1, 129) <= input(37);
output(1, 130) <= input(38);
output(1, 131) <= input(39);
output(1, 132) <= input(40);
output(1, 133) <= input(41);
output(1, 134) <= input(42);
output(1, 135) <= input(43);
output(1, 136) <= input(44);
output(1, 137) <= input(45);
output(1, 138) <= input(46);
output(1, 139) <= input(47);
output(1, 140) <= input(48);
output(1, 141) <= input(49);
output(1, 142) <= input(50);
output(1, 143) <= input(51);
output(1, 144) <= input(37);
output(1, 145) <= input(38);
output(1, 146) <= input(39);
output(1, 147) <= input(40);
output(1, 148) <= input(41);
output(1, 149) <= input(42);
output(1, 150) <= input(43);
output(1, 151) <= input(44);
output(1, 152) <= input(45);
output(1, 153) <= input(46);
output(1, 154) <= input(47);
output(1, 155) <= input(48);
output(1, 156) <= input(49);
output(1, 157) <= input(50);
output(1, 158) <= input(51);
output(1, 159) <= input(52);
output(1, 160) <= input(7);
output(1, 161) <= input(8);
output(1, 162) <= input(9);
output(1, 163) <= input(10);
output(1, 164) <= input(11);
output(1, 165) <= input(12);
output(1, 166) <= input(13);
output(1, 167) <= input(14);
output(1, 168) <= input(15);
output(1, 169) <= input(16);
output(1, 170) <= input(17);
output(1, 171) <= input(18);
output(1, 172) <= input(19);
output(1, 173) <= input(20);
output(1, 174) <= input(21);
output(1, 175) <= input(22);
output(1, 176) <= input(8);
output(1, 177) <= input(9);
output(1, 178) <= input(10);
output(1, 179) <= input(11);
output(1, 180) <= input(12);
output(1, 181) <= input(13);
output(1, 182) <= input(14);
output(1, 183) <= input(15);
output(1, 184) <= input(16);
output(1, 185) <= input(17);
output(1, 186) <= input(18);
output(1, 187) <= input(19);
output(1, 188) <= input(20);
output(1, 189) <= input(21);
output(1, 190) <= input(22);
output(1, 191) <= input(23);
output(1, 192) <= input(9);
output(1, 193) <= input(10);
output(1, 194) <= input(11);
output(1, 195) <= input(12);
output(1, 196) <= input(13);
output(1, 197) <= input(14);
output(1, 198) <= input(15);
output(1, 199) <= input(16);
output(1, 200) <= input(17);
output(1, 201) <= input(18);
output(1, 202) <= input(19);
output(1, 203) <= input(20);
output(1, 204) <= input(21);
output(1, 205) <= input(22);
output(1, 206) <= input(23);
output(1, 207) <= input(24);
output(1, 208) <= input(10);
output(1, 209) <= input(11);
output(1, 210) <= input(12);
output(1, 211) <= input(13);
output(1, 212) <= input(14);
output(1, 213) <= input(15);
output(1, 214) <= input(16);
output(1, 215) <= input(17);
output(1, 216) <= input(18);
output(1, 217) <= input(19);
output(1, 218) <= input(20);
output(1, 219) <= input(21);
output(1, 220) <= input(22);
output(1, 221) <= input(23);
output(1, 222) <= input(24);
output(1, 223) <= input(25);
output(1, 224) <= input(11);
output(1, 225) <= input(12);
output(1, 226) <= input(13);
output(1, 227) <= input(14);
output(1, 228) <= input(15);
output(1, 229) <= input(16);
output(1, 230) <= input(17);
output(1, 231) <= input(18);
output(1, 232) <= input(19);
output(1, 233) <= input(20);
output(1, 234) <= input(21);
output(1, 235) <= input(22);
output(1, 236) <= input(23);
output(1, 237) <= input(24);
output(1, 238) <= input(25);
output(1, 239) <= input(26);
output(1, 240) <= input(12);
output(1, 241) <= input(13);
output(1, 242) <= input(14);
output(1, 243) <= input(15);
output(1, 244) <= input(16);
output(1, 245) <= input(17);
output(1, 246) <= input(18);
output(1, 247) <= input(19);
output(1, 248) <= input(20);
output(1, 249) <= input(21);
output(1, 250) <= input(22);
output(1, 251) <= input(23);
output(1, 252) <= input(24);
output(1, 253) <= input(25);
output(1, 254) <= input(26);
output(1, 255) <= input(27);
output(2, 0) <= input(53);
output(2, 1) <= input(54);
output(2, 2) <= input(55);
output(2, 3) <= input(56);
output(2, 4) <= input(57);
output(2, 5) <= input(58);
output(2, 6) <= input(33);
output(2, 7) <= input(34);
output(2, 8) <= input(35);
output(2, 9) <= input(36);
output(2, 10) <= input(37);
output(2, 11) <= input(38);
output(2, 12) <= input(39);
output(2, 13) <= input(40);
output(2, 14) <= input(41);
output(2, 15) <= input(42);
output(2, 16) <= input(54);
output(2, 17) <= input(55);
output(2, 18) <= input(56);
output(2, 19) <= input(57);
output(2, 20) <= input(58);
output(2, 21) <= input(33);
output(2, 22) <= input(34);
output(2, 23) <= input(35);
output(2, 24) <= input(36);
output(2, 25) <= input(37);
output(2, 26) <= input(38);
output(2, 27) <= input(39);
output(2, 28) <= input(40);
output(2, 29) <= input(41);
output(2, 30) <= input(42);
output(2, 31) <= input(43);
output(2, 32) <= input(31);
output(2, 33) <= input(32);
output(2, 34) <= input(0);
output(2, 35) <= input(1);
output(2, 36) <= input(2);
output(2, 37) <= input(3);
output(2, 38) <= input(4);
output(2, 39) <= input(5);
output(2, 40) <= input(6);
output(2, 41) <= input(7);
output(2, 42) <= input(8);
output(2, 43) <= input(9);
output(2, 44) <= input(10);
output(2, 45) <= input(11);
output(2, 46) <= input(12);
output(2, 47) <= input(13);
output(2, 48) <= input(32);
output(2, 49) <= input(0);
output(2, 50) <= input(1);
output(2, 51) <= input(2);
output(2, 52) <= input(3);
output(2, 53) <= input(4);
output(2, 54) <= input(5);
output(2, 55) <= input(6);
output(2, 56) <= input(7);
output(2, 57) <= input(8);
output(2, 58) <= input(9);
output(2, 59) <= input(10);
output(2, 60) <= input(11);
output(2, 61) <= input(12);
output(2, 62) <= input(13);
output(2, 63) <= input(14);
output(2, 64) <= input(0);
output(2, 65) <= input(1);
output(2, 66) <= input(2);
output(2, 67) <= input(3);
output(2, 68) <= input(4);
output(2, 69) <= input(5);
output(2, 70) <= input(6);
output(2, 71) <= input(7);
output(2, 72) <= input(8);
output(2, 73) <= input(9);
output(2, 74) <= input(10);
output(2, 75) <= input(11);
output(2, 76) <= input(12);
output(2, 77) <= input(13);
output(2, 78) <= input(14);
output(2, 79) <= input(15);
output(2, 80) <= input(57);
output(2, 81) <= input(58);
output(2, 82) <= input(33);
output(2, 83) <= input(34);
output(2, 84) <= input(35);
output(2, 85) <= input(36);
output(2, 86) <= input(37);
output(2, 87) <= input(38);
output(2, 88) <= input(39);
output(2, 89) <= input(40);
output(2, 90) <= input(41);
output(2, 91) <= input(42);
output(2, 92) <= input(43);
output(2, 93) <= input(44);
output(2, 94) <= input(45);
output(2, 95) <= input(46);
output(2, 96) <= input(58);
output(2, 97) <= input(33);
output(2, 98) <= input(34);
output(2, 99) <= input(35);
output(2, 100) <= input(36);
output(2, 101) <= input(37);
output(2, 102) <= input(38);
output(2, 103) <= input(39);
output(2, 104) <= input(40);
output(2, 105) <= input(41);
output(2, 106) <= input(42);
output(2, 107) <= input(43);
output(2, 108) <= input(44);
output(2, 109) <= input(45);
output(2, 110) <= input(46);
output(2, 111) <= input(47);
output(2, 112) <= input(33);
output(2, 113) <= input(34);
output(2, 114) <= input(35);
output(2, 115) <= input(36);
output(2, 116) <= input(37);
output(2, 117) <= input(38);
output(2, 118) <= input(39);
output(2, 119) <= input(40);
output(2, 120) <= input(41);
output(2, 121) <= input(42);
output(2, 122) <= input(43);
output(2, 123) <= input(44);
output(2, 124) <= input(45);
output(2, 125) <= input(46);
output(2, 126) <= input(47);
output(2, 127) <= input(48);
output(2, 128) <= input(3);
output(2, 129) <= input(4);
output(2, 130) <= input(5);
output(2, 131) <= input(6);
output(2, 132) <= input(7);
output(2, 133) <= input(8);
output(2, 134) <= input(9);
output(2, 135) <= input(10);
output(2, 136) <= input(11);
output(2, 137) <= input(12);
output(2, 138) <= input(13);
output(2, 139) <= input(14);
output(2, 140) <= input(15);
output(2, 141) <= input(16);
output(2, 142) <= input(17);
output(2, 143) <= input(18);
output(2, 144) <= input(4);
output(2, 145) <= input(5);
output(2, 146) <= input(6);
output(2, 147) <= input(7);
output(2, 148) <= input(8);
output(2, 149) <= input(9);
output(2, 150) <= input(10);
output(2, 151) <= input(11);
output(2, 152) <= input(12);
output(2, 153) <= input(13);
output(2, 154) <= input(14);
output(2, 155) <= input(15);
output(2, 156) <= input(16);
output(2, 157) <= input(17);
output(2, 158) <= input(18);
output(2, 159) <= input(19);
output(2, 160) <= input(35);
output(2, 161) <= input(36);
output(2, 162) <= input(37);
output(2, 163) <= input(38);
output(2, 164) <= input(39);
output(2, 165) <= input(40);
output(2, 166) <= input(41);
output(2, 167) <= input(42);
output(2, 168) <= input(43);
output(2, 169) <= input(44);
output(2, 170) <= input(45);
output(2, 171) <= input(46);
output(2, 172) <= input(47);
output(2, 173) <= input(48);
output(2, 174) <= input(49);
output(2, 175) <= input(50);
output(2, 176) <= input(36);
output(2, 177) <= input(37);
output(2, 178) <= input(38);
output(2, 179) <= input(39);
output(2, 180) <= input(40);
output(2, 181) <= input(41);
output(2, 182) <= input(42);
output(2, 183) <= input(43);
output(2, 184) <= input(44);
output(2, 185) <= input(45);
output(2, 186) <= input(46);
output(2, 187) <= input(47);
output(2, 188) <= input(48);
output(2, 189) <= input(49);
output(2, 190) <= input(50);
output(2, 191) <= input(51);
output(2, 192) <= input(37);
output(2, 193) <= input(38);
output(2, 194) <= input(39);
output(2, 195) <= input(40);
output(2, 196) <= input(41);
output(2, 197) <= input(42);
output(2, 198) <= input(43);
output(2, 199) <= input(44);
output(2, 200) <= input(45);
output(2, 201) <= input(46);
output(2, 202) <= input(47);
output(2, 203) <= input(48);
output(2, 204) <= input(49);
output(2, 205) <= input(50);
output(2, 206) <= input(51);
output(2, 207) <= input(52);
output(2, 208) <= input(7);
output(2, 209) <= input(8);
output(2, 210) <= input(9);
output(2, 211) <= input(10);
output(2, 212) <= input(11);
output(2, 213) <= input(12);
output(2, 214) <= input(13);
output(2, 215) <= input(14);
output(2, 216) <= input(15);
output(2, 217) <= input(16);
output(2, 218) <= input(17);
output(2, 219) <= input(18);
output(2, 220) <= input(19);
output(2, 221) <= input(20);
output(2, 222) <= input(21);
output(2, 223) <= input(22);
output(2, 224) <= input(8);
output(2, 225) <= input(9);
output(2, 226) <= input(10);
output(2, 227) <= input(11);
output(2, 228) <= input(12);
output(2, 229) <= input(13);
output(2, 230) <= input(14);
output(2, 231) <= input(15);
output(2, 232) <= input(16);
output(2, 233) <= input(17);
output(2, 234) <= input(18);
output(2, 235) <= input(19);
output(2, 236) <= input(20);
output(2, 237) <= input(21);
output(2, 238) <= input(22);
output(2, 239) <= input(23);
output(2, 240) <= input(9);
output(2, 241) <= input(10);
output(2, 242) <= input(11);
output(2, 243) <= input(12);
output(2, 244) <= input(13);
output(2, 245) <= input(14);
output(2, 246) <= input(15);
output(2, 247) <= input(16);
output(2, 248) <= input(17);
output(2, 249) <= input(18);
output(2, 250) <= input(19);
output(2, 251) <= input(20);
output(2, 252) <= input(21);
output(2, 253) <= input(22);
output(2, 254) <= input(23);
output(2, 255) <= input(24);
output(3, 0) <= input(59);
output(3, 1) <= input(60);
output(3, 2) <= input(61);
output(3, 3) <= input(31);
output(3, 4) <= input(32);
output(3, 5) <= input(0);
output(3, 6) <= input(1);
output(3, 7) <= input(2);
output(3, 8) <= input(3);
output(3, 9) <= input(4);
output(3, 10) <= input(5);
output(3, 11) <= input(6);
output(3, 12) <= input(7);
output(3, 13) <= input(8);
output(3, 14) <= input(9);
output(3, 15) <= input(10);
output(3, 16) <= input(62);
output(3, 17) <= input(53);
output(3, 18) <= input(54);
output(3, 19) <= input(55);
output(3, 20) <= input(56);
output(3, 21) <= input(57);
output(3, 22) <= input(58);
output(3, 23) <= input(33);
output(3, 24) <= input(34);
output(3, 25) <= input(35);
output(3, 26) <= input(36);
output(3, 27) <= input(37);
output(3, 28) <= input(38);
output(3, 29) <= input(39);
output(3, 30) <= input(40);
output(3, 31) <= input(41);
output(3, 32) <= input(53);
output(3, 33) <= input(54);
output(3, 34) <= input(55);
output(3, 35) <= input(56);
output(3, 36) <= input(57);
output(3, 37) <= input(58);
output(3, 38) <= input(33);
output(3, 39) <= input(34);
output(3, 40) <= input(35);
output(3, 41) <= input(36);
output(3, 42) <= input(37);
output(3, 43) <= input(38);
output(3, 44) <= input(39);
output(3, 45) <= input(40);
output(3, 46) <= input(41);
output(3, 47) <= input(42);
output(3, 48) <= input(61);
output(3, 49) <= input(31);
output(3, 50) <= input(32);
output(3, 51) <= input(0);
output(3, 52) <= input(1);
output(3, 53) <= input(2);
output(3, 54) <= input(3);
output(3, 55) <= input(4);
output(3, 56) <= input(5);
output(3, 57) <= input(6);
output(3, 58) <= input(7);
output(3, 59) <= input(8);
output(3, 60) <= input(9);
output(3, 61) <= input(10);
output(3, 62) <= input(11);
output(3, 63) <= input(12);
output(3, 64) <= input(31);
output(3, 65) <= input(32);
output(3, 66) <= input(0);
output(3, 67) <= input(1);
output(3, 68) <= input(2);
output(3, 69) <= input(3);
output(3, 70) <= input(4);
output(3, 71) <= input(5);
output(3, 72) <= input(6);
output(3, 73) <= input(7);
output(3, 74) <= input(8);
output(3, 75) <= input(9);
output(3, 76) <= input(10);
output(3, 77) <= input(11);
output(3, 78) <= input(12);
output(3, 79) <= input(13);
output(3, 80) <= input(55);
output(3, 81) <= input(56);
output(3, 82) <= input(57);
output(3, 83) <= input(58);
output(3, 84) <= input(33);
output(3, 85) <= input(34);
output(3, 86) <= input(35);
output(3, 87) <= input(36);
output(3, 88) <= input(37);
output(3, 89) <= input(38);
output(3, 90) <= input(39);
output(3, 91) <= input(40);
output(3, 92) <= input(41);
output(3, 93) <= input(42);
output(3, 94) <= input(43);
output(3, 95) <= input(44);
output(3, 96) <= input(56);
output(3, 97) <= input(57);
output(3, 98) <= input(58);
output(3, 99) <= input(33);
output(3, 100) <= input(34);
output(3, 101) <= input(35);
output(3, 102) <= input(36);
output(3, 103) <= input(37);
output(3, 104) <= input(38);
output(3, 105) <= input(39);
output(3, 106) <= input(40);
output(3, 107) <= input(41);
output(3, 108) <= input(42);
output(3, 109) <= input(43);
output(3, 110) <= input(44);
output(3, 111) <= input(45);
output(3, 112) <= input(0);
output(3, 113) <= input(1);
output(3, 114) <= input(2);
output(3, 115) <= input(3);
output(3, 116) <= input(4);
output(3, 117) <= input(5);
output(3, 118) <= input(6);
output(3, 119) <= input(7);
output(3, 120) <= input(8);
output(3, 121) <= input(9);
output(3, 122) <= input(10);
output(3, 123) <= input(11);
output(3, 124) <= input(12);
output(3, 125) <= input(13);
output(3, 126) <= input(14);
output(3, 127) <= input(15);
output(3, 128) <= input(57);
output(3, 129) <= input(58);
output(3, 130) <= input(33);
output(3, 131) <= input(34);
output(3, 132) <= input(35);
output(3, 133) <= input(36);
output(3, 134) <= input(37);
output(3, 135) <= input(38);
output(3, 136) <= input(39);
output(3, 137) <= input(40);
output(3, 138) <= input(41);
output(3, 139) <= input(42);
output(3, 140) <= input(43);
output(3, 141) <= input(44);
output(3, 142) <= input(45);
output(3, 143) <= input(46);
output(3, 144) <= input(58);
output(3, 145) <= input(33);
output(3, 146) <= input(34);
output(3, 147) <= input(35);
output(3, 148) <= input(36);
output(3, 149) <= input(37);
output(3, 150) <= input(38);
output(3, 151) <= input(39);
output(3, 152) <= input(40);
output(3, 153) <= input(41);
output(3, 154) <= input(42);
output(3, 155) <= input(43);
output(3, 156) <= input(44);
output(3, 157) <= input(45);
output(3, 158) <= input(46);
output(3, 159) <= input(47);
output(3, 160) <= input(2);
output(3, 161) <= input(3);
output(3, 162) <= input(4);
output(3, 163) <= input(5);
output(3, 164) <= input(6);
output(3, 165) <= input(7);
output(3, 166) <= input(8);
output(3, 167) <= input(9);
output(3, 168) <= input(10);
output(3, 169) <= input(11);
output(3, 170) <= input(12);
output(3, 171) <= input(13);
output(3, 172) <= input(14);
output(3, 173) <= input(15);
output(3, 174) <= input(16);
output(3, 175) <= input(17);
output(3, 176) <= input(3);
output(3, 177) <= input(4);
output(3, 178) <= input(5);
output(3, 179) <= input(6);
output(3, 180) <= input(7);
output(3, 181) <= input(8);
output(3, 182) <= input(9);
output(3, 183) <= input(10);
output(3, 184) <= input(11);
output(3, 185) <= input(12);
output(3, 186) <= input(13);
output(3, 187) <= input(14);
output(3, 188) <= input(15);
output(3, 189) <= input(16);
output(3, 190) <= input(17);
output(3, 191) <= input(18);
output(3, 192) <= input(34);
output(3, 193) <= input(35);
output(3, 194) <= input(36);
output(3, 195) <= input(37);
output(3, 196) <= input(38);
output(3, 197) <= input(39);
output(3, 198) <= input(40);
output(3, 199) <= input(41);
output(3, 200) <= input(42);
output(3, 201) <= input(43);
output(3, 202) <= input(44);
output(3, 203) <= input(45);
output(3, 204) <= input(46);
output(3, 205) <= input(47);
output(3, 206) <= input(48);
output(3, 207) <= input(49);
output(3, 208) <= input(35);
output(3, 209) <= input(36);
output(3, 210) <= input(37);
output(3, 211) <= input(38);
output(3, 212) <= input(39);
output(3, 213) <= input(40);
output(3, 214) <= input(41);
output(3, 215) <= input(42);
output(3, 216) <= input(43);
output(3, 217) <= input(44);
output(3, 218) <= input(45);
output(3, 219) <= input(46);
output(3, 220) <= input(47);
output(3, 221) <= input(48);
output(3, 222) <= input(49);
output(3, 223) <= input(50);
output(3, 224) <= input(5);
output(3, 225) <= input(6);
output(3, 226) <= input(7);
output(3, 227) <= input(8);
output(3, 228) <= input(9);
output(3, 229) <= input(10);
output(3, 230) <= input(11);
output(3, 231) <= input(12);
output(3, 232) <= input(13);
output(3, 233) <= input(14);
output(3, 234) <= input(15);
output(3, 235) <= input(16);
output(3, 236) <= input(17);
output(3, 237) <= input(18);
output(3, 238) <= input(19);
output(3, 239) <= input(20);
output(3, 240) <= input(6);
output(3, 241) <= input(7);
output(3, 242) <= input(8);
output(3, 243) <= input(9);
output(3, 244) <= input(10);
output(3, 245) <= input(11);
output(3, 246) <= input(12);
output(3, 247) <= input(13);
output(3, 248) <= input(14);
output(3, 249) <= input(15);
output(3, 250) <= input(16);
output(3, 251) <= input(17);
output(3, 252) <= input(18);
output(3, 253) <= input(19);
output(3, 254) <= input(20);
output(3, 255) <= input(21);
output(4, 0) <= input(63);
output(4, 1) <= input(64);
output(4, 2) <= input(62);
output(4, 3) <= input(53);
output(4, 4) <= input(54);
output(4, 5) <= input(55);
output(4, 6) <= input(56);
output(4, 7) <= input(57);
output(4, 8) <= input(58);
output(4, 9) <= input(33);
output(4, 10) <= input(34);
output(4, 11) <= input(35);
output(4, 12) <= input(36);
output(4, 13) <= input(37);
output(4, 14) <= input(38);
output(4, 15) <= input(39);
output(4, 16) <= input(65);
output(4, 17) <= input(59);
output(4, 18) <= input(60);
output(4, 19) <= input(61);
output(4, 20) <= input(31);
output(4, 21) <= input(32);
output(4, 22) <= input(0);
output(4, 23) <= input(1);
output(4, 24) <= input(2);
output(4, 25) <= input(3);
output(4, 26) <= input(4);
output(4, 27) <= input(5);
output(4, 28) <= input(6);
output(4, 29) <= input(7);
output(4, 30) <= input(8);
output(4, 31) <= input(9);
output(4, 32) <= input(64);
output(4, 33) <= input(62);
output(4, 34) <= input(53);
output(4, 35) <= input(54);
output(4, 36) <= input(55);
output(4, 37) <= input(56);
output(4, 38) <= input(57);
output(4, 39) <= input(58);
output(4, 40) <= input(33);
output(4, 41) <= input(34);
output(4, 42) <= input(35);
output(4, 43) <= input(36);
output(4, 44) <= input(37);
output(4, 45) <= input(38);
output(4, 46) <= input(39);
output(4, 47) <= input(40);
output(4, 48) <= input(62);
output(4, 49) <= input(53);
output(4, 50) <= input(54);
output(4, 51) <= input(55);
output(4, 52) <= input(56);
output(4, 53) <= input(57);
output(4, 54) <= input(58);
output(4, 55) <= input(33);
output(4, 56) <= input(34);
output(4, 57) <= input(35);
output(4, 58) <= input(36);
output(4, 59) <= input(37);
output(4, 60) <= input(38);
output(4, 61) <= input(39);
output(4, 62) <= input(40);
output(4, 63) <= input(41);
output(4, 64) <= input(60);
output(4, 65) <= input(61);
output(4, 66) <= input(31);
output(4, 67) <= input(32);
output(4, 68) <= input(0);
output(4, 69) <= input(1);
output(4, 70) <= input(2);
output(4, 71) <= input(3);
output(4, 72) <= input(4);
output(4, 73) <= input(5);
output(4, 74) <= input(6);
output(4, 75) <= input(7);
output(4, 76) <= input(8);
output(4, 77) <= input(9);
output(4, 78) <= input(10);
output(4, 79) <= input(11);
output(4, 80) <= input(53);
output(4, 81) <= input(54);
output(4, 82) <= input(55);
output(4, 83) <= input(56);
output(4, 84) <= input(57);
output(4, 85) <= input(58);
output(4, 86) <= input(33);
output(4, 87) <= input(34);
output(4, 88) <= input(35);
output(4, 89) <= input(36);
output(4, 90) <= input(37);
output(4, 91) <= input(38);
output(4, 92) <= input(39);
output(4, 93) <= input(40);
output(4, 94) <= input(41);
output(4, 95) <= input(42);
output(4, 96) <= input(61);
output(4, 97) <= input(31);
output(4, 98) <= input(32);
output(4, 99) <= input(0);
output(4, 100) <= input(1);
output(4, 101) <= input(2);
output(4, 102) <= input(3);
output(4, 103) <= input(4);
output(4, 104) <= input(5);
output(4, 105) <= input(6);
output(4, 106) <= input(7);
output(4, 107) <= input(8);
output(4, 108) <= input(9);
output(4, 109) <= input(10);
output(4, 110) <= input(11);
output(4, 111) <= input(12);
output(4, 112) <= input(31);
output(4, 113) <= input(32);
output(4, 114) <= input(0);
output(4, 115) <= input(1);
output(4, 116) <= input(2);
output(4, 117) <= input(3);
output(4, 118) <= input(4);
output(4, 119) <= input(5);
output(4, 120) <= input(6);
output(4, 121) <= input(7);
output(4, 122) <= input(8);
output(4, 123) <= input(9);
output(4, 124) <= input(10);
output(4, 125) <= input(11);
output(4, 126) <= input(12);
output(4, 127) <= input(13);
output(4, 128) <= input(55);
output(4, 129) <= input(56);
output(4, 130) <= input(57);
output(4, 131) <= input(58);
output(4, 132) <= input(33);
output(4, 133) <= input(34);
output(4, 134) <= input(35);
output(4, 135) <= input(36);
output(4, 136) <= input(37);
output(4, 137) <= input(38);
output(4, 138) <= input(39);
output(4, 139) <= input(40);
output(4, 140) <= input(41);
output(4, 141) <= input(42);
output(4, 142) <= input(43);
output(4, 143) <= input(44);
output(4, 144) <= input(32);
output(4, 145) <= input(0);
output(4, 146) <= input(1);
output(4, 147) <= input(2);
output(4, 148) <= input(3);
output(4, 149) <= input(4);
output(4, 150) <= input(5);
output(4, 151) <= input(6);
output(4, 152) <= input(7);
output(4, 153) <= input(8);
output(4, 154) <= input(9);
output(4, 155) <= input(10);
output(4, 156) <= input(11);
output(4, 157) <= input(12);
output(4, 158) <= input(13);
output(4, 159) <= input(14);
output(4, 160) <= input(56);
output(4, 161) <= input(57);
output(4, 162) <= input(58);
output(4, 163) <= input(33);
output(4, 164) <= input(34);
output(4, 165) <= input(35);
output(4, 166) <= input(36);
output(4, 167) <= input(37);
output(4, 168) <= input(38);
output(4, 169) <= input(39);
output(4, 170) <= input(40);
output(4, 171) <= input(41);
output(4, 172) <= input(42);
output(4, 173) <= input(43);
output(4, 174) <= input(44);
output(4, 175) <= input(45);
output(4, 176) <= input(57);
output(4, 177) <= input(58);
output(4, 178) <= input(33);
output(4, 179) <= input(34);
output(4, 180) <= input(35);
output(4, 181) <= input(36);
output(4, 182) <= input(37);
output(4, 183) <= input(38);
output(4, 184) <= input(39);
output(4, 185) <= input(40);
output(4, 186) <= input(41);
output(4, 187) <= input(42);
output(4, 188) <= input(43);
output(4, 189) <= input(44);
output(4, 190) <= input(45);
output(4, 191) <= input(46);
output(4, 192) <= input(1);
output(4, 193) <= input(2);
output(4, 194) <= input(3);
output(4, 195) <= input(4);
output(4, 196) <= input(5);
output(4, 197) <= input(6);
output(4, 198) <= input(7);
output(4, 199) <= input(8);
output(4, 200) <= input(9);
output(4, 201) <= input(10);
output(4, 202) <= input(11);
output(4, 203) <= input(12);
output(4, 204) <= input(13);
output(4, 205) <= input(14);
output(4, 206) <= input(15);
output(4, 207) <= input(16);
output(4, 208) <= input(58);
output(4, 209) <= input(33);
output(4, 210) <= input(34);
output(4, 211) <= input(35);
output(4, 212) <= input(36);
output(4, 213) <= input(37);
output(4, 214) <= input(38);
output(4, 215) <= input(39);
output(4, 216) <= input(40);
output(4, 217) <= input(41);
output(4, 218) <= input(42);
output(4, 219) <= input(43);
output(4, 220) <= input(44);
output(4, 221) <= input(45);
output(4, 222) <= input(46);
output(4, 223) <= input(47);
output(4, 224) <= input(2);
output(4, 225) <= input(3);
output(4, 226) <= input(4);
output(4, 227) <= input(5);
output(4, 228) <= input(6);
output(4, 229) <= input(7);
output(4, 230) <= input(8);
output(4, 231) <= input(9);
output(4, 232) <= input(10);
output(4, 233) <= input(11);
output(4, 234) <= input(12);
output(4, 235) <= input(13);
output(4, 236) <= input(14);
output(4, 237) <= input(15);
output(4, 238) <= input(16);
output(4, 239) <= input(17);
output(4, 240) <= input(3);
output(4, 241) <= input(4);
output(4, 242) <= input(5);
output(4, 243) <= input(6);
output(4, 244) <= input(7);
output(4, 245) <= input(8);
output(4, 246) <= input(9);
output(4, 247) <= input(10);
output(4, 248) <= input(11);
output(4, 249) <= input(12);
output(4, 250) <= input(13);
output(4, 251) <= input(14);
output(4, 252) <= input(15);
output(4, 253) <= input(16);
output(4, 254) <= input(17);
output(4, 255) <= input(18);
output(5, 0) <= input(66);
output(5, 1) <= input(63);
output(5, 2) <= input(64);
output(5, 3) <= input(62);
output(5, 4) <= input(53);
output(5, 5) <= input(54);
output(5, 6) <= input(55);
output(5, 7) <= input(56);
output(5, 8) <= input(57);
output(5, 9) <= input(58);
output(5, 10) <= input(33);
output(5, 11) <= input(34);
output(5, 12) <= input(35);
output(5, 13) <= input(36);
output(5, 14) <= input(37);
output(5, 15) <= input(38);
output(5, 16) <= input(67);
output(5, 17) <= input(65);
output(5, 18) <= input(59);
output(5, 19) <= input(60);
output(5, 20) <= input(61);
output(5, 21) <= input(31);
output(5, 22) <= input(32);
output(5, 23) <= input(0);
output(5, 24) <= input(1);
output(5, 25) <= input(2);
output(5, 26) <= input(3);
output(5, 27) <= input(4);
output(5, 28) <= input(5);
output(5, 29) <= input(6);
output(5, 30) <= input(7);
output(5, 31) <= input(8);
output(5, 32) <= input(63);
output(5, 33) <= input(64);
output(5, 34) <= input(62);
output(5, 35) <= input(53);
output(5, 36) <= input(54);
output(5, 37) <= input(55);
output(5, 38) <= input(56);
output(5, 39) <= input(57);
output(5, 40) <= input(58);
output(5, 41) <= input(33);
output(5, 42) <= input(34);
output(5, 43) <= input(35);
output(5, 44) <= input(36);
output(5, 45) <= input(37);
output(5, 46) <= input(38);
output(5, 47) <= input(39);
output(5, 48) <= input(65);
output(5, 49) <= input(59);
output(5, 50) <= input(60);
output(5, 51) <= input(61);
output(5, 52) <= input(31);
output(5, 53) <= input(32);
output(5, 54) <= input(0);
output(5, 55) <= input(1);
output(5, 56) <= input(2);
output(5, 57) <= input(3);
output(5, 58) <= input(4);
output(5, 59) <= input(5);
output(5, 60) <= input(6);
output(5, 61) <= input(7);
output(5, 62) <= input(8);
output(5, 63) <= input(9);
output(5, 64) <= input(64);
output(5, 65) <= input(62);
output(5, 66) <= input(53);
output(5, 67) <= input(54);
output(5, 68) <= input(55);
output(5, 69) <= input(56);
output(5, 70) <= input(57);
output(5, 71) <= input(58);
output(5, 72) <= input(33);
output(5, 73) <= input(34);
output(5, 74) <= input(35);
output(5, 75) <= input(36);
output(5, 76) <= input(37);
output(5, 77) <= input(38);
output(5, 78) <= input(39);
output(5, 79) <= input(40);
output(5, 80) <= input(59);
output(5, 81) <= input(60);
output(5, 82) <= input(61);
output(5, 83) <= input(31);
output(5, 84) <= input(32);
output(5, 85) <= input(0);
output(5, 86) <= input(1);
output(5, 87) <= input(2);
output(5, 88) <= input(3);
output(5, 89) <= input(4);
output(5, 90) <= input(5);
output(5, 91) <= input(6);
output(5, 92) <= input(7);
output(5, 93) <= input(8);
output(5, 94) <= input(9);
output(5, 95) <= input(10);
output(5, 96) <= input(62);
output(5, 97) <= input(53);
output(5, 98) <= input(54);
output(5, 99) <= input(55);
output(5, 100) <= input(56);
output(5, 101) <= input(57);
output(5, 102) <= input(58);
output(5, 103) <= input(33);
output(5, 104) <= input(34);
output(5, 105) <= input(35);
output(5, 106) <= input(36);
output(5, 107) <= input(37);
output(5, 108) <= input(38);
output(5, 109) <= input(39);
output(5, 110) <= input(40);
output(5, 111) <= input(41);
output(5, 112) <= input(53);
output(5, 113) <= input(54);
output(5, 114) <= input(55);
output(5, 115) <= input(56);
output(5, 116) <= input(57);
output(5, 117) <= input(58);
output(5, 118) <= input(33);
output(5, 119) <= input(34);
output(5, 120) <= input(35);
output(5, 121) <= input(36);
output(5, 122) <= input(37);
output(5, 123) <= input(38);
output(5, 124) <= input(39);
output(5, 125) <= input(40);
output(5, 126) <= input(41);
output(5, 127) <= input(42);
output(5, 128) <= input(61);
output(5, 129) <= input(31);
output(5, 130) <= input(32);
output(5, 131) <= input(0);
output(5, 132) <= input(1);
output(5, 133) <= input(2);
output(5, 134) <= input(3);
output(5, 135) <= input(4);
output(5, 136) <= input(5);
output(5, 137) <= input(6);
output(5, 138) <= input(7);
output(5, 139) <= input(8);
output(5, 140) <= input(9);
output(5, 141) <= input(10);
output(5, 142) <= input(11);
output(5, 143) <= input(12);
output(5, 144) <= input(54);
output(5, 145) <= input(55);
output(5, 146) <= input(56);
output(5, 147) <= input(57);
output(5, 148) <= input(58);
output(5, 149) <= input(33);
output(5, 150) <= input(34);
output(5, 151) <= input(35);
output(5, 152) <= input(36);
output(5, 153) <= input(37);
output(5, 154) <= input(38);
output(5, 155) <= input(39);
output(5, 156) <= input(40);
output(5, 157) <= input(41);
output(5, 158) <= input(42);
output(5, 159) <= input(43);
output(5, 160) <= input(31);
output(5, 161) <= input(32);
output(5, 162) <= input(0);
output(5, 163) <= input(1);
output(5, 164) <= input(2);
output(5, 165) <= input(3);
output(5, 166) <= input(4);
output(5, 167) <= input(5);
output(5, 168) <= input(6);
output(5, 169) <= input(7);
output(5, 170) <= input(8);
output(5, 171) <= input(9);
output(5, 172) <= input(10);
output(5, 173) <= input(11);
output(5, 174) <= input(12);
output(5, 175) <= input(13);
output(5, 176) <= input(55);
output(5, 177) <= input(56);
output(5, 178) <= input(57);
output(5, 179) <= input(58);
output(5, 180) <= input(33);
output(5, 181) <= input(34);
output(5, 182) <= input(35);
output(5, 183) <= input(36);
output(5, 184) <= input(37);
output(5, 185) <= input(38);
output(5, 186) <= input(39);
output(5, 187) <= input(40);
output(5, 188) <= input(41);
output(5, 189) <= input(42);
output(5, 190) <= input(43);
output(5, 191) <= input(44);
output(5, 192) <= input(32);
output(5, 193) <= input(0);
output(5, 194) <= input(1);
output(5, 195) <= input(2);
output(5, 196) <= input(3);
output(5, 197) <= input(4);
output(5, 198) <= input(5);
output(5, 199) <= input(6);
output(5, 200) <= input(7);
output(5, 201) <= input(8);
output(5, 202) <= input(9);
output(5, 203) <= input(10);
output(5, 204) <= input(11);
output(5, 205) <= input(12);
output(5, 206) <= input(13);
output(5, 207) <= input(14);
output(5, 208) <= input(56);
output(5, 209) <= input(57);
output(5, 210) <= input(58);
output(5, 211) <= input(33);
output(5, 212) <= input(34);
output(5, 213) <= input(35);
output(5, 214) <= input(36);
output(5, 215) <= input(37);
output(5, 216) <= input(38);
output(5, 217) <= input(39);
output(5, 218) <= input(40);
output(5, 219) <= input(41);
output(5, 220) <= input(42);
output(5, 221) <= input(43);
output(5, 222) <= input(44);
output(5, 223) <= input(45);
output(5, 224) <= input(0);
output(5, 225) <= input(1);
output(5, 226) <= input(2);
output(5, 227) <= input(3);
output(5, 228) <= input(4);
output(5, 229) <= input(5);
output(5, 230) <= input(6);
output(5, 231) <= input(7);
output(5, 232) <= input(8);
output(5, 233) <= input(9);
output(5, 234) <= input(10);
output(5, 235) <= input(11);
output(5, 236) <= input(12);
output(5, 237) <= input(13);
output(5, 238) <= input(14);
output(5, 239) <= input(15);
output(5, 240) <= input(1);
output(5, 241) <= input(2);
output(5, 242) <= input(3);
output(5, 243) <= input(4);
output(5, 244) <= input(5);
output(5, 245) <= input(6);
output(5, 246) <= input(7);
output(5, 247) <= input(8);
output(5, 248) <= input(9);
output(5, 249) <= input(10);
output(5, 250) <= input(11);
output(5, 251) <= input(12);
output(5, 252) <= input(13);
output(5, 253) <= input(14);
output(5, 254) <= input(15);
output(5, 255) <= input(16);
when "0001" =>
output(0, 0) <= input(0);
output(0, 1) <= input(1);
output(0, 2) <= input(2);
output(0, 3) <= input(3);
output(0, 4) <= input(4);
output(0, 5) <= input(5);
output(0, 6) <= input(6);
output(0, 7) <= input(7);
output(0, 8) <= input(8);
output(0, 9) <= input(9);
output(0, 10) <= input(10);
output(0, 11) <= input(11);
output(0, 12) <= input(12);
output(0, 13) <= input(13);
output(0, 14) <= input(14);
output(0, 15) <= input(15);
output(0, 16) <= input(16);
output(0, 17) <= input(17);
output(0, 18) <= input(18);
output(0, 19) <= input(19);
output(0, 20) <= input(20);
output(0, 21) <= input(21);
output(0, 22) <= input(22);
output(0, 23) <= input(23);
output(0, 24) <= input(24);
output(0, 25) <= input(25);
output(0, 26) <= input(26);
output(0, 27) <= input(27);
output(0, 28) <= input(28);
output(0, 29) <= input(29);
output(0, 30) <= input(30);
output(0, 31) <= input(31);
output(0, 32) <= input(1);
output(0, 33) <= input(2);
output(0, 34) <= input(3);
output(0, 35) <= input(4);
output(0, 36) <= input(5);
output(0, 37) <= input(6);
output(0, 38) <= input(7);
output(0, 39) <= input(8);
output(0, 40) <= input(9);
output(0, 41) <= input(10);
output(0, 42) <= input(11);
output(0, 43) <= input(12);
output(0, 44) <= input(13);
output(0, 45) <= input(14);
output(0, 46) <= input(15);
output(0, 47) <= input(32);
output(0, 48) <= input(17);
output(0, 49) <= input(18);
output(0, 50) <= input(19);
output(0, 51) <= input(20);
output(0, 52) <= input(21);
output(0, 53) <= input(22);
output(0, 54) <= input(23);
output(0, 55) <= input(24);
output(0, 56) <= input(25);
output(0, 57) <= input(26);
output(0, 58) <= input(27);
output(0, 59) <= input(28);
output(0, 60) <= input(29);
output(0, 61) <= input(30);
output(0, 62) <= input(31);
output(0, 63) <= input(33);
output(0, 64) <= input(2);
output(0, 65) <= input(3);
output(0, 66) <= input(4);
output(0, 67) <= input(5);
output(0, 68) <= input(6);
output(0, 69) <= input(7);
output(0, 70) <= input(8);
output(0, 71) <= input(9);
output(0, 72) <= input(10);
output(0, 73) <= input(11);
output(0, 74) <= input(12);
output(0, 75) <= input(13);
output(0, 76) <= input(14);
output(0, 77) <= input(15);
output(0, 78) <= input(32);
output(0, 79) <= input(34);
output(0, 80) <= input(18);
output(0, 81) <= input(19);
output(0, 82) <= input(20);
output(0, 83) <= input(21);
output(0, 84) <= input(22);
output(0, 85) <= input(23);
output(0, 86) <= input(24);
output(0, 87) <= input(25);
output(0, 88) <= input(26);
output(0, 89) <= input(27);
output(0, 90) <= input(28);
output(0, 91) <= input(29);
output(0, 92) <= input(30);
output(0, 93) <= input(31);
output(0, 94) <= input(33);
output(0, 95) <= input(35);
output(0, 96) <= input(3);
output(0, 97) <= input(4);
output(0, 98) <= input(5);
output(0, 99) <= input(6);
output(0, 100) <= input(7);
output(0, 101) <= input(8);
output(0, 102) <= input(9);
output(0, 103) <= input(10);
output(0, 104) <= input(11);
output(0, 105) <= input(12);
output(0, 106) <= input(13);
output(0, 107) <= input(14);
output(0, 108) <= input(15);
output(0, 109) <= input(32);
output(0, 110) <= input(34);
output(0, 111) <= input(36);
output(0, 112) <= input(19);
output(0, 113) <= input(20);
output(0, 114) <= input(21);
output(0, 115) <= input(22);
output(0, 116) <= input(23);
output(0, 117) <= input(24);
output(0, 118) <= input(25);
output(0, 119) <= input(26);
output(0, 120) <= input(27);
output(0, 121) <= input(28);
output(0, 122) <= input(29);
output(0, 123) <= input(30);
output(0, 124) <= input(31);
output(0, 125) <= input(33);
output(0, 126) <= input(35);
output(0, 127) <= input(37);
output(0, 128) <= input(4);
output(0, 129) <= input(5);
output(0, 130) <= input(6);
output(0, 131) <= input(7);
output(0, 132) <= input(8);
output(0, 133) <= input(9);
output(0, 134) <= input(10);
output(0, 135) <= input(11);
output(0, 136) <= input(12);
output(0, 137) <= input(13);
output(0, 138) <= input(14);
output(0, 139) <= input(15);
output(0, 140) <= input(32);
output(0, 141) <= input(34);
output(0, 142) <= input(36);
output(0, 143) <= input(38);
output(0, 144) <= input(20);
output(0, 145) <= input(21);
output(0, 146) <= input(22);
output(0, 147) <= input(23);
output(0, 148) <= input(24);
output(0, 149) <= input(25);
output(0, 150) <= input(26);
output(0, 151) <= input(27);
output(0, 152) <= input(28);
output(0, 153) <= input(29);
output(0, 154) <= input(30);
output(0, 155) <= input(31);
output(0, 156) <= input(33);
output(0, 157) <= input(35);
output(0, 158) <= input(37);
output(0, 159) <= input(39);
output(0, 160) <= input(5);
output(0, 161) <= input(6);
output(0, 162) <= input(7);
output(0, 163) <= input(8);
output(0, 164) <= input(9);
output(0, 165) <= input(10);
output(0, 166) <= input(11);
output(0, 167) <= input(12);
output(0, 168) <= input(13);
output(0, 169) <= input(14);
output(0, 170) <= input(15);
output(0, 171) <= input(32);
output(0, 172) <= input(34);
output(0, 173) <= input(36);
output(0, 174) <= input(38);
output(0, 175) <= input(40);
output(0, 176) <= input(21);
output(0, 177) <= input(22);
output(0, 178) <= input(23);
output(0, 179) <= input(24);
output(0, 180) <= input(25);
output(0, 181) <= input(26);
output(0, 182) <= input(27);
output(0, 183) <= input(28);
output(0, 184) <= input(29);
output(0, 185) <= input(30);
output(0, 186) <= input(31);
output(0, 187) <= input(33);
output(0, 188) <= input(35);
output(0, 189) <= input(37);
output(0, 190) <= input(39);
output(0, 191) <= input(41);
output(0, 192) <= input(6);
output(0, 193) <= input(7);
output(0, 194) <= input(8);
output(0, 195) <= input(9);
output(0, 196) <= input(10);
output(0, 197) <= input(11);
output(0, 198) <= input(12);
output(0, 199) <= input(13);
output(0, 200) <= input(14);
output(0, 201) <= input(15);
output(0, 202) <= input(32);
output(0, 203) <= input(34);
output(0, 204) <= input(36);
output(0, 205) <= input(38);
output(0, 206) <= input(40);
output(0, 207) <= input(42);
output(0, 208) <= input(22);
output(0, 209) <= input(23);
output(0, 210) <= input(24);
output(0, 211) <= input(25);
output(0, 212) <= input(26);
output(0, 213) <= input(27);
output(0, 214) <= input(28);
output(0, 215) <= input(29);
output(0, 216) <= input(30);
output(0, 217) <= input(31);
output(0, 218) <= input(33);
output(0, 219) <= input(35);
output(0, 220) <= input(37);
output(0, 221) <= input(39);
output(0, 222) <= input(41);
output(0, 223) <= input(43);
output(0, 224) <= input(7);
output(0, 225) <= input(8);
output(0, 226) <= input(9);
output(0, 227) <= input(10);
output(0, 228) <= input(11);
output(0, 229) <= input(12);
output(0, 230) <= input(13);
output(0, 231) <= input(14);
output(0, 232) <= input(15);
output(0, 233) <= input(32);
output(0, 234) <= input(34);
output(0, 235) <= input(36);
output(0, 236) <= input(38);
output(0, 237) <= input(40);
output(0, 238) <= input(42);
output(0, 239) <= input(44);
output(0, 240) <= input(23);
output(0, 241) <= input(24);
output(0, 242) <= input(25);
output(0, 243) <= input(26);
output(0, 244) <= input(27);
output(0, 245) <= input(28);
output(0, 246) <= input(29);
output(0, 247) <= input(30);
output(0, 248) <= input(31);
output(0, 249) <= input(33);
output(0, 250) <= input(35);
output(0, 251) <= input(37);
output(0, 252) <= input(39);
output(0, 253) <= input(41);
output(0, 254) <= input(43);
output(0, 255) <= input(45);
output(1, 0) <= input(46);
output(1, 1) <= input(47);
output(1, 2) <= input(16);
output(1, 3) <= input(17);
output(1, 4) <= input(18);
output(1, 5) <= input(19);
output(1, 6) <= input(20);
output(1, 7) <= input(21);
output(1, 8) <= input(22);
output(1, 9) <= input(23);
output(1, 10) <= input(24);
output(1, 11) <= input(25);
output(1, 12) <= input(26);
output(1, 13) <= input(27);
output(1, 14) <= input(28);
output(1, 15) <= input(29);
output(1, 16) <= input(48);
output(1, 17) <= input(0);
output(1, 18) <= input(1);
output(1, 19) <= input(2);
output(1, 20) <= input(3);
output(1, 21) <= input(4);
output(1, 22) <= input(5);
output(1, 23) <= input(6);
output(1, 24) <= input(7);
output(1, 25) <= input(8);
output(1, 26) <= input(9);
output(1, 27) <= input(10);
output(1, 28) <= input(11);
output(1, 29) <= input(12);
output(1, 30) <= input(13);
output(1, 31) <= input(14);
output(1, 32) <= input(47);
output(1, 33) <= input(16);
output(1, 34) <= input(17);
output(1, 35) <= input(18);
output(1, 36) <= input(19);
output(1, 37) <= input(20);
output(1, 38) <= input(21);
output(1, 39) <= input(22);
output(1, 40) <= input(23);
output(1, 41) <= input(24);
output(1, 42) <= input(25);
output(1, 43) <= input(26);
output(1, 44) <= input(27);
output(1, 45) <= input(28);
output(1, 46) <= input(29);
output(1, 47) <= input(30);
output(1, 48) <= input(0);
output(1, 49) <= input(1);
output(1, 50) <= input(2);
output(1, 51) <= input(3);
output(1, 52) <= input(4);
output(1, 53) <= input(5);
output(1, 54) <= input(6);
output(1, 55) <= input(7);
output(1, 56) <= input(8);
output(1, 57) <= input(9);
output(1, 58) <= input(10);
output(1, 59) <= input(11);
output(1, 60) <= input(12);
output(1, 61) <= input(13);
output(1, 62) <= input(14);
output(1, 63) <= input(15);
output(1, 64) <= input(16);
output(1, 65) <= input(17);
output(1, 66) <= input(18);
output(1, 67) <= input(19);
output(1, 68) <= input(20);
output(1, 69) <= input(21);
output(1, 70) <= input(22);
output(1, 71) <= input(23);
output(1, 72) <= input(24);
output(1, 73) <= input(25);
output(1, 74) <= input(26);
output(1, 75) <= input(27);
output(1, 76) <= input(28);
output(1, 77) <= input(29);
output(1, 78) <= input(30);
output(1, 79) <= input(31);
output(1, 80) <= input(1);
output(1, 81) <= input(2);
output(1, 82) <= input(3);
output(1, 83) <= input(4);
output(1, 84) <= input(5);
output(1, 85) <= input(6);
output(1, 86) <= input(7);
output(1, 87) <= input(8);
output(1, 88) <= input(9);
output(1, 89) <= input(10);
output(1, 90) <= input(11);
output(1, 91) <= input(12);
output(1, 92) <= input(13);
output(1, 93) <= input(14);
output(1, 94) <= input(15);
output(1, 95) <= input(32);
output(1, 96) <= input(17);
output(1, 97) <= input(18);
output(1, 98) <= input(19);
output(1, 99) <= input(20);
output(1, 100) <= input(21);
output(1, 101) <= input(22);
output(1, 102) <= input(23);
output(1, 103) <= input(24);
output(1, 104) <= input(25);
output(1, 105) <= input(26);
output(1, 106) <= input(27);
output(1, 107) <= input(28);
output(1, 108) <= input(29);
output(1, 109) <= input(30);
output(1, 110) <= input(31);
output(1, 111) <= input(33);
output(1, 112) <= input(2);
output(1, 113) <= input(3);
output(1, 114) <= input(4);
output(1, 115) <= input(5);
output(1, 116) <= input(6);
output(1, 117) <= input(7);
output(1, 118) <= input(8);
output(1, 119) <= input(9);
output(1, 120) <= input(10);
output(1, 121) <= input(11);
output(1, 122) <= input(12);
output(1, 123) <= input(13);
output(1, 124) <= input(14);
output(1, 125) <= input(15);
output(1, 126) <= input(32);
output(1, 127) <= input(34);
output(1, 128) <= input(2);
output(1, 129) <= input(3);
output(1, 130) <= input(4);
output(1, 131) <= input(5);
output(1, 132) <= input(6);
output(1, 133) <= input(7);
output(1, 134) <= input(8);
output(1, 135) <= input(9);
output(1, 136) <= input(10);
output(1, 137) <= input(11);
output(1, 138) <= input(12);
output(1, 139) <= input(13);
output(1, 140) <= input(14);
output(1, 141) <= input(15);
output(1, 142) <= input(32);
output(1, 143) <= input(34);
output(1, 144) <= input(18);
output(1, 145) <= input(19);
output(1, 146) <= input(20);
output(1, 147) <= input(21);
output(1, 148) <= input(22);
output(1, 149) <= input(23);
output(1, 150) <= input(24);
output(1, 151) <= input(25);
output(1, 152) <= input(26);
output(1, 153) <= input(27);
output(1, 154) <= input(28);
output(1, 155) <= input(29);
output(1, 156) <= input(30);
output(1, 157) <= input(31);
output(1, 158) <= input(33);
output(1, 159) <= input(35);
output(1, 160) <= input(3);
output(1, 161) <= input(4);
output(1, 162) <= input(5);
output(1, 163) <= input(6);
output(1, 164) <= input(7);
output(1, 165) <= input(8);
output(1, 166) <= input(9);
output(1, 167) <= input(10);
output(1, 168) <= input(11);
output(1, 169) <= input(12);
output(1, 170) <= input(13);
output(1, 171) <= input(14);
output(1, 172) <= input(15);
output(1, 173) <= input(32);
output(1, 174) <= input(34);
output(1, 175) <= input(36);
output(1, 176) <= input(19);
output(1, 177) <= input(20);
output(1, 178) <= input(21);
output(1, 179) <= input(22);
output(1, 180) <= input(23);
output(1, 181) <= input(24);
output(1, 182) <= input(25);
output(1, 183) <= input(26);
output(1, 184) <= input(27);
output(1, 185) <= input(28);
output(1, 186) <= input(29);
output(1, 187) <= input(30);
output(1, 188) <= input(31);
output(1, 189) <= input(33);
output(1, 190) <= input(35);
output(1, 191) <= input(37);
output(1, 192) <= input(4);
output(1, 193) <= input(5);
output(1, 194) <= input(6);
output(1, 195) <= input(7);
output(1, 196) <= input(8);
output(1, 197) <= input(9);
output(1, 198) <= input(10);
output(1, 199) <= input(11);
output(1, 200) <= input(12);
output(1, 201) <= input(13);
output(1, 202) <= input(14);
output(1, 203) <= input(15);
output(1, 204) <= input(32);
output(1, 205) <= input(34);
output(1, 206) <= input(36);
output(1, 207) <= input(38);
output(1, 208) <= input(20);
output(1, 209) <= input(21);
output(1, 210) <= input(22);
output(1, 211) <= input(23);
output(1, 212) <= input(24);
output(1, 213) <= input(25);
output(1, 214) <= input(26);
output(1, 215) <= input(27);
output(1, 216) <= input(28);
output(1, 217) <= input(29);
output(1, 218) <= input(30);
output(1, 219) <= input(31);
output(1, 220) <= input(33);
output(1, 221) <= input(35);
output(1, 222) <= input(37);
output(1, 223) <= input(39);
output(1, 224) <= input(5);
output(1, 225) <= input(6);
output(1, 226) <= input(7);
output(1, 227) <= input(8);
output(1, 228) <= input(9);
output(1, 229) <= input(10);
output(1, 230) <= input(11);
output(1, 231) <= input(12);
output(1, 232) <= input(13);
output(1, 233) <= input(14);
output(1, 234) <= input(15);
output(1, 235) <= input(32);
output(1, 236) <= input(34);
output(1, 237) <= input(36);
output(1, 238) <= input(38);
output(1, 239) <= input(40);
output(1, 240) <= input(21);
output(1, 241) <= input(22);
output(1, 242) <= input(23);
output(1, 243) <= input(24);
output(1, 244) <= input(25);
output(1, 245) <= input(26);
output(1, 246) <= input(27);
output(1, 247) <= input(28);
output(1, 248) <= input(29);
output(1, 249) <= input(30);
output(1, 250) <= input(31);
output(1, 251) <= input(33);
output(1, 252) <= input(35);
output(1, 253) <= input(37);
output(1, 254) <= input(39);
output(1, 255) <= input(41);
output(2, 0) <= input(49);
output(2, 1) <= input(46);
output(2, 2) <= input(47);
output(2, 3) <= input(16);
output(2, 4) <= input(17);
output(2, 5) <= input(18);
output(2, 6) <= input(19);
output(2, 7) <= input(20);
output(2, 8) <= input(21);
output(2, 9) <= input(22);
output(2, 10) <= input(23);
output(2, 11) <= input(24);
output(2, 12) <= input(25);
output(2, 13) <= input(26);
output(2, 14) <= input(27);
output(2, 15) <= input(28);
output(2, 16) <= input(50);
output(2, 17) <= input(48);
output(2, 18) <= input(0);
output(2, 19) <= input(1);
output(2, 20) <= input(2);
output(2, 21) <= input(3);
output(2, 22) <= input(4);
output(2, 23) <= input(5);
output(2, 24) <= input(6);
output(2, 25) <= input(7);
output(2, 26) <= input(8);
output(2, 27) <= input(9);
output(2, 28) <= input(10);
output(2, 29) <= input(11);
output(2, 30) <= input(12);
output(2, 31) <= input(13);
output(2, 32) <= input(46);
output(2, 33) <= input(47);
output(2, 34) <= input(16);
output(2, 35) <= input(17);
output(2, 36) <= input(18);
output(2, 37) <= input(19);
output(2, 38) <= input(20);
output(2, 39) <= input(21);
output(2, 40) <= input(22);
output(2, 41) <= input(23);
output(2, 42) <= input(24);
output(2, 43) <= input(25);
output(2, 44) <= input(26);
output(2, 45) <= input(27);
output(2, 46) <= input(28);
output(2, 47) <= input(29);
output(2, 48) <= input(48);
output(2, 49) <= input(0);
output(2, 50) <= input(1);
output(2, 51) <= input(2);
output(2, 52) <= input(3);
output(2, 53) <= input(4);
output(2, 54) <= input(5);
output(2, 55) <= input(6);
output(2, 56) <= input(7);
output(2, 57) <= input(8);
output(2, 58) <= input(9);
output(2, 59) <= input(10);
output(2, 60) <= input(11);
output(2, 61) <= input(12);
output(2, 62) <= input(13);
output(2, 63) <= input(14);
output(2, 64) <= input(48);
output(2, 65) <= input(0);
output(2, 66) <= input(1);
output(2, 67) <= input(2);
output(2, 68) <= input(3);
output(2, 69) <= input(4);
output(2, 70) <= input(5);
output(2, 71) <= input(6);
output(2, 72) <= input(7);
output(2, 73) <= input(8);
output(2, 74) <= input(9);
output(2, 75) <= input(10);
output(2, 76) <= input(11);
output(2, 77) <= input(12);
output(2, 78) <= input(13);
output(2, 79) <= input(14);
output(2, 80) <= input(47);
output(2, 81) <= input(16);
output(2, 82) <= input(17);
output(2, 83) <= input(18);
output(2, 84) <= input(19);
output(2, 85) <= input(20);
output(2, 86) <= input(21);
output(2, 87) <= input(22);
output(2, 88) <= input(23);
output(2, 89) <= input(24);
output(2, 90) <= input(25);
output(2, 91) <= input(26);
output(2, 92) <= input(27);
output(2, 93) <= input(28);
output(2, 94) <= input(29);
output(2, 95) <= input(30);
output(2, 96) <= input(0);
output(2, 97) <= input(1);
output(2, 98) <= input(2);
output(2, 99) <= input(3);
output(2, 100) <= input(4);
output(2, 101) <= input(5);
output(2, 102) <= input(6);
output(2, 103) <= input(7);
output(2, 104) <= input(8);
output(2, 105) <= input(9);
output(2, 106) <= input(10);
output(2, 107) <= input(11);
output(2, 108) <= input(12);
output(2, 109) <= input(13);
output(2, 110) <= input(14);
output(2, 111) <= input(15);
output(2, 112) <= input(16);
output(2, 113) <= input(17);
output(2, 114) <= input(18);
output(2, 115) <= input(19);
output(2, 116) <= input(20);
output(2, 117) <= input(21);
output(2, 118) <= input(22);
output(2, 119) <= input(23);
output(2, 120) <= input(24);
output(2, 121) <= input(25);
output(2, 122) <= input(26);
output(2, 123) <= input(27);
output(2, 124) <= input(28);
output(2, 125) <= input(29);
output(2, 126) <= input(30);
output(2, 127) <= input(31);
output(2, 128) <= input(16);
output(2, 129) <= input(17);
output(2, 130) <= input(18);
output(2, 131) <= input(19);
output(2, 132) <= input(20);
output(2, 133) <= input(21);
output(2, 134) <= input(22);
output(2, 135) <= input(23);
output(2, 136) <= input(24);
output(2, 137) <= input(25);
output(2, 138) <= input(26);
output(2, 139) <= input(27);
output(2, 140) <= input(28);
output(2, 141) <= input(29);
output(2, 142) <= input(30);
output(2, 143) <= input(31);
output(2, 144) <= input(1);
output(2, 145) <= input(2);
output(2, 146) <= input(3);
output(2, 147) <= input(4);
output(2, 148) <= input(5);
output(2, 149) <= input(6);
output(2, 150) <= input(7);
output(2, 151) <= input(8);
output(2, 152) <= input(9);
output(2, 153) <= input(10);
output(2, 154) <= input(11);
output(2, 155) <= input(12);
output(2, 156) <= input(13);
output(2, 157) <= input(14);
output(2, 158) <= input(15);
output(2, 159) <= input(32);
output(2, 160) <= input(17);
output(2, 161) <= input(18);
output(2, 162) <= input(19);
output(2, 163) <= input(20);
output(2, 164) <= input(21);
output(2, 165) <= input(22);
output(2, 166) <= input(23);
output(2, 167) <= input(24);
output(2, 168) <= input(25);
output(2, 169) <= input(26);
output(2, 170) <= input(27);
output(2, 171) <= input(28);
output(2, 172) <= input(29);
output(2, 173) <= input(30);
output(2, 174) <= input(31);
output(2, 175) <= input(33);
output(2, 176) <= input(2);
output(2, 177) <= input(3);
output(2, 178) <= input(4);
output(2, 179) <= input(5);
output(2, 180) <= input(6);
output(2, 181) <= input(7);
output(2, 182) <= input(8);
output(2, 183) <= input(9);
output(2, 184) <= input(10);
output(2, 185) <= input(11);
output(2, 186) <= input(12);
output(2, 187) <= input(13);
output(2, 188) <= input(14);
output(2, 189) <= input(15);
output(2, 190) <= input(32);
output(2, 191) <= input(34);
output(2, 192) <= input(2);
output(2, 193) <= input(3);
output(2, 194) <= input(4);
output(2, 195) <= input(5);
output(2, 196) <= input(6);
output(2, 197) <= input(7);
output(2, 198) <= input(8);
output(2, 199) <= input(9);
output(2, 200) <= input(10);
output(2, 201) <= input(11);
output(2, 202) <= input(12);
output(2, 203) <= input(13);
output(2, 204) <= input(14);
output(2, 205) <= input(15);
output(2, 206) <= input(32);
output(2, 207) <= input(34);
output(2, 208) <= input(18);
output(2, 209) <= input(19);
output(2, 210) <= input(20);
output(2, 211) <= input(21);
output(2, 212) <= input(22);
output(2, 213) <= input(23);
output(2, 214) <= input(24);
output(2, 215) <= input(25);
output(2, 216) <= input(26);
output(2, 217) <= input(27);
output(2, 218) <= input(28);
output(2, 219) <= input(29);
output(2, 220) <= input(30);
output(2, 221) <= input(31);
output(2, 222) <= input(33);
output(2, 223) <= input(35);
output(2, 224) <= input(3);
output(2, 225) <= input(4);
output(2, 226) <= input(5);
output(2, 227) <= input(6);
output(2, 228) <= input(7);
output(2, 229) <= input(8);
output(2, 230) <= input(9);
output(2, 231) <= input(10);
output(2, 232) <= input(11);
output(2, 233) <= input(12);
output(2, 234) <= input(13);
output(2, 235) <= input(14);
output(2, 236) <= input(15);
output(2, 237) <= input(32);
output(2, 238) <= input(34);
output(2, 239) <= input(36);
output(2, 240) <= input(19);
output(2, 241) <= input(20);
output(2, 242) <= input(21);
output(2, 243) <= input(22);
output(2, 244) <= input(23);
output(2, 245) <= input(24);
output(2, 246) <= input(25);
output(2, 247) <= input(26);
output(2, 248) <= input(27);
output(2, 249) <= input(28);
output(2, 250) <= input(29);
output(2, 251) <= input(30);
output(2, 252) <= input(31);
output(2, 253) <= input(33);
output(2, 254) <= input(35);
output(2, 255) <= input(37);
output(3, 0) <= input(51);
output(3, 1) <= input(49);
output(3, 2) <= input(46);
output(3, 3) <= input(47);
output(3, 4) <= input(16);
output(3, 5) <= input(17);
output(3, 6) <= input(18);
output(3, 7) <= input(19);
output(3, 8) <= input(20);
output(3, 9) <= input(21);
output(3, 10) <= input(22);
output(3, 11) <= input(23);
output(3, 12) <= input(24);
output(3, 13) <= input(25);
output(3, 14) <= input(26);
output(3, 15) <= input(27);
output(3, 16) <= input(52);
output(3, 17) <= input(50);
output(3, 18) <= input(48);
output(3, 19) <= input(0);
output(3, 20) <= input(1);
output(3, 21) <= input(2);
output(3, 22) <= input(3);
output(3, 23) <= input(4);
output(3, 24) <= input(5);
output(3, 25) <= input(6);
output(3, 26) <= input(7);
output(3, 27) <= input(8);
output(3, 28) <= input(9);
output(3, 29) <= input(10);
output(3, 30) <= input(11);
output(3, 31) <= input(12);
output(3, 32) <= input(52);
output(3, 33) <= input(50);
output(3, 34) <= input(48);
output(3, 35) <= input(0);
output(3, 36) <= input(1);
output(3, 37) <= input(2);
output(3, 38) <= input(3);
output(3, 39) <= input(4);
output(3, 40) <= input(5);
output(3, 41) <= input(6);
output(3, 42) <= input(7);
output(3, 43) <= input(8);
output(3, 44) <= input(9);
output(3, 45) <= input(10);
output(3, 46) <= input(11);
output(3, 47) <= input(12);
output(3, 48) <= input(49);
output(3, 49) <= input(46);
output(3, 50) <= input(47);
output(3, 51) <= input(16);
output(3, 52) <= input(17);
output(3, 53) <= input(18);
output(3, 54) <= input(19);
output(3, 55) <= input(20);
output(3, 56) <= input(21);
output(3, 57) <= input(22);
output(3, 58) <= input(23);
output(3, 59) <= input(24);
output(3, 60) <= input(25);
output(3, 61) <= input(26);
output(3, 62) <= input(27);
output(3, 63) <= input(28);
output(3, 64) <= input(50);
output(3, 65) <= input(48);
output(3, 66) <= input(0);
output(3, 67) <= input(1);
output(3, 68) <= input(2);
output(3, 69) <= input(3);
output(3, 70) <= input(4);
output(3, 71) <= input(5);
output(3, 72) <= input(6);
output(3, 73) <= input(7);
output(3, 74) <= input(8);
output(3, 75) <= input(9);
output(3, 76) <= input(10);
output(3, 77) <= input(11);
output(3, 78) <= input(12);
output(3, 79) <= input(13);
output(3, 80) <= input(50);
output(3, 81) <= input(48);
output(3, 82) <= input(0);
output(3, 83) <= input(1);
output(3, 84) <= input(2);
output(3, 85) <= input(3);
output(3, 86) <= input(4);
output(3, 87) <= input(5);
output(3, 88) <= input(6);
output(3, 89) <= input(7);
output(3, 90) <= input(8);
output(3, 91) <= input(9);
output(3, 92) <= input(10);
output(3, 93) <= input(11);
output(3, 94) <= input(12);
output(3, 95) <= input(13);
output(3, 96) <= input(46);
output(3, 97) <= input(47);
output(3, 98) <= input(16);
output(3, 99) <= input(17);
output(3, 100) <= input(18);
output(3, 101) <= input(19);
output(3, 102) <= input(20);
output(3, 103) <= input(21);
output(3, 104) <= input(22);
output(3, 105) <= input(23);
output(3, 106) <= input(24);
output(3, 107) <= input(25);
output(3, 108) <= input(26);
output(3, 109) <= input(27);
output(3, 110) <= input(28);
output(3, 111) <= input(29);
output(3, 112) <= input(48);
output(3, 113) <= input(0);
output(3, 114) <= input(1);
output(3, 115) <= input(2);
output(3, 116) <= input(3);
output(3, 117) <= input(4);
output(3, 118) <= input(5);
output(3, 119) <= input(6);
output(3, 120) <= input(7);
output(3, 121) <= input(8);
output(3, 122) <= input(9);
output(3, 123) <= input(10);
output(3, 124) <= input(11);
output(3, 125) <= input(12);
output(3, 126) <= input(13);
output(3, 127) <= input(14);
output(3, 128) <= input(48);
output(3, 129) <= input(0);
output(3, 130) <= input(1);
output(3, 131) <= input(2);
output(3, 132) <= input(3);
output(3, 133) <= input(4);
output(3, 134) <= input(5);
output(3, 135) <= input(6);
output(3, 136) <= input(7);
output(3, 137) <= input(8);
output(3, 138) <= input(9);
output(3, 139) <= input(10);
output(3, 140) <= input(11);
output(3, 141) <= input(12);
output(3, 142) <= input(13);
output(3, 143) <= input(14);
output(3, 144) <= input(47);
output(3, 145) <= input(16);
output(3, 146) <= input(17);
output(3, 147) <= input(18);
output(3, 148) <= input(19);
output(3, 149) <= input(20);
output(3, 150) <= input(21);
output(3, 151) <= input(22);
output(3, 152) <= input(23);
output(3, 153) <= input(24);
output(3, 154) <= input(25);
output(3, 155) <= input(26);
output(3, 156) <= input(27);
output(3, 157) <= input(28);
output(3, 158) <= input(29);
output(3, 159) <= input(30);
output(3, 160) <= input(47);
output(3, 161) <= input(16);
output(3, 162) <= input(17);
output(3, 163) <= input(18);
output(3, 164) <= input(19);
output(3, 165) <= input(20);
output(3, 166) <= input(21);
output(3, 167) <= input(22);
output(3, 168) <= input(23);
output(3, 169) <= input(24);
output(3, 170) <= input(25);
output(3, 171) <= input(26);
output(3, 172) <= input(27);
output(3, 173) <= input(28);
output(3, 174) <= input(29);
output(3, 175) <= input(30);
output(3, 176) <= input(0);
output(3, 177) <= input(1);
output(3, 178) <= input(2);
output(3, 179) <= input(3);
output(3, 180) <= input(4);
output(3, 181) <= input(5);
output(3, 182) <= input(6);
output(3, 183) <= input(7);
output(3, 184) <= input(8);
output(3, 185) <= input(9);
output(3, 186) <= input(10);
output(3, 187) <= input(11);
output(3, 188) <= input(12);
output(3, 189) <= input(13);
output(3, 190) <= input(14);
output(3, 191) <= input(15);
output(3, 192) <= input(16);
output(3, 193) <= input(17);
output(3, 194) <= input(18);
output(3, 195) <= input(19);
output(3, 196) <= input(20);
output(3, 197) <= input(21);
output(3, 198) <= input(22);
output(3, 199) <= input(23);
output(3, 200) <= input(24);
output(3, 201) <= input(25);
output(3, 202) <= input(26);
output(3, 203) <= input(27);
output(3, 204) <= input(28);
output(3, 205) <= input(29);
output(3, 206) <= input(30);
output(3, 207) <= input(31);
output(3, 208) <= input(16);
output(3, 209) <= input(17);
output(3, 210) <= input(18);
output(3, 211) <= input(19);
output(3, 212) <= input(20);
output(3, 213) <= input(21);
output(3, 214) <= input(22);
output(3, 215) <= input(23);
output(3, 216) <= input(24);
output(3, 217) <= input(25);
output(3, 218) <= input(26);
output(3, 219) <= input(27);
output(3, 220) <= input(28);
output(3, 221) <= input(29);
output(3, 222) <= input(30);
output(3, 223) <= input(31);
output(3, 224) <= input(1);
output(3, 225) <= input(2);
output(3, 226) <= input(3);
output(3, 227) <= input(4);
output(3, 228) <= input(5);
output(3, 229) <= input(6);
output(3, 230) <= input(7);
output(3, 231) <= input(8);
output(3, 232) <= input(9);
output(3, 233) <= input(10);
output(3, 234) <= input(11);
output(3, 235) <= input(12);
output(3, 236) <= input(13);
output(3, 237) <= input(14);
output(3, 238) <= input(15);
output(3, 239) <= input(32);
output(3, 240) <= input(17);
output(3, 241) <= input(18);
output(3, 242) <= input(19);
output(3, 243) <= input(20);
output(3, 244) <= input(21);
output(3, 245) <= input(22);
output(3, 246) <= input(23);
output(3, 247) <= input(24);
output(3, 248) <= input(25);
output(3, 249) <= input(26);
output(3, 250) <= input(27);
output(3, 251) <= input(28);
output(3, 252) <= input(29);
output(3, 253) <= input(30);
output(3, 254) <= input(31);
output(3, 255) <= input(33);
output(4, 0) <= input(53);
output(4, 1) <= input(51);
output(4, 2) <= input(49);
output(4, 3) <= input(46);
output(4, 4) <= input(47);
output(4, 5) <= input(16);
output(4, 6) <= input(17);
output(4, 7) <= input(18);
output(4, 8) <= input(19);
output(4, 9) <= input(20);
output(4, 10) <= input(21);
output(4, 11) <= input(22);
output(4, 12) <= input(23);
output(4, 13) <= input(24);
output(4, 14) <= input(25);
output(4, 15) <= input(26);
output(4, 16) <= input(54);
output(4, 17) <= input(52);
output(4, 18) <= input(50);
output(4, 19) <= input(48);
output(4, 20) <= input(0);
output(4, 21) <= input(1);
output(4, 22) <= input(2);
output(4, 23) <= input(3);
output(4, 24) <= input(4);
output(4, 25) <= input(5);
output(4, 26) <= input(6);
output(4, 27) <= input(7);
output(4, 28) <= input(8);
output(4, 29) <= input(9);
output(4, 30) <= input(10);
output(4, 31) <= input(11);
output(4, 32) <= input(54);
output(4, 33) <= input(52);
output(4, 34) <= input(50);
output(4, 35) <= input(48);
output(4, 36) <= input(0);
output(4, 37) <= input(1);
output(4, 38) <= input(2);
output(4, 39) <= input(3);
output(4, 40) <= input(4);
output(4, 41) <= input(5);
output(4, 42) <= input(6);
output(4, 43) <= input(7);
output(4, 44) <= input(8);
output(4, 45) <= input(9);
output(4, 46) <= input(10);
output(4, 47) <= input(11);
output(4, 48) <= input(51);
output(4, 49) <= input(49);
output(4, 50) <= input(46);
output(4, 51) <= input(47);
output(4, 52) <= input(16);
output(4, 53) <= input(17);
output(4, 54) <= input(18);
output(4, 55) <= input(19);
output(4, 56) <= input(20);
output(4, 57) <= input(21);
output(4, 58) <= input(22);
output(4, 59) <= input(23);
output(4, 60) <= input(24);
output(4, 61) <= input(25);
output(4, 62) <= input(26);
output(4, 63) <= input(27);
output(4, 64) <= input(51);
output(4, 65) <= input(49);
output(4, 66) <= input(46);
output(4, 67) <= input(47);
output(4, 68) <= input(16);
output(4, 69) <= input(17);
output(4, 70) <= input(18);
output(4, 71) <= input(19);
output(4, 72) <= input(20);
output(4, 73) <= input(21);
output(4, 74) <= input(22);
output(4, 75) <= input(23);
output(4, 76) <= input(24);
output(4, 77) <= input(25);
output(4, 78) <= input(26);
output(4, 79) <= input(27);
output(4, 80) <= input(52);
output(4, 81) <= input(50);
output(4, 82) <= input(48);
output(4, 83) <= input(0);
output(4, 84) <= input(1);
output(4, 85) <= input(2);
output(4, 86) <= input(3);
output(4, 87) <= input(4);
output(4, 88) <= input(5);
output(4, 89) <= input(6);
output(4, 90) <= input(7);
output(4, 91) <= input(8);
output(4, 92) <= input(9);
output(4, 93) <= input(10);
output(4, 94) <= input(11);
output(4, 95) <= input(12);
output(4, 96) <= input(52);
output(4, 97) <= input(50);
output(4, 98) <= input(48);
output(4, 99) <= input(0);
output(4, 100) <= input(1);
output(4, 101) <= input(2);
output(4, 102) <= input(3);
output(4, 103) <= input(4);
output(4, 104) <= input(5);
output(4, 105) <= input(6);
output(4, 106) <= input(7);
output(4, 107) <= input(8);
output(4, 108) <= input(9);
output(4, 109) <= input(10);
output(4, 110) <= input(11);
output(4, 111) <= input(12);
output(4, 112) <= input(49);
output(4, 113) <= input(46);
output(4, 114) <= input(47);
output(4, 115) <= input(16);
output(4, 116) <= input(17);
output(4, 117) <= input(18);
output(4, 118) <= input(19);
output(4, 119) <= input(20);
output(4, 120) <= input(21);
output(4, 121) <= input(22);
output(4, 122) <= input(23);
output(4, 123) <= input(24);
output(4, 124) <= input(25);
output(4, 125) <= input(26);
output(4, 126) <= input(27);
output(4, 127) <= input(28);
output(4, 128) <= input(49);
output(4, 129) <= input(46);
output(4, 130) <= input(47);
output(4, 131) <= input(16);
output(4, 132) <= input(17);
output(4, 133) <= input(18);
output(4, 134) <= input(19);
output(4, 135) <= input(20);
output(4, 136) <= input(21);
output(4, 137) <= input(22);
output(4, 138) <= input(23);
output(4, 139) <= input(24);
output(4, 140) <= input(25);
output(4, 141) <= input(26);
output(4, 142) <= input(27);
output(4, 143) <= input(28);
output(4, 144) <= input(50);
output(4, 145) <= input(48);
output(4, 146) <= input(0);
output(4, 147) <= input(1);
output(4, 148) <= input(2);
output(4, 149) <= input(3);
output(4, 150) <= input(4);
output(4, 151) <= input(5);
output(4, 152) <= input(6);
output(4, 153) <= input(7);
output(4, 154) <= input(8);
output(4, 155) <= input(9);
output(4, 156) <= input(10);
output(4, 157) <= input(11);
output(4, 158) <= input(12);
output(4, 159) <= input(13);
output(4, 160) <= input(50);
output(4, 161) <= input(48);
output(4, 162) <= input(0);
output(4, 163) <= input(1);
output(4, 164) <= input(2);
output(4, 165) <= input(3);
output(4, 166) <= input(4);
output(4, 167) <= input(5);
output(4, 168) <= input(6);
output(4, 169) <= input(7);
output(4, 170) <= input(8);
output(4, 171) <= input(9);
output(4, 172) <= input(10);
output(4, 173) <= input(11);
output(4, 174) <= input(12);
output(4, 175) <= input(13);
output(4, 176) <= input(46);
output(4, 177) <= input(47);
output(4, 178) <= input(16);
output(4, 179) <= input(17);
output(4, 180) <= input(18);
output(4, 181) <= input(19);
output(4, 182) <= input(20);
output(4, 183) <= input(21);
output(4, 184) <= input(22);
output(4, 185) <= input(23);
output(4, 186) <= input(24);
output(4, 187) <= input(25);
output(4, 188) <= input(26);
output(4, 189) <= input(27);
output(4, 190) <= input(28);
output(4, 191) <= input(29);
output(4, 192) <= input(46);
output(4, 193) <= input(47);
output(4, 194) <= input(16);
output(4, 195) <= input(17);
output(4, 196) <= input(18);
output(4, 197) <= input(19);
output(4, 198) <= input(20);
output(4, 199) <= input(21);
output(4, 200) <= input(22);
output(4, 201) <= input(23);
output(4, 202) <= input(24);
output(4, 203) <= input(25);
output(4, 204) <= input(26);
output(4, 205) <= input(27);
output(4, 206) <= input(28);
output(4, 207) <= input(29);
output(4, 208) <= input(48);
output(4, 209) <= input(0);
output(4, 210) <= input(1);
output(4, 211) <= input(2);
output(4, 212) <= input(3);
output(4, 213) <= input(4);
output(4, 214) <= input(5);
output(4, 215) <= input(6);
output(4, 216) <= input(7);
output(4, 217) <= input(8);
output(4, 218) <= input(9);
output(4, 219) <= input(10);
output(4, 220) <= input(11);
output(4, 221) <= input(12);
output(4, 222) <= input(13);
output(4, 223) <= input(14);
output(4, 224) <= input(48);
output(4, 225) <= input(0);
output(4, 226) <= input(1);
output(4, 227) <= input(2);
output(4, 228) <= input(3);
output(4, 229) <= input(4);
output(4, 230) <= input(5);
output(4, 231) <= input(6);
output(4, 232) <= input(7);
output(4, 233) <= input(8);
output(4, 234) <= input(9);
output(4, 235) <= input(10);
output(4, 236) <= input(11);
output(4, 237) <= input(12);
output(4, 238) <= input(13);
output(4, 239) <= input(14);
output(4, 240) <= input(47);
output(4, 241) <= input(16);
output(4, 242) <= input(17);
output(4, 243) <= input(18);
output(4, 244) <= input(19);
output(4, 245) <= input(20);
output(4, 246) <= input(21);
output(4, 247) <= input(22);
output(4, 248) <= input(23);
output(4, 249) <= input(24);
output(4, 250) <= input(25);
output(4, 251) <= input(26);
output(4, 252) <= input(27);
output(4, 253) <= input(28);
output(4, 254) <= input(29);
output(4, 255) <= input(30);
output(5, 0) <= input(55);
output(5, 1) <= input(53);
output(5, 2) <= input(51);
output(5, 3) <= input(49);
output(5, 4) <= input(46);
output(5, 5) <= input(47);
output(5, 6) <= input(16);
output(5, 7) <= input(17);
output(5, 8) <= input(18);
output(5, 9) <= input(19);
output(5, 10) <= input(20);
output(5, 11) <= input(21);
output(5, 12) <= input(22);
output(5, 13) <= input(23);
output(5, 14) <= input(24);
output(5, 15) <= input(25);
output(5, 16) <= input(55);
output(5, 17) <= input(53);
output(5, 18) <= input(51);
output(5, 19) <= input(49);
output(5, 20) <= input(46);
output(5, 21) <= input(47);
output(5, 22) <= input(16);
output(5, 23) <= input(17);
output(5, 24) <= input(18);
output(5, 25) <= input(19);
output(5, 26) <= input(20);
output(5, 27) <= input(21);
output(5, 28) <= input(22);
output(5, 29) <= input(23);
output(5, 30) <= input(24);
output(5, 31) <= input(25);
output(5, 32) <= input(56);
output(5, 33) <= input(54);
output(5, 34) <= input(52);
output(5, 35) <= input(50);
output(5, 36) <= input(48);
output(5, 37) <= input(0);
output(5, 38) <= input(1);
output(5, 39) <= input(2);
output(5, 40) <= input(3);
output(5, 41) <= input(4);
output(5, 42) <= input(5);
output(5, 43) <= input(6);
output(5, 44) <= input(7);
output(5, 45) <= input(8);
output(5, 46) <= input(9);
output(5, 47) <= input(10);
output(5, 48) <= input(56);
output(5, 49) <= input(54);
output(5, 50) <= input(52);
output(5, 51) <= input(50);
output(5, 52) <= input(48);
output(5, 53) <= input(0);
output(5, 54) <= input(1);
output(5, 55) <= input(2);
output(5, 56) <= input(3);
output(5, 57) <= input(4);
output(5, 58) <= input(5);
output(5, 59) <= input(6);
output(5, 60) <= input(7);
output(5, 61) <= input(8);
output(5, 62) <= input(9);
output(5, 63) <= input(10);
output(5, 64) <= input(56);
output(5, 65) <= input(54);
output(5, 66) <= input(52);
output(5, 67) <= input(50);
output(5, 68) <= input(48);
output(5, 69) <= input(0);
output(5, 70) <= input(1);
output(5, 71) <= input(2);
output(5, 72) <= input(3);
output(5, 73) <= input(4);
output(5, 74) <= input(5);
output(5, 75) <= input(6);
output(5, 76) <= input(7);
output(5, 77) <= input(8);
output(5, 78) <= input(9);
output(5, 79) <= input(10);
output(5, 80) <= input(53);
output(5, 81) <= input(51);
output(5, 82) <= input(49);
output(5, 83) <= input(46);
output(5, 84) <= input(47);
output(5, 85) <= input(16);
output(5, 86) <= input(17);
output(5, 87) <= input(18);
output(5, 88) <= input(19);
output(5, 89) <= input(20);
output(5, 90) <= input(21);
output(5, 91) <= input(22);
output(5, 92) <= input(23);
output(5, 93) <= input(24);
output(5, 94) <= input(25);
output(5, 95) <= input(26);
output(5, 96) <= input(53);
output(5, 97) <= input(51);
output(5, 98) <= input(49);
output(5, 99) <= input(46);
output(5, 100) <= input(47);
output(5, 101) <= input(16);
output(5, 102) <= input(17);
output(5, 103) <= input(18);
output(5, 104) <= input(19);
output(5, 105) <= input(20);
output(5, 106) <= input(21);
output(5, 107) <= input(22);
output(5, 108) <= input(23);
output(5, 109) <= input(24);
output(5, 110) <= input(25);
output(5, 111) <= input(26);
output(5, 112) <= input(54);
output(5, 113) <= input(52);
output(5, 114) <= input(50);
output(5, 115) <= input(48);
output(5, 116) <= input(0);
output(5, 117) <= input(1);
output(5, 118) <= input(2);
output(5, 119) <= input(3);
output(5, 120) <= input(4);
output(5, 121) <= input(5);
output(5, 122) <= input(6);
output(5, 123) <= input(7);
output(5, 124) <= input(8);
output(5, 125) <= input(9);
output(5, 126) <= input(10);
output(5, 127) <= input(11);
output(5, 128) <= input(54);
output(5, 129) <= input(52);
output(5, 130) <= input(50);
output(5, 131) <= input(48);
output(5, 132) <= input(0);
output(5, 133) <= input(1);
output(5, 134) <= input(2);
output(5, 135) <= input(3);
output(5, 136) <= input(4);
output(5, 137) <= input(5);
output(5, 138) <= input(6);
output(5, 139) <= input(7);
output(5, 140) <= input(8);
output(5, 141) <= input(9);
output(5, 142) <= input(10);
output(5, 143) <= input(11);
output(5, 144) <= input(54);
output(5, 145) <= input(52);
output(5, 146) <= input(50);
output(5, 147) <= input(48);
output(5, 148) <= input(0);
output(5, 149) <= input(1);
output(5, 150) <= input(2);
output(5, 151) <= input(3);
output(5, 152) <= input(4);
output(5, 153) <= input(5);
output(5, 154) <= input(6);
output(5, 155) <= input(7);
output(5, 156) <= input(8);
output(5, 157) <= input(9);
output(5, 158) <= input(10);
output(5, 159) <= input(11);
output(5, 160) <= input(51);
output(5, 161) <= input(49);
output(5, 162) <= input(46);
output(5, 163) <= input(47);
output(5, 164) <= input(16);
output(5, 165) <= input(17);
output(5, 166) <= input(18);
output(5, 167) <= input(19);
output(5, 168) <= input(20);
output(5, 169) <= input(21);
output(5, 170) <= input(22);
output(5, 171) <= input(23);
output(5, 172) <= input(24);
output(5, 173) <= input(25);
output(5, 174) <= input(26);
output(5, 175) <= input(27);
output(5, 176) <= input(51);
output(5, 177) <= input(49);
output(5, 178) <= input(46);
output(5, 179) <= input(47);
output(5, 180) <= input(16);
output(5, 181) <= input(17);
output(5, 182) <= input(18);
output(5, 183) <= input(19);
output(5, 184) <= input(20);
output(5, 185) <= input(21);
output(5, 186) <= input(22);
output(5, 187) <= input(23);
output(5, 188) <= input(24);
output(5, 189) <= input(25);
output(5, 190) <= input(26);
output(5, 191) <= input(27);
output(5, 192) <= input(51);
output(5, 193) <= input(49);
output(5, 194) <= input(46);
output(5, 195) <= input(47);
output(5, 196) <= input(16);
output(5, 197) <= input(17);
output(5, 198) <= input(18);
output(5, 199) <= input(19);
output(5, 200) <= input(20);
output(5, 201) <= input(21);
output(5, 202) <= input(22);
output(5, 203) <= input(23);
output(5, 204) <= input(24);
output(5, 205) <= input(25);
output(5, 206) <= input(26);
output(5, 207) <= input(27);
output(5, 208) <= input(52);
output(5, 209) <= input(50);
output(5, 210) <= input(48);
output(5, 211) <= input(0);
output(5, 212) <= input(1);
output(5, 213) <= input(2);
output(5, 214) <= input(3);
output(5, 215) <= input(4);
output(5, 216) <= input(5);
output(5, 217) <= input(6);
output(5, 218) <= input(7);
output(5, 219) <= input(8);
output(5, 220) <= input(9);
output(5, 221) <= input(10);
output(5, 222) <= input(11);
output(5, 223) <= input(12);
output(5, 224) <= input(52);
output(5, 225) <= input(50);
output(5, 226) <= input(48);
output(5, 227) <= input(0);
output(5, 228) <= input(1);
output(5, 229) <= input(2);
output(5, 230) <= input(3);
output(5, 231) <= input(4);
output(5, 232) <= input(5);
output(5, 233) <= input(6);
output(5, 234) <= input(7);
output(5, 235) <= input(8);
output(5, 236) <= input(9);
output(5, 237) <= input(10);
output(5, 238) <= input(11);
output(5, 239) <= input(12);
output(5, 240) <= input(49);
output(5, 241) <= input(46);
output(5, 242) <= input(47);
output(5, 243) <= input(16);
output(5, 244) <= input(17);
output(5, 245) <= input(18);
output(5, 246) <= input(19);
output(5, 247) <= input(20);
output(5, 248) <= input(21);
output(5, 249) <= input(22);
output(5, 250) <= input(23);
output(5, 251) <= input(24);
output(5, 252) <= input(25);
output(5, 253) <= input(26);
output(5, 254) <= input(27);
output(5, 255) <= input(28);
when "0010" =>
output(0, 0) <= input(0);
output(0, 1) <= input(1);
output(0, 2) <= input(2);
output(0, 3) <= input(3);
output(0, 4) <= input(4);
output(0, 5) <= input(5);
output(0, 6) <= input(6);
output(0, 7) <= input(7);
output(0, 8) <= input(8);
output(0, 9) <= input(9);
output(0, 10) <= input(10);
output(0, 11) <= input(11);
output(0, 12) <= input(12);
output(0, 13) <= input(13);
output(0, 14) <= input(14);
output(0, 15) <= input(15);
output(0, 16) <= input(0);
output(0, 17) <= input(1);
output(0, 18) <= input(2);
output(0, 19) <= input(3);
output(0, 20) <= input(4);
output(0, 21) <= input(5);
output(0, 22) <= input(6);
output(0, 23) <= input(7);
output(0, 24) <= input(8);
output(0, 25) <= input(9);
output(0, 26) <= input(10);
output(0, 27) <= input(11);
output(0, 28) <= input(12);
output(0, 29) <= input(13);
output(0, 30) <= input(14);
output(0, 31) <= input(15);
output(0, 32) <= input(0);
output(0, 33) <= input(1);
output(0, 34) <= input(2);
output(0, 35) <= input(3);
output(0, 36) <= input(4);
output(0, 37) <= input(5);
output(0, 38) <= input(6);
output(0, 39) <= input(7);
output(0, 40) <= input(8);
output(0, 41) <= input(9);
output(0, 42) <= input(10);
output(0, 43) <= input(11);
output(0, 44) <= input(12);
output(0, 45) <= input(13);
output(0, 46) <= input(14);
output(0, 47) <= input(15);
output(0, 48) <= input(16);
output(0, 49) <= input(17);
output(0, 50) <= input(18);
output(0, 51) <= input(19);
output(0, 52) <= input(20);
output(0, 53) <= input(21);
output(0, 54) <= input(22);
output(0, 55) <= input(23);
output(0, 56) <= input(24);
output(0, 57) <= input(25);
output(0, 58) <= input(26);
output(0, 59) <= input(27);
output(0, 60) <= input(28);
output(0, 61) <= input(29);
output(0, 62) <= input(30);
output(0, 63) <= input(31);
output(0, 64) <= input(16);
output(0, 65) <= input(17);
output(0, 66) <= input(18);
output(0, 67) <= input(19);
output(0, 68) <= input(20);
output(0, 69) <= input(21);
output(0, 70) <= input(22);
output(0, 71) <= input(23);
output(0, 72) <= input(24);
output(0, 73) <= input(25);
output(0, 74) <= input(26);
output(0, 75) <= input(27);
output(0, 76) <= input(28);
output(0, 77) <= input(29);
output(0, 78) <= input(30);
output(0, 79) <= input(31);
output(0, 80) <= input(16);
output(0, 81) <= input(17);
output(0, 82) <= input(18);
output(0, 83) <= input(19);
output(0, 84) <= input(20);
output(0, 85) <= input(21);
output(0, 86) <= input(22);
output(0, 87) <= input(23);
output(0, 88) <= input(24);
output(0, 89) <= input(25);
output(0, 90) <= input(26);
output(0, 91) <= input(27);
output(0, 92) <= input(28);
output(0, 93) <= input(29);
output(0, 94) <= input(30);
output(0, 95) <= input(31);
output(0, 96) <= input(16);
output(0, 97) <= input(17);
output(0, 98) <= input(18);
output(0, 99) <= input(19);
output(0, 100) <= input(20);
output(0, 101) <= input(21);
output(0, 102) <= input(22);
output(0, 103) <= input(23);
output(0, 104) <= input(24);
output(0, 105) <= input(25);
output(0, 106) <= input(26);
output(0, 107) <= input(27);
output(0, 108) <= input(28);
output(0, 109) <= input(29);
output(0, 110) <= input(30);
output(0, 111) <= input(31);
output(0, 112) <= input(1);
output(0, 113) <= input(2);
output(0, 114) <= input(3);
output(0, 115) <= input(4);
output(0, 116) <= input(5);
output(0, 117) <= input(6);
output(0, 118) <= input(7);
output(0, 119) <= input(8);
output(0, 120) <= input(9);
output(0, 121) <= input(10);
output(0, 122) <= input(11);
output(0, 123) <= input(12);
output(0, 124) <= input(13);
output(0, 125) <= input(14);
output(0, 126) <= input(15);
output(0, 127) <= input(32);
output(0, 128) <= input(1);
output(0, 129) <= input(2);
output(0, 130) <= input(3);
output(0, 131) <= input(4);
output(0, 132) <= input(5);
output(0, 133) <= input(6);
output(0, 134) <= input(7);
output(0, 135) <= input(8);
output(0, 136) <= input(9);
output(0, 137) <= input(10);
output(0, 138) <= input(11);
output(0, 139) <= input(12);
output(0, 140) <= input(13);
output(0, 141) <= input(14);
output(0, 142) <= input(15);
output(0, 143) <= input(32);
output(0, 144) <= input(1);
output(0, 145) <= input(2);
output(0, 146) <= input(3);
output(0, 147) <= input(4);
output(0, 148) <= input(5);
output(0, 149) <= input(6);
output(0, 150) <= input(7);
output(0, 151) <= input(8);
output(0, 152) <= input(9);
output(0, 153) <= input(10);
output(0, 154) <= input(11);
output(0, 155) <= input(12);
output(0, 156) <= input(13);
output(0, 157) <= input(14);
output(0, 158) <= input(15);
output(0, 159) <= input(32);
output(0, 160) <= input(1);
output(0, 161) <= input(2);
output(0, 162) <= input(3);
output(0, 163) <= input(4);
output(0, 164) <= input(5);
output(0, 165) <= input(6);
output(0, 166) <= input(7);
output(0, 167) <= input(8);
output(0, 168) <= input(9);
output(0, 169) <= input(10);
output(0, 170) <= input(11);
output(0, 171) <= input(12);
output(0, 172) <= input(13);
output(0, 173) <= input(14);
output(0, 174) <= input(15);
output(0, 175) <= input(32);
output(0, 176) <= input(17);
output(0, 177) <= input(18);
output(0, 178) <= input(19);
output(0, 179) <= input(20);
output(0, 180) <= input(21);
output(0, 181) <= input(22);
output(0, 182) <= input(23);
output(0, 183) <= input(24);
output(0, 184) <= input(25);
output(0, 185) <= input(26);
output(0, 186) <= input(27);
output(0, 187) <= input(28);
output(0, 188) <= input(29);
output(0, 189) <= input(30);
output(0, 190) <= input(31);
output(0, 191) <= input(33);
output(0, 192) <= input(17);
output(0, 193) <= input(18);
output(0, 194) <= input(19);
output(0, 195) <= input(20);
output(0, 196) <= input(21);
output(0, 197) <= input(22);
output(0, 198) <= input(23);
output(0, 199) <= input(24);
output(0, 200) <= input(25);
output(0, 201) <= input(26);
output(0, 202) <= input(27);
output(0, 203) <= input(28);
output(0, 204) <= input(29);
output(0, 205) <= input(30);
output(0, 206) <= input(31);
output(0, 207) <= input(33);
output(0, 208) <= input(17);
output(0, 209) <= input(18);
output(0, 210) <= input(19);
output(0, 211) <= input(20);
output(0, 212) <= input(21);
output(0, 213) <= input(22);
output(0, 214) <= input(23);
output(0, 215) <= input(24);
output(0, 216) <= input(25);
output(0, 217) <= input(26);
output(0, 218) <= input(27);
output(0, 219) <= input(28);
output(0, 220) <= input(29);
output(0, 221) <= input(30);
output(0, 222) <= input(31);
output(0, 223) <= input(33);
output(0, 224) <= input(17);
output(0, 225) <= input(18);
output(0, 226) <= input(19);
output(0, 227) <= input(20);
output(0, 228) <= input(21);
output(0, 229) <= input(22);
output(0, 230) <= input(23);
output(0, 231) <= input(24);
output(0, 232) <= input(25);
output(0, 233) <= input(26);
output(0, 234) <= input(27);
output(0, 235) <= input(28);
output(0, 236) <= input(29);
output(0, 237) <= input(30);
output(0, 238) <= input(31);
output(0, 239) <= input(33);
output(0, 240) <= input(2);
output(0, 241) <= input(3);
output(0, 242) <= input(4);
output(0, 243) <= input(5);
output(0, 244) <= input(6);
output(0, 245) <= input(7);
output(0, 246) <= input(8);
output(0, 247) <= input(9);
output(0, 248) <= input(10);
output(0, 249) <= input(11);
output(0, 250) <= input(12);
output(0, 251) <= input(13);
output(0, 252) <= input(14);
output(0, 253) <= input(15);
output(0, 254) <= input(32);
output(0, 255) <= input(34);
output(1, 0) <= input(35);
output(1, 1) <= input(16);
output(1, 2) <= input(17);
output(1, 3) <= input(18);
output(1, 4) <= input(19);
output(1, 5) <= input(20);
output(1, 6) <= input(21);
output(1, 7) <= input(22);
output(1, 8) <= input(23);
output(1, 9) <= input(24);
output(1, 10) <= input(25);
output(1, 11) <= input(26);
output(1, 12) <= input(27);
output(1, 13) <= input(28);
output(1, 14) <= input(29);
output(1, 15) <= input(30);
output(1, 16) <= input(35);
output(1, 17) <= input(16);
output(1, 18) <= input(17);
output(1, 19) <= input(18);
output(1, 20) <= input(19);
output(1, 21) <= input(20);
output(1, 22) <= input(21);
output(1, 23) <= input(22);
output(1, 24) <= input(23);
output(1, 25) <= input(24);
output(1, 26) <= input(25);
output(1, 27) <= input(26);
output(1, 28) <= input(27);
output(1, 29) <= input(28);
output(1, 30) <= input(29);
output(1, 31) <= input(30);
output(1, 32) <= input(35);
output(1, 33) <= input(16);
output(1, 34) <= input(17);
output(1, 35) <= input(18);
output(1, 36) <= input(19);
output(1, 37) <= input(20);
output(1, 38) <= input(21);
output(1, 39) <= input(22);
output(1, 40) <= input(23);
output(1, 41) <= input(24);
output(1, 42) <= input(25);
output(1, 43) <= input(26);
output(1, 44) <= input(27);
output(1, 45) <= input(28);
output(1, 46) <= input(29);
output(1, 47) <= input(30);
output(1, 48) <= input(35);
output(1, 49) <= input(16);
output(1, 50) <= input(17);
output(1, 51) <= input(18);
output(1, 52) <= input(19);
output(1, 53) <= input(20);
output(1, 54) <= input(21);
output(1, 55) <= input(22);
output(1, 56) <= input(23);
output(1, 57) <= input(24);
output(1, 58) <= input(25);
output(1, 59) <= input(26);
output(1, 60) <= input(27);
output(1, 61) <= input(28);
output(1, 62) <= input(29);
output(1, 63) <= input(30);
output(1, 64) <= input(35);
output(1, 65) <= input(16);
output(1, 66) <= input(17);
output(1, 67) <= input(18);
output(1, 68) <= input(19);
output(1, 69) <= input(20);
output(1, 70) <= input(21);
output(1, 71) <= input(22);
output(1, 72) <= input(23);
output(1, 73) <= input(24);
output(1, 74) <= input(25);
output(1, 75) <= input(26);
output(1, 76) <= input(27);
output(1, 77) <= input(28);
output(1, 78) <= input(29);
output(1, 79) <= input(30);
output(1, 80) <= input(0);
output(1, 81) <= input(1);
output(1, 82) <= input(2);
output(1, 83) <= input(3);
output(1, 84) <= input(4);
output(1, 85) <= input(5);
output(1, 86) <= input(6);
output(1, 87) <= input(7);
output(1, 88) <= input(8);
output(1, 89) <= input(9);
output(1, 90) <= input(10);
output(1, 91) <= input(11);
output(1, 92) <= input(12);
output(1, 93) <= input(13);
output(1, 94) <= input(14);
output(1, 95) <= input(15);
output(1, 96) <= input(0);
output(1, 97) <= input(1);
output(1, 98) <= input(2);
output(1, 99) <= input(3);
output(1, 100) <= input(4);
output(1, 101) <= input(5);
output(1, 102) <= input(6);
output(1, 103) <= input(7);
output(1, 104) <= input(8);
output(1, 105) <= input(9);
output(1, 106) <= input(10);
output(1, 107) <= input(11);
output(1, 108) <= input(12);
output(1, 109) <= input(13);
output(1, 110) <= input(14);
output(1, 111) <= input(15);
output(1, 112) <= input(0);
output(1, 113) <= input(1);
output(1, 114) <= input(2);
output(1, 115) <= input(3);
output(1, 116) <= input(4);
output(1, 117) <= input(5);
output(1, 118) <= input(6);
output(1, 119) <= input(7);
output(1, 120) <= input(8);
output(1, 121) <= input(9);
output(1, 122) <= input(10);
output(1, 123) <= input(11);
output(1, 124) <= input(12);
output(1, 125) <= input(13);
output(1, 126) <= input(14);
output(1, 127) <= input(15);
output(1, 128) <= input(0);
output(1, 129) <= input(1);
output(1, 130) <= input(2);
output(1, 131) <= input(3);
output(1, 132) <= input(4);
output(1, 133) <= input(5);
output(1, 134) <= input(6);
output(1, 135) <= input(7);
output(1, 136) <= input(8);
output(1, 137) <= input(9);
output(1, 138) <= input(10);
output(1, 139) <= input(11);
output(1, 140) <= input(12);
output(1, 141) <= input(13);
output(1, 142) <= input(14);
output(1, 143) <= input(15);
output(1, 144) <= input(0);
output(1, 145) <= input(1);
output(1, 146) <= input(2);
output(1, 147) <= input(3);
output(1, 148) <= input(4);
output(1, 149) <= input(5);
output(1, 150) <= input(6);
output(1, 151) <= input(7);
output(1, 152) <= input(8);
output(1, 153) <= input(9);
output(1, 154) <= input(10);
output(1, 155) <= input(11);
output(1, 156) <= input(12);
output(1, 157) <= input(13);
output(1, 158) <= input(14);
output(1, 159) <= input(15);
output(1, 160) <= input(16);
output(1, 161) <= input(17);
output(1, 162) <= input(18);
output(1, 163) <= input(19);
output(1, 164) <= input(20);
output(1, 165) <= input(21);
output(1, 166) <= input(22);
output(1, 167) <= input(23);
output(1, 168) <= input(24);
output(1, 169) <= input(25);
output(1, 170) <= input(26);
output(1, 171) <= input(27);
output(1, 172) <= input(28);
output(1, 173) <= input(29);
output(1, 174) <= input(30);
output(1, 175) <= input(31);
output(1, 176) <= input(16);
output(1, 177) <= input(17);
output(1, 178) <= input(18);
output(1, 179) <= input(19);
output(1, 180) <= input(20);
output(1, 181) <= input(21);
output(1, 182) <= input(22);
output(1, 183) <= input(23);
output(1, 184) <= input(24);
output(1, 185) <= input(25);
output(1, 186) <= input(26);
output(1, 187) <= input(27);
output(1, 188) <= input(28);
output(1, 189) <= input(29);
output(1, 190) <= input(30);
output(1, 191) <= input(31);
output(1, 192) <= input(16);
output(1, 193) <= input(17);
output(1, 194) <= input(18);
output(1, 195) <= input(19);
output(1, 196) <= input(20);
output(1, 197) <= input(21);
output(1, 198) <= input(22);
output(1, 199) <= input(23);
output(1, 200) <= input(24);
output(1, 201) <= input(25);
output(1, 202) <= input(26);
output(1, 203) <= input(27);
output(1, 204) <= input(28);
output(1, 205) <= input(29);
output(1, 206) <= input(30);
output(1, 207) <= input(31);
output(1, 208) <= input(16);
output(1, 209) <= input(17);
output(1, 210) <= input(18);
output(1, 211) <= input(19);
output(1, 212) <= input(20);
output(1, 213) <= input(21);
output(1, 214) <= input(22);
output(1, 215) <= input(23);
output(1, 216) <= input(24);
output(1, 217) <= input(25);
output(1, 218) <= input(26);
output(1, 219) <= input(27);
output(1, 220) <= input(28);
output(1, 221) <= input(29);
output(1, 222) <= input(30);
output(1, 223) <= input(31);
output(1, 224) <= input(16);
output(1, 225) <= input(17);
output(1, 226) <= input(18);
output(1, 227) <= input(19);
output(1, 228) <= input(20);
output(1, 229) <= input(21);
output(1, 230) <= input(22);
output(1, 231) <= input(23);
output(1, 232) <= input(24);
output(1, 233) <= input(25);
output(1, 234) <= input(26);
output(1, 235) <= input(27);
output(1, 236) <= input(28);
output(1, 237) <= input(29);
output(1, 238) <= input(30);
output(1, 239) <= input(31);
output(1, 240) <= input(1);
output(1, 241) <= input(2);
output(1, 242) <= input(3);
output(1, 243) <= input(4);
output(1, 244) <= input(5);
output(1, 245) <= input(6);
output(1, 246) <= input(7);
output(1, 247) <= input(8);
output(1, 248) <= input(9);
output(1, 249) <= input(10);
output(1, 250) <= input(11);
output(1, 251) <= input(12);
output(1, 252) <= input(13);
output(1, 253) <= input(14);
output(1, 254) <= input(15);
output(1, 255) <= input(32);
output(2, 0) <= input(36);
output(2, 1) <= input(0);
output(2, 2) <= input(1);
output(2, 3) <= input(2);
output(2, 4) <= input(3);
output(2, 5) <= input(4);
output(2, 6) <= input(5);
output(2, 7) <= input(6);
output(2, 8) <= input(7);
output(2, 9) <= input(8);
output(2, 10) <= input(9);
output(2, 11) <= input(10);
output(2, 12) <= input(11);
output(2, 13) <= input(12);
output(2, 14) <= input(13);
output(2, 15) <= input(14);
output(2, 16) <= input(36);
output(2, 17) <= input(0);
output(2, 18) <= input(1);
output(2, 19) <= input(2);
output(2, 20) <= input(3);
output(2, 21) <= input(4);
output(2, 22) <= input(5);
output(2, 23) <= input(6);
output(2, 24) <= input(7);
output(2, 25) <= input(8);
output(2, 26) <= input(9);
output(2, 27) <= input(10);
output(2, 28) <= input(11);
output(2, 29) <= input(12);
output(2, 30) <= input(13);
output(2, 31) <= input(14);
output(2, 32) <= input(36);
output(2, 33) <= input(0);
output(2, 34) <= input(1);
output(2, 35) <= input(2);
output(2, 36) <= input(3);
output(2, 37) <= input(4);
output(2, 38) <= input(5);
output(2, 39) <= input(6);
output(2, 40) <= input(7);
output(2, 41) <= input(8);
output(2, 42) <= input(9);
output(2, 43) <= input(10);
output(2, 44) <= input(11);
output(2, 45) <= input(12);
output(2, 46) <= input(13);
output(2, 47) <= input(14);
output(2, 48) <= input(36);
output(2, 49) <= input(0);
output(2, 50) <= input(1);
output(2, 51) <= input(2);
output(2, 52) <= input(3);
output(2, 53) <= input(4);
output(2, 54) <= input(5);
output(2, 55) <= input(6);
output(2, 56) <= input(7);
output(2, 57) <= input(8);
output(2, 58) <= input(9);
output(2, 59) <= input(10);
output(2, 60) <= input(11);
output(2, 61) <= input(12);
output(2, 62) <= input(13);
output(2, 63) <= input(14);
output(2, 64) <= input(36);
output(2, 65) <= input(0);
output(2, 66) <= input(1);
output(2, 67) <= input(2);
output(2, 68) <= input(3);
output(2, 69) <= input(4);
output(2, 70) <= input(5);
output(2, 71) <= input(6);
output(2, 72) <= input(7);
output(2, 73) <= input(8);
output(2, 74) <= input(9);
output(2, 75) <= input(10);
output(2, 76) <= input(11);
output(2, 77) <= input(12);
output(2, 78) <= input(13);
output(2, 79) <= input(14);
output(2, 80) <= input(36);
output(2, 81) <= input(0);
output(2, 82) <= input(1);
output(2, 83) <= input(2);
output(2, 84) <= input(3);
output(2, 85) <= input(4);
output(2, 86) <= input(5);
output(2, 87) <= input(6);
output(2, 88) <= input(7);
output(2, 89) <= input(8);
output(2, 90) <= input(9);
output(2, 91) <= input(10);
output(2, 92) <= input(11);
output(2, 93) <= input(12);
output(2, 94) <= input(13);
output(2, 95) <= input(14);
output(2, 96) <= input(36);
output(2, 97) <= input(0);
output(2, 98) <= input(1);
output(2, 99) <= input(2);
output(2, 100) <= input(3);
output(2, 101) <= input(4);
output(2, 102) <= input(5);
output(2, 103) <= input(6);
output(2, 104) <= input(7);
output(2, 105) <= input(8);
output(2, 106) <= input(9);
output(2, 107) <= input(10);
output(2, 108) <= input(11);
output(2, 109) <= input(12);
output(2, 110) <= input(13);
output(2, 111) <= input(14);
output(2, 112) <= input(35);
output(2, 113) <= input(16);
output(2, 114) <= input(17);
output(2, 115) <= input(18);
output(2, 116) <= input(19);
output(2, 117) <= input(20);
output(2, 118) <= input(21);
output(2, 119) <= input(22);
output(2, 120) <= input(23);
output(2, 121) <= input(24);
output(2, 122) <= input(25);
output(2, 123) <= input(26);
output(2, 124) <= input(27);
output(2, 125) <= input(28);
output(2, 126) <= input(29);
output(2, 127) <= input(30);
output(2, 128) <= input(35);
output(2, 129) <= input(16);
output(2, 130) <= input(17);
output(2, 131) <= input(18);
output(2, 132) <= input(19);
output(2, 133) <= input(20);
output(2, 134) <= input(21);
output(2, 135) <= input(22);
output(2, 136) <= input(23);
output(2, 137) <= input(24);
output(2, 138) <= input(25);
output(2, 139) <= input(26);
output(2, 140) <= input(27);
output(2, 141) <= input(28);
output(2, 142) <= input(29);
output(2, 143) <= input(30);
output(2, 144) <= input(35);
output(2, 145) <= input(16);
output(2, 146) <= input(17);
output(2, 147) <= input(18);
output(2, 148) <= input(19);
output(2, 149) <= input(20);
output(2, 150) <= input(21);
output(2, 151) <= input(22);
output(2, 152) <= input(23);
output(2, 153) <= input(24);
output(2, 154) <= input(25);
output(2, 155) <= input(26);
output(2, 156) <= input(27);
output(2, 157) <= input(28);
output(2, 158) <= input(29);
output(2, 159) <= input(30);
output(2, 160) <= input(35);
output(2, 161) <= input(16);
output(2, 162) <= input(17);
output(2, 163) <= input(18);
output(2, 164) <= input(19);
output(2, 165) <= input(20);
output(2, 166) <= input(21);
output(2, 167) <= input(22);
output(2, 168) <= input(23);
output(2, 169) <= input(24);
output(2, 170) <= input(25);
output(2, 171) <= input(26);
output(2, 172) <= input(27);
output(2, 173) <= input(28);
output(2, 174) <= input(29);
output(2, 175) <= input(30);
output(2, 176) <= input(35);
output(2, 177) <= input(16);
output(2, 178) <= input(17);
output(2, 179) <= input(18);
output(2, 180) <= input(19);
output(2, 181) <= input(20);
output(2, 182) <= input(21);
output(2, 183) <= input(22);
output(2, 184) <= input(23);
output(2, 185) <= input(24);
output(2, 186) <= input(25);
output(2, 187) <= input(26);
output(2, 188) <= input(27);
output(2, 189) <= input(28);
output(2, 190) <= input(29);
output(2, 191) <= input(30);
output(2, 192) <= input(35);
output(2, 193) <= input(16);
output(2, 194) <= input(17);
output(2, 195) <= input(18);
output(2, 196) <= input(19);
output(2, 197) <= input(20);
output(2, 198) <= input(21);
output(2, 199) <= input(22);
output(2, 200) <= input(23);
output(2, 201) <= input(24);
output(2, 202) <= input(25);
output(2, 203) <= input(26);
output(2, 204) <= input(27);
output(2, 205) <= input(28);
output(2, 206) <= input(29);
output(2, 207) <= input(30);
output(2, 208) <= input(35);
output(2, 209) <= input(16);
output(2, 210) <= input(17);
output(2, 211) <= input(18);
output(2, 212) <= input(19);
output(2, 213) <= input(20);
output(2, 214) <= input(21);
output(2, 215) <= input(22);
output(2, 216) <= input(23);
output(2, 217) <= input(24);
output(2, 218) <= input(25);
output(2, 219) <= input(26);
output(2, 220) <= input(27);
output(2, 221) <= input(28);
output(2, 222) <= input(29);
output(2, 223) <= input(30);
output(2, 224) <= input(35);
output(2, 225) <= input(16);
output(2, 226) <= input(17);
output(2, 227) <= input(18);
output(2, 228) <= input(19);
output(2, 229) <= input(20);
output(2, 230) <= input(21);
output(2, 231) <= input(22);
output(2, 232) <= input(23);
output(2, 233) <= input(24);
output(2, 234) <= input(25);
output(2, 235) <= input(26);
output(2, 236) <= input(27);
output(2, 237) <= input(28);
output(2, 238) <= input(29);
output(2, 239) <= input(30);
output(2, 240) <= input(0);
output(2, 241) <= input(1);
output(2, 242) <= input(2);
output(2, 243) <= input(3);
output(2, 244) <= input(4);
output(2, 245) <= input(5);
output(2, 246) <= input(6);
output(2, 247) <= input(7);
output(2, 248) <= input(8);
output(2, 249) <= input(9);
output(2, 250) <= input(10);
output(2, 251) <= input(11);
output(2, 252) <= input(12);
output(2, 253) <= input(13);
output(2, 254) <= input(14);
output(2, 255) <= input(15);
output(3, 0) <= input(37);
output(3, 1) <= input(35);
output(3, 2) <= input(16);
output(3, 3) <= input(17);
output(3, 4) <= input(18);
output(3, 5) <= input(19);
output(3, 6) <= input(20);
output(3, 7) <= input(21);
output(3, 8) <= input(22);
output(3, 9) <= input(23);
output(3, 10) <= input(24);
output(3, 11) <= input(25);
output(3, 12) <= input(26);
output(3, 13) <= input(27);
output(3, 14) <= input(28);
output(3, 15) <= input(29);
output(3, 16) <= input(37);
output(3, 17) <= input(35);
output(3, 18) <= input(16);
output(3, 19) <= input(17);
output(3, 20) <= input(18);
output(3, 21) <= input(19);
output(3, 22) <= input(20);
output(3, 23) <= input(21);
output(3, 24) <= input(22);
output(3, 25) <= input(23);
output(3, 26) <= input(24);
output(3, 27) <= input(25);
output(3, 28) <= input(26);
output(3, 29) <= input(27);
output(3, 30) <= input(28);
output(3, 31) <= input(29);
output(3, 32) <= input(37);
output(3, 33) <= input(35);
output(3, 34) <= input(16);
output(3, 35) <= input(17);
output(3, 36) <= input(18);
output(3, 37) <= input(19);
output(3, 38) <= input(20);
output(3, 39) <= input(21);
output(3, 40) <= input(22);
output(3, 41) <= input(23);
output(3, 42) <= input(24);
output(3, 43) <= input(25);
output(3, 44) <= input(26);
output(3, 45) <= input(27);
output(3, 46) <= input(28);
output(3, 47) <= input(29);
output(3, 48) <= input(37);
output(3, 49) <= input(35);
output(3, 50) <= input(16);
output(3, 51) <= input(17);
output(3, 52) <= input(18);
output(3, 53) <= input(19);
output(3, 54) <= input(20);
output(3, 55) <= input(21);
output(3, 56) <= input(22);
output(3, 57) <= input(23);
output(3, 58) <= input(24);
output(3, 59) <= input(25);
output(3, 60) <= input(26);
output(3, 61) <= input(27);
output(3, 62) <= input(28);
output(3, 63) <= input(29);
output(3, 64) <= input(37);
output(3, 65) <= input(35);
output(3, 66) <= input(16);
output(3, 67) <= input(17);
output(3, 68) <= input(18);
output(3, 69) <= input(19);
output(3, 70) <= input(20);
output(3, 71) <= input(21);
output(3, 72) <= input(22);
output(3, 73) <= input(23);
output(3, 74) <= input(24);
output(3, 75) <= input(25);
output(3, 76) <= input(26);
output(3, 77) <= input(27);
output(3, 78) <= input(28);
output(3, 79) <= input(29);
output(3, 80) <= input(37);
output(3, 81) <= input(35);
output(3, 82) <= input(16);
output(3, 83) <= input(17);
output(3, 84) <= input(18);
output(3, 85) <= input(19);
output(3, 86) <= input(20);
output(3, 87) <= input(21);
output(3, 88) <= input(22);
output(3, 89) <= input(23);
output(3, 90) <= input(24);
output(3, 91) <= input(25);
output(3, 92) <= input(26);
output(3, 93) <= input(27);
output(3, 94) <= input(28);
output(3, 95) <= input(29);
output(3, 96) <= input(37);
output(3, 97) <= input(35);
output(3, 98) <= input(16);
output(3, 99) <= input(17);
output(3, 100) <= input(18);
output(3, 101) <= input(19);
output(3, 102) <= input(20);
output(3, 103) <= input(21);
output(3, 104) <= input(22);
output(3, 105) <= input(23);
output(3, 106) <= input(24);
output(3, 107) <= input(25);
output(3, 108) <= input(26);
output(3, 109) <= input(27);
output(3, 110) <= input(28);
output(3, 111) <= input(29);
output(3, 112) <= input(37);
output(3, 113) <= input(35);
output(3, 114) <= input(16);
output(3, 115) <= input(17);
output(3, 116) <= input(18);
output(3, 117) <= input(19);
output(3, 118) <= input(20);
output(3, 119) <= input(21);
output(3, 120) <= input(22);
output(3, 121) <= input(23);
output(3, 122) <= input(24);
output(3, 123) <= input(25);
output(3, 124) <= input(26);
output(3, 125) <= input(27);
output(3, 126) <= input(28);
output(3, 127) <= input(29);
output(3, 128) <= input(37);
output(3, 129) <= input(35);
output(3, 130) <= input(16);
output(3, 131) <= input(17);
output(3, 132) <= input(18);
output(3, 133) <= input(19);
output(3, 134) <= input(20);
output(3, 135) <= input(21);
output(3, 136) <= input(22);
output(3, 137) <= input(23);
output(3, 138) <= input(24);
output(3, 139) <= input(25);
output(3, 140) <= input(26);
output(3, 141) <= input(27);
output(3, 142) <= input(28);
output(3, 143) <= input(29);
output(3, 144) <= input(37);
output(3, 145) <= input(35);
output(3, 146) <= input(16);
output(3, 147) <= input(17);
output(3, 148) <= input(18);
output(3, 149) <= input(19);
output(3, 150) <= input(20);
output(3, 151) <= input(21);
output(3, 152) <= input(22);
output(3, 153) <= input(23);
output(3, 154) <= input(24);
output(3, 155) <= input(25);
output(3, 156) <= input(26);
output(3, 157) <= input(27);
output(3, 158) <= input(28);
output(3, 159) <= input(29);
output(3, 160) <= input(37);
output(3, 161) <= input(35);
output(3, 162) <= input(16);
output(3, 163) <= input(17);
output(3, 164) <= input(18);
output(3, 165) <= input(19);
output(3, 166) <= input(20);
output(3, 167) <= input(21);
output(3, 168) <= input(22);
output(3, 169) <= input(23);
output(3, 170) <= input(24);
output(3, 171) <= input(25);
output(3, 172) <= input(26);
output(3, 173) <= input(27);
output(3, 174) <= input(28);
output(3, 175) <= input(29);
output(3, 176) <= input(37);
output(3, 177) <= input(35);
output(3, 178) <= input(16);
output(3, 179) <= input(17);
output(3, 180) <= input(18);
output(3, 181) <= input(19);
output(3, 182) <= input(20);
output(3, 183) <= input(21);
output(3, 184) <= input(22);
output(3, 185) <= input(23);
output(3, 186) <= input(24);
output(3, 187) <= input(25);
output(3, 188) <= input(26);
output(3, 189) <= input(27);
output(3, 190) <= input(28);
output(3, 191) <= input(29);
output(3, 192) <= input(37);
output(3, 193) <= input(35);
output(3, 194) <= input(16);
output(3, 195) <= input(17);
output(3, 196) <= input(18);
output(3, 197) <= input(19);
output(3, 198) <= input(20);
output(3, 199) <= input(21);
output(3, 200) <= input(22);
output(3, 201) <= input(23);
output(3, 202) <= input(24);
output(3, 203) <= input(25);
output(3, 204) <= input(26);
output(3, 205) <= input(27);
output(3, 206) <= input(28);
output(3, 207) <= input(29);
output(3, 208) <= input(37);
output(3, 209) <= input(35);
output(3, 210) <= input(16);
output(3, 211) <= input(17);
output(3, 212) <= input(18);
output(3, 213) <= input(19);
output(3, 214) <= input(20);
output(3, 215) <= input(21);
output(3, 216) <= input(22);
output(3, 217) <= input(23);
output(3, 218) <= input(24);
output(3, 219) <= input(25);
output(3, 220) <= input(26);
output(3, 221) <= input(27);
output(3, 222) <= input(28);
output(3, 223) <= input(29);
output(3, 224) <= input(37);
output(3, 225) <= input(35);
output(3, 226) <= input(16);
output(3, 227) <= input(17);
output(3, 228) <= input(18);
output(3, 229) <= input(19);
output(3, 230) <= input(20);
output(3, 231) <= input(21);
output(3, 232) <= input(22);
output(3, 233) <= input(23);
output(3, 234) <= input(24);
output(3, 235) <= input(25);
output(3, 236) <= input(26);
output(3, 237) <= input(27);
output(3, 238) <= input(28);
output(3, 239) <= input(29);
output(3, 240) <= input(36);
output(3, 241) <= input(0);
output(3, 242) <= input(1);
output(3, 243) <= input(2);
output(3, 244) <= input(3);
output(3, 245) <= input(4);
output(3, 246) <= input(5);
output(3, 247) <= input(6);
output(3, 248) <= input(7);
output(3, 249) <= input(8);
output(3, 250) <= input(9);
output(3, 251) <= input(10);
output(3, 252) <= input(11);
output(3, 253) <= input(12);
output(3, 254) <= input(13);
output(3, 255) <= input(14);
output(4, 0) <= input(38);
output(4, 1) <= input(36);
output(4, 2) <= input(0);
output(4, 3) <= input(1);
output(4, 4) <= input(2);
output(4, 5) <= input(3);
output(4, 6) <= input(4);
output(4, 7) <= input(5);
output(4, 8) <= input(6);
output(4, 9) <= input(7);
output(4, 10) <= input(8);
output(4, 11) <= input(9);
output(4, 12) <= input(10);
output(4, 13) <= input(11);
output(4, 14) <= input(12);
output(4, 15) <= input(13);
output(4, 16) <= input(38);
output(4, 17) <= input(36);
output(4, 18) <= input(0);
output(4, 19) <= input(1);
output(4, 20) <= input(2);
output(4, 21) <= input(3);
output(4, 22) <= input(4);
output(4, 23) <= input(5);
output(4, 24) <= input(6);
output(4, 25) <= input(7);
output(4, 26) <= input(8);
output(4, 27) <= input(9);
output(4, 28) <= input(10);
output(4, 29) <= input(11);
output(4, 30) <= input(12);
output(4, 31) <= input(13);
output(4, 32) <= input(38);
output(4, 33) <= input(36);
output(4, 34) <= input(0);
output(4, 35) <= input(1);
output(4, 36) <= input(2);
output(4, 37) <= input(3);
output(4, 38) <= input(4);
output(4, 39) <= input(5);
output(4, 40) <= input(6);
output(4, 41) <= input(7);
output(4, 42) <= input(8);
output(4, 43) <= input(9);
output(4, 44) <= input(10);
output(4, 45) <= input(11);
output(4, 46) <= input(12);
output(4, 47) <= input(13);
output(4, 48) <= input(38);
output(4, 49) <= input(36);
output(4, 50) <= input(0);
output(4, 51) <= input(1);
output(4, 52) <= input(2);
output(4, 53) <= input(3);
output(4, 54) <= input(4);
output(4, 55) <= input(5);
output(4, 56) <= input(6);
output(4, 57) <= input(7);
output(4, 58) <= input(8);
output(4, 59) <= input(9);
output(4, 60) <= input(10);
output(4, 61) <= input(11);
output(4, 62) <= input(12);
output(4, 63) <= input(13);
output(4, 64) <= input(38);
output(4, 65) <= input(36);
output(4, 66) <= input(0);
output(4, 67) <= input(1);
output(4, 68) <= input(2);
output(4, 69) <= input(3);
output(4, 70) <= input(4);
output(4, 71) <= input(5);
output(4, 72) <= input(6);
output(4, 73) <= input(7);
output(4, 74) <= input(8);
output(4, 75) <= input(9);
output(4, 76) <= input(10);
output(4, 77) <= input(11);
output(4, 78) <= input(12);
output(4, 79) <= input(13);
output(4, 80) <= input(38);
output(4, 81) <= input(36);
output(4, 82) <= input(0);
output(4, 83) <= input(1);
output(4, 84) <= input(2);
output(4, 85) <= input(3);
output(4, 86) <= input(4);
output(4, 87) <= input(5);
output(4, 88) <= input(6);
output(4, 89) <= input(7);
output(4, 90) <= input(8);
output(4, 91) <= input(9);
output(4, 92) <= input(10);
output(4, 93) <= input(11);
output(4, 94) <= input(12);
output(4, 95) <= input(13);
output(4, 96) <= input(38);
output(4, 97) <= input(36);
output(4, 98) <= input(0);
output(4, 99) <= input(1);
output(4, 100) <= input(2);
output(4, 101) <= input(3);
output(4, 102) <= input(4);
output(4, 103) <= input(5);
output(4, 104) <= input(6);
output(4, 105) <= input(7);
output(4, 106) <= input(8);
output(4, 107) <= input(9);
output(4, 108) <= input(10);
output(4, 109) <= input(11);
output(4, 110) <= input(12);
output(4, 111) <= input(13);
output(4, 112) <= input(38);
output(4, 113) <= input(36);
output(4, 114) <= input(0);
output(4, 115) <= input(1);
output(4, 116) <= input(2);
output(4, 117) <= input(3);
output(4, 118) <= input(4);
output(4, 119) <= input(5);
output(4, 120) <= input(6);
output(4, 121) <= input(7);
output(4, 122) <= input(8);
output(4, 123) <= input(9);
output(4, 124) <= input(10);
output(4, 125) <= input(11);
output(4, 126) <= input(12);
output(4, 127) <= input(13);
output(4, 128) <= input(38);
output(4, 129) <= input(36);
output(4, 130) <= input(0);
output(4, 131) <= input(1);
output(4, 132) <= input(2);
output(4, 133) <= input(3);
output(4, 134) <= input(4);
output(4, 135) <= input(5);
output(4, 136) <= input(6);
output(4, 137) <= input(7);
output(4, 138) <= input(8);
output(4, 139) <= input(9);
output(4, 140) <= input(10);
output(4, 141) <= input(11);
output(4, 142) <= input(12);
output(4, 143) <= input(13);
output(4, 144) <= input(38);
output(4, 145) <= input(36);
output(4, 146) <= input(0);
output(4, 147) <= input(1);
output(4, 148) <= input(2);
output(4, 149) <= input(3);
output(4, 150) <= input(4);
output(4, 151) <= input(5);
output(4, 152) <= input(6);
output(4, 153) <= input(7);
output(4, 154) <= input(8);
output(4, 155) <= input(9);
output(4, 156) <= input(10);
output(4, 157) <= input(11);
output(4, 158) <= input(12);
output(4, 159) <= input(13);
output(4, 160) <= input(38);
output(4, 161) <= input(36);
output(4, 162) <= input(0);
output(4, 163) <= input(1);
output(4, 164) <= input(2);
output(4, 165) <= input(3);
output(4, 166) <= input(4);
output(4, 167) <= input(5);
output(4, 168) <= input(6);
output(4, 169) <= input(7);
output(4, 170) <= input(8);
output(4, 171) <= input(9);
output(4, 172) <= input(10);
output(4, 173) <= input(11);
output(4, 174) <= input(12);
output(4, 175) <= input(13);
output(4, 176) <= input(38);
output(4, 177) <= input(36);
output(4, 178) <= input(0);
output(4, 179) <= input(1);
output(4, 180) <= input(2);
output(4, 181) <= input(3);
output(4, 182) <= input(4);
output(4, 183) <= input(5);
output(4, 184) <= input(6);
output(4, 185) <= input(7);
output(4, 186) <= input(8);
output(4, 187) <= input(9);
output(4, 188) <= input(10);
output(4, 189) <= input(11);
output(4, 190) <= input(12);
output(4, 191) <= input(13);
output(4, 192) <= input(38);
output(4, 193) <= input(36);
output(4, 194) <= input(0);
output(4, 195) <= input(1);
output(4, 196) <= input(2);
output(4, 197) <= input(3);
output(4, 198) <= input(4);
output(4, 199) <= input(5);
output(4, 200) <= input(6);
output(4, 201) <= input(7);
output(4, 202) <= input(8);
output(4, 203) <= input(9);
output(4, 204) <= input(10);
output(4, 205) <= input(11);
output(4, 206) <= input(12);
output(4, 207) <= input(13);
output(4, 208) <= input(38);
output(4, 209) <= input(36);
output(4, 210) <= input(0);
output(4, 211) <= input(1);
output(4, 212) <= input(2);
output(4, 213) <= input(3);
output(4, 214) <= input(4);
output(4, 215) <= input(5);
output(4, 216) <= input(6);
output(4, 217) <= input(7);
output(4, 218) <= input(8);
output(4, 219) <= input(9);
output(4, 220) <= input(10);
output(4, 221) <= input(11);
output(4, 222) <= input(12);
output(4, 223) <= input(13);
output(4, 224) <= input(38);
output(4, 225) <= input(36);
output(4, 226) <= input(0);
output(4, 227) <= input(1);
output(4, 228) <= input(2);
output(4, 229) <= input(3);
output(4, 230) <= input(4);
output(4, 231) <= input(5);
output(4, 232) <= input(6);
output(4, 233) <= input(7);
output(4, 234) <= input(8);
output(4, 235) <= input(9);
output(4, 236) <= input(10);
output(4, 237) <= input(11);
output(4, 238) <= input(12);
output(4, 239) <= input(13);
output(4, 240) <= input(38);
output(4, 241) <= input(36);
output(4, 242) <= input(0);
output(4, 243) <= input(1);
output(4, 244) <= input(2);
output(4, 245) <= input(3);
output(4, 246) <= input(4);
output(4, 247) <= input(5);
output(4, 248) <= input(6);
output(4, 249) <= input(7);
output(4, 250) <= input(8);
output(4, 251) <= input(9);
output(4, 252) <= input(10);
output(4, 253) <= input(11);
output(4, 254) <= input(12);
output(4, 255) <= input(13);
output(5, 0) <= input(39);
output(5, 1) <= input(38);
output(5, 2) <= input(36);
output(5, 3) <= input(0);
output(5, 4) <= input(1);
output(5, 5) <= input(2);
output(5, 6) <= input(3);
output(5, 7) <= input(4);
output(5, 8) <= input(5);
output(5, 9) <= input(6);
output(5, 10) <= input(7);
output(5, 11) <= input(8);
output(5, 12) <= input(9);
output(5, 13) <= input(10);
output(5, 14) <= input(11);
output(5, 15) <= input(12);
output(5, 16) <= input(39);
output(5, 17) <= input(38);
output(5, 18) <= input(36);
output(5, 19) <= input(0);
output(5, 20) <= input(1);
output(5, 21) <= input(2);
output(5, 22) <= input(3);
output(5, 23) <= input(4);
output(5, 24) <= input(5);
output(5, 25) <= input(6);
output(5, 26) <= input(7);
output(5, 27) <= input(8);
output(5, 28) <= input(9);
output(5, 29) <= input(10);
output(5, 30) <= input(11);
output(5, 31) <= input(12);
output(5, 32) <= input(39);
output(5, 33) <= input(38);
output(5, 34) <= input(36);
output(5, 35) <= input(0);
output(5, 36) <= input(1);
output(5, 37) <= input(2);
output(5, 38) <= input(3);
output(5, 39) <= input(4);
output(5, 40) <= input(5);
output(5, 41) <= input(6);
output(5, 42) <= input(7);
output(5, 43) <= input(8);
output(5, 44) <= input(9);
output(5, 45) <= input(10);
output(5, 46) <= input(11);
output(5, 47) <= input(12);
output(5, 48) <= input(39);
output(5, 49) <= input(38);
output(5, 50) <= input(36);
output(5, 51) <= input(0);
output(5, 52) <= input(1);
output(5, 53) <= input(2);
output(5, 54) <= input(3);
output(5, 55) <= input(4);
output(5, 56) <= input(5);
output(5, 57) <= input(6);
output(5, 58) <= input(7);
output(5, 59) <= input(8);
output(5, 60) <= input(9);
output(5, 61) <= input(10);
output(5, 62) <= input(11);
output(5, 63) <= input(12);
output(5, 64) <= input(39);
output(5, 65) <= input(38);
output(5, 66) <= input(36);
output(5, 67) <= input(0);
output(5, 68) <= input(1);
output(5, 69) <= input(2);
output(5, 70) <= input(3);
output(5, 71) <= input(4);
output(5, 72) <= input(5);
output(5, 73) <= input(6);
output(5, 74) <= input(7);
output(5, 75) <= input(8);
output(5, 76) <= input(9);
output(5, 77) <= input(10);
output(5, 78) <= input(11);
output(5, 79) <= input(12);
output(5, 80) <= input(39);
output(5, 81) <= input(38);
output(5, 82) <= input(36);
output(5, 83) <= input(0);
output(5, 84) <= input(1);
output(5, 85) <= input(2);
output(5, 86) <= input(3);
output(5, 87) <= input(4);
output(5, 88) <= input(5);
output(5, 89) <= input(6);
output(5, 90) <= input(7);
output(5, 91) <= input(8);
output(5, 92) <= input(9);
output(5, 93) <= input(10);
output(5, 94) <= input(11);
output(5, 95) <= input(12);
output(5, 96) <= input(39);
output(5, 97) <= input(38);
output(5, 98) <= input(36);
output(5, 99) <= input(0);
output(5, 100) <= input(1);
output(5, 101) <= input(2);
output(5, 102) <= input(3);
output(5, 103) <= input(4);
output(5, 104) <= input(5);
output(5, 105) <= input(6);
output(5, 106) <= input(7);
output(5, 107) <= input(8);
output(5, 108) <= input(9);
output(5, 109) <= input(10);
output(5, 110) <= input(11);
output(5, 111) <= input(12);
output(5, 112) <= input(39);
output(5, 113) <= input(38);
output(5, 114) <= input(36);
output(5, 115) <= input(0);
output(5, 116) <= input(1);
output(5, 117) <= input(2);
output(5, 118) <= input(3);
output(5, 119) <= input(4);
output(5, 120) <= input(5);
output(5, 121) <= input(6);
output(5, 122) <= input(7);
output(5, 123) <= input(8);
output(5, 124) <= input(9);
output(5, 125) <= input(10);
output(5, 126) <= input(11);
output(5, 127) <= input(12);
output(5, 128) <= input(39);
output(5, 129) <= input(38);
output(5, 130) <= input(36);
output(5, 131) <= input(0);
output(5, 132) <= input(1);
output(5, 133) <= input(2);
output(5, 134) <= input(3);
output(5, 135) <= input(4);
output(5, 136) <= input(5);
output(5, 137) <= input(6);
output(5, 138) <= input(7);
output(5, 139) <= input(8);
output(5, 140) <= input(9);
output(5, 141) <= input(10);
output(5, 142) <= input(11);
output(5, 143) <= input(12);
output(5, 144) <= input(39);
output(5, 145) <= input(38);
output(5, 146) <= input(36);
output(5, 147) <= input(0);
output(5, 148) <= input(1);
output(5, 149) <= input(2);
output(5, 150) <= input(3);
output(5, 151) <= input(4);
output(5, 152) <= input(5);
output(5, 153) <= input(6);
output(5, 154) <= input(7);
output(5, 155) <= input(8);
output(5, 156) <= input(9);
output(5, 157) <= input(10);
output(5, 158) <= input(11);
output(5, 159) <= input(12);
output(5, 160) <= input(39);
output(5, 161) <= input(38);
output(5, 162) <= input(36);
output(5, 163) <= input(0);
output(5, 164) <= input(1);
output(5, 165) <= input(2);
output(5, 166) <= input(3);
output(5, 167) <= input(4);
output(5, 168) <= input(5);
output(5, 169) <= input(6);
output(5, 170) <= input(7);
output(5, 171) <= input(8);
output(5, 172) <= input(9);
output(5, 173) <= input(10);
output(5, 174) <= input(11);
output(5, 175) <= input(12);
output(5, 176) <= input(39);
output(5, 177) <= input(38);
output(5, 178) <= input(36);
output(5, 179) <= input(0);
output(5, 180) <= input(1);
output(5, 181) <= input(2);
output(5, 182) <= input(3);
output(5, 183) <= input(4);
output(5, 184) <= input(5);
output(5, 185) <= input(6);
output(5, 186) <= input(7);
output(5, 187) <= input(8);
output(5, 188) <= input(9);
output(5, 189) <= input(10);
output(5, 190) <= input(11);
output(5, 191) <= input(12);
output(5, 192) <= input(39);
output(5, 193) <= input(38);
output(5, 194) <= input(36);
output(5, 195) <= input(0);
output(5, 196) <= input(1);
output(5, 197) <= input(2);
output(5, 198) <= input(3);
output(5, 199) <= input(4);
output(5, 200) <= input(5);
output(5, 201) <= input(6);
output(5, 202) <= input(7);
output(5, 203) <= input(8);
output(5, 204) <= input(9);
output(5, 205) <= input(10);
output(5, 206) <= input(11);
output(5, 207) <= input(12);
output(5, 208) <= input(39);
output(5, 209) <= input(38);
output(5, 210) <= input(36);
output(5, 211) <= input(0);
output(5, 212) <= input(1);
output(5, 213) <= input(2);
output(5, 214) <= input(3);
output(5, 215) <= input(4);
output(5, 216) <= input(5);
output(5, 217) <= input(6);
output(5, 218) <= input(7);
output(5, 219) <= input(8);
output(5, 220) <= input(9);
output(5, 221) <= input(10);
output(5, 222) <= input(11);
output(5, 223) <= input(12);
output(5, 224) <= input(39);
output(5, 225) <= input(38);
output(5, 226) <= input(36);
output(5, 227) <= input(0);
output(5, 228) <= input(1);
output(5, 229) <= input(2);
output(5, 230) <= input(3);
output(5, 231) <= input(4);
output(5, 232) <= input(5);
output(5, 233) <= input(6);
output(5, 234) <= input(7);
output(5, 235) <= input(8);
output(5, 236) <= input(9);
output(5, 237) <= input(10);
output(5, 238) <= input(11);
output(5, 239) <= input(12);
output(5, 240) <= input(39);
output(5, 241) <= input(38);
output(5, 242) <= input(36);
output(5, 243) <= input(0);
output(5, 244) <= input(1);
output(5, 245) <= input(2);
output(5, 246) <= input(3);
output(5, 247) <= input(4);
output(5, 248) <= input(5);
output(5, 249) <= input(6);
output(5, 250) <= input(7);
output(5, 251) <= input(8);
output(5, 252) <= input(9);
output(5, 253) <= input(10);
output(5, 254) <= input(11);
output(5, 255) <= input(12);
output(6, 0) <= input(40);
output(6, 1) <= input(41);
output(6, 2) <= input(37);
output(6, 3) <= input(35);
output(6, 4) <= input(16);
output(6, 5) <= input(17);
output(6, 6) <= input(18);
output(6, 7) <= input(19);
output(6, 8) <= input(20);
output(6, 9) <= input(21);
output(6, 10) <= input(22);
output(6, 11) <= input(23);
output(6, 12) <= input(24);
output(6, 13) <= input(25);
output(6, 14) <= input(26);
output(6, 15) <= input(27);
output(6, 16) <= input(40);
output(6, 17) <= input(41);
output(6, 18) <= input(37);
output(6, 19) <= input(35);
output(6, 20) <= input(16);
output(6, 21) <= input(17);
output(6, 22) <= input(18);
output(6, 23) <= input(19);
output(6, 24) <= input(20);
output(6, 25) <= input(21);
output(6, 26) <= input(22);
output(6, 27) <= input(23);
output(6, 28) <= input(24);
output(6, 29) <= input(25);
output(6, 30) <= input(26);
output(6, 31) <= input(27);
output(6, 32) <= input(40);
output(6, 33) <= input(41);
output(6, 34) <= input(37);
output(6, 35) <= input(35);
output(6, 36) <= input(16);
output(6, 37) <= input(17);
output(6, 38) <= input(18);
output(6, 39) <= input(19);
output(6, 40) <= input(20);
output(6, 41) <= input(21);
output(6, 42) <= input(22);
output(6, 43) <= input(23);
output(6, 44) <= input(24);
output(6, 45) <= input(25);
output(6, 46) <= input(26);
output(6, 47) <= input(27);
output(6, 48) <= input(40);
output(6, 49) <= input(41);
output(6, 50) <= input(37);
output(6, 51) <= input(35);
output(6, 52) <= input(16);
output(6, 53) <= input(17);
output(6, 54) <= input(18);
output(6, 55) <= input(19);
output(6, 56) <= input(20);
output(6, 57) <= input(21);
output(6, 58) <= input(22);
output(6, 59) <= input(23);
output(6, 60) <= input(24);
output(6, 61) <= input(25);
output(6, 62) <= input(26);
output(6, 63) <= input(27);
output(6, 64) <= input(40);
output(6, 65) <= input(41);
output(6, 66) <= input(37);
output(6, 67) <= input(35);
output(6, 68) <= input(16);
output(6, 69) <= input(17);
output(6, 70) <= input(18);
output(6, 71) <= input(19);
output(6, 72) <= input(20);
output(6, 73) <= input(21);
output(6, 74) <= input(22);
output(6, 75) <= input(23);
output(6, 76) <= input(24);
output(6, 77) <= input(25);
output(6, 78) <= input(26);
output(6, 79) <= input(27);
output(6, 80) <= input(40);
output(6, 81) <= input(41);
output(6, 82) <= input(37);
output(6, 83) <= input(35);
output(6, 84) <= input(16);
output(6, 85) <= input(17);
output(6, 86) <= input(18);
output(6, 87) <= input(19);
output(6, 88) <= input(20);
output(6, 89) <= input(21);
output(6, 90) <= input(22);
output(6, 91) <= input(23);
output(6, 92) <= input(24);
output(6, 93) <= input(25);
output(6, 94) <= input(26);
output(6, 95) <= input(27);
output(6, 96) <= input(40);
output(6, 97) <= input(41);
output(6, 98) <= input(37);
output(6, 99) <= input(35);
output(6, 100) <= input(16);
output(6, 101) <= input(17);
output(6, 102) <= input(18);
output(6, 103) <= input(19);
output(6, 104) <= input(20);
output(6, 105) <= input(21);
output(6, 106) <= input(22);
output(6, 107) <= input(23);
output(6, 108) <= input(24);
output(6, 109) <= input(25);
output(6, 110) <= input(26);
output(6, 111) <= input(27);
output(6, 112) <= input(40);
output(6, 113) <= input(41);
output(6, 114) <= input(37);
output(6, 115) <= input(35);
output(6, 116) <= input(16);
output(6, 117) <= input(17);
output(6, 118) <= input(18);
output(6, 119) <= input(19);
output(6, 120) <= input(20);
output(6, 121) <= input(21);
output(6, 122) <= input(22);
output(6, 123) <= input(23);
output(6, 124) <= input(24);
output(6, 125) <= input(25);
output(6, 126) <= input(26);
output(6, 127) <= input(27);
output(6, 128) <= input(42);
output(6, 129) <= input(39);
output(6, 130) <= input(38);
output(6, 131) <= input(36);
output(6, 132) <= input(0);
output(6, 133) <= input(1);
output(6, 134) <= input(2);
output(6, 135) <= input(3);
output(6, 136) <= input(4);
output(6, 137) <= input(5);
output(6, 138) <= input(6);
output(6, 139) <= input(7);
output(6, 140) <= input(8);
output(6, 141) <= input(9);
output(6, 142) <= input(10);
output(6, 143) <= input(11);
output(6, 144) <= input(42);
output(6, 145) <= input(39);
output(6, 146) <= input(38);
output(6, 147) <= input(36);
output(6, 148) <= input(0);
output(6, 149) <= input(1);
output(6, 150) <= input(2);
output(6, 151) <= input(3);
output(6, 152) <= input(4);
output(6, 153) <= input(5);
output(6, 154) <= input(6);
output(6, 155) <= input(7);
output(6, 156) <= input(8);
output(6, 157) <= input(9);
output(6, 158) <= input(10);
output(6, 159) <= input(11);
output(6, 160) <= input(42);
output(6, 161) <= input(39);
output(6, 162) <= input(38);
output(6, 163) <= input(36);
output(6, 164) <= input(0);
output(6, 165) <= input(1);
output(6, 166) <= input(2);
output(6, 167) <= input(3);
output(6, 168) <= input(4);
output(6, 169) <= input(5);
output(6, 170) <= input(6);
output(6, 171) <= input(7);
output(6, 172) <= input(8);
output(6, 173) <= input(9);
output(6, 174) <= input(10);
output(6, 175) <= input(11);
output(6, 176) <= input(42);
output(6, 177) <= input(39);
output(6, 178) <= input(38);
output(6, 179) <= input(36);
output(6, 180) <= input(0);
output(6, 181) <= input(1);
output(6, 182) <= input(2);
output(6, 183) <= input(3);
output(6, 184) <= input(4);
output(6, 185) <= input(5);
output(6, 186) <= input(6);
output(6, 187) <= input(7);
output(6, 188) <= input(8);
output(6, 189) <= input(9);
output(6, 190) <= input(10);
output(6, 191) <= input(11);
output(6, 192) <= input(42);
output(6, 193) <= input(39);
output(6, 194) <= input(38);
output(6, 195) <= input(36);
output(6, 196) <= input(0);
output(6, 197) <= input(1);
output(6, 198) <= input(2);
output(6, 199) <= input(3);
output(6, 200) <= input(4);
output(6, 201) <= input(5);
output(6, 202) <= input(6);
output(6, 203) <= input(7);
output(6, 204) <= input(8);
output(6, 205) <= input(9);
output(6, 206) <= input(10);
output(6, 207) <= input(11);
output(6, 208) <= input(42);
output(6, 209) <= input(39);
output(6, 210) <= input(38);
output(6, 211) <= input(36);
output(6, 212) <= input(0);
output(6, 213) <= input(1);
output(6, 214) <= input(2);
output(6, 215) <= input(3);
output(6, 216) <= input(4);
output(6, 217) <= input(5);
output(6, 218) <= input(6);
output(6, 219) <= input(7);
output(6, 220) <= input(8);
output(6, 221) <= input(9);
output(6, 222) <= input(10);
output(6, 223) <= input(11);
output(6, 224) <= input(42);
output(6, 225) <= input(39);
output(6, 226) <= input(38);
output(6, 227) <= input(36);
output(6, 228) <= input(0);
output(6, 229) <= input(1);
output(6, 230) <= input(2);
output(6, 231) <= input(3);
output(6, 232) <= input(4);
output(6, 233) <= input(5);
output(6, 234) <= input(6);
output(6, 235) <= input(7);
output(6, 236) <= input(8);
output(6, 237) <= input(9);
output(6, 238) <= input(10);
output(6, 239) <= input(11);
output(6, 240) <= input(42);
output(6, 241) <= input(39);
output(6, 242) <= input(38);
output(6, 243) <= input(36);
output(6, 244) <= input(0);
output(6, 245) <= input(1);
output(6, 246) <= input(2);
output(6, 247) <= input(3);
output(6, 248) <= input(4);
output(6, 249) <= input(5);
output(6, 250) <= input(6);
output(6, 251) <= input(7);
output(6, 252) <= input(8);
output(6, 253) <= input(9);
output(6, 254) <= input(10);
output(6, 255) <= input(11);
output(7, 0) <= input(42);
output(7, 1) <= input(39);
output(7, 2) <= input(38);
output(7, 3) <= input(36);
output(7, 4) <= input(0);
output(7, 5) <= input(1);
output(7, 6) <= input(2);
output(7, 7) <= input(3);
output(7, 8) <= input(4);
output(7, 9) <= input(5);
output(7, 10) <= input(6);
output(7, 11) <= input(7);
output(7, 12) <= input(8);
output(7, 13) <= input(9);
output(7, 14) <= input(10);
output(7, 15) <= input(11);
output(7, 16) <= input(42);
output(7, 17) <= input(39);
output(7, 18) <= input(38);
output(7, 19) <= input(36);
output(7, 20) <= input(0);
output(7, 21) <= input(1);
output(7, 22) <= input(2);
output(7, 23) <= input(3);
output(7, 24) <= input(4);
output(7, 25) <= input(5);
output(7, 26) <= input(6);
output(7, 27) <= input(7);
output(7, 28) <= input(8);
output(7, 29) <= input(9);
output(7, 30) <= input(10);
output(7, 31) <= input(11);
output(7, 32) <= input(42);
output(7, 33) <= input(39);
output(7, 34) <= input(38);
output(7, 35) <= input(36);
output(7, 36) <= input(0);
output(7, 37) <= input(1);
output(7, 38) <= input(2);
output(7, 39) <= input(3);
output(7, 40) <= input(4);
output(7, 41) <= input(5);
output(7, 42) <= input(6);
output(7, 43) <= input(7);
output(7, 44) <= input(8);
output(7, 45) <= input(9);
output(7, 46) <= input(10);
output(7, 47) <= input(11);
output(7, 48) <= input(42);
output(7, 49) <= input(39);
output(7, 50) <= input(38);
output(7, 51) <= input(36);
output(7, 52) <= input(0);
output(7, 53) <= input(1);
output(7, 54) <= input(2);
output(7, 55) <= input(3);
output(7, 56) <= input(4);
output(7, 57) <= input(5);
output(7, 58) <= input(6);
output(7, 59) <= input(7);
output(7, 60) <= input(8);
output(7, 61) <= input(9);
output(7, 62) <= input(10);
output(7, 63) <= input(11);
output(7, 64) <= input(42);
output(7, 65) <= input(39);
output(7, 66) <= input(38);
output(7, 67) <= input(36);
output(7, 68) <= input(0);
output(7, 69) <= input(1);
output(7, 70) <= input(2);
output(7, 71) <= input(3);
output(7, 72) <= input(4);
output(7, 73) <= input(5);
output(7, 74) <= input(6);
output(7, 75) <= input(7);
output(7, 76) <= input(8);
output(7, 77) <= input(9);
output(7, 78) <= input(10);
output(7, 79) <= input(11);
output(7, 80) <= input(43);
output(7, 81) <= input(40);
output(7, 82) <= input(41);
output(7, 83) <= input(37);
output(7, 84) <= input(35);
output(7, 85) <= input(16);
output(7, 86) <= input(17);
output(7, 87) <= input(18);
output(7, 88) <= input(19);
output(7, 89) <= input(20);
output(7, 90) <= input(21);
output(7, 91) <= input(22);
output(7, 92) <= input(23);
output(7, 93) <= input(24);
output(7, 94) <= input(25);
output(7, 95) <= input(26);
output(7, 96) <= input(43);
output(7, 97) <= input(40);
output(7, 98) <= input(41);
output(7, 99) <= input(37);
output(7, 100) <= input(35);
output(7, 101) <= input(16);
output(7, 102) <= input(17);
output(7, 103) <= input(18);
output(7, 104) <= input(19);
output(7, 105) <= input(20);
output(7, 106) <= input(21);
output(7, 107) <= input(22);
output(7, 108) <= input(23);
output(7, 109) <= input(24);
output(7, 110) <= input(25);
output(7, 111) <= input(26);
output(7, 112) <= input(43);
output(7, 113) <= input(40);
output(7, 114) <= input(41);
output(7, 115) <= input(37);
output(7, 116) <= input(35);
output(7, 117) <= input(16);
output(7, 118) <= input(17);
output(7, 119) <= input(18);
output(7, 120) <= input(19);
output(7, 121) <= input(20);
output(7, 122) <= input(21);
output(7, 123) <= input(22);
output(7, 124) <= input(23);
output(7, 125) <= input(24);
output(7, 126) <= input(25);
output(7, 127) <= input(26);
output(7, 128) <= input(43);
output(7, 129) <= input(40);
output(7, 130) <= input(41);
output(7, 131) <= input(37);
output(7, 132) <= input(35);
output(7, 133) <= input(16);
output(7, 134) <= input(17);
output(7, 135) <= input(18);
output(7, 136) <= input(19);
output(7, 137) <= input(20);
output(7, 138) <= input(21);
output(7, 139) <= input(22);
output(7, 140) <= input(23);
output(7, 141) <= input(24);
output(7, 142) <= input(25);
output(7, 143) <= input(26);
output(7, 144) <= input(43);
output(7, 145) <= input(40);
output(7, 146) <= input(41);
output(7, 147) <= input(37);
output(7, 148) <= input(35);
output(7, 149) <= input(16);
output(7, 150) <= input(17);
output(7, 151) <= input(18);
output(7, 152) <= input(19);
output(7, 153) <= input(20);
output(7, 154) <= input(21);
output(7, 155) <= input(22);
output(7, 156) <= input(23);
output(7, 157) <= input(24);
output(7, 158) <= input(25);
output(7, 159) <= input(26);
output(7, 160) <= input(44);
output(7, 161) <= input(42);
output(7, 162) <= input(39);
output(7, 163) <= input(38);
output(7, 164) <= input(36);
output(7, 165) <= input(0);
output(7, 166) <= input(1);
output(7, 167) <= input(2);
output(7, 168) <= input(3);
output(7, 169) <= input(4);
output(7, 170) <= input(5);
output(7, 171) <= input(6);
output(7, 172) <= input(7);
output(7, 173) <= input(8);
output(7, 174) <= input(9);
output(7, 175) <= input(10);
output(7, 176) <= input(44);
output(7, 177) <= input(42);
output(7, 178) <= input(39);
output(7, 179) <= input(38);
output(7, 180) <= input(36);
output(7, 181) <= input(0);
output(7, 182) <= input(1);
output(7, 183) <= input(2);
output(7, 184) <= input(3);
output(7, 185) <= input(4);
output(7, 186) <= input(5);
output(7, 187) <= input(6);
output(7, 188) <= input(7);
output(7, 189) <= input(8);
output(7, 190) <= input(9);
output(7, 191) <= input(10);
output(7, 192) <= input(44);
output(7, 193) <= input(42);
output(7, 194) <= input(39);
output(7, 195) <= input(38);
output(7, 196) <= input(36);
output(7, 197) <= input(0);
output(7, 198) <= input(1);
output(7, 199) <= input(2);
output(7, 200) <= input(3);
output(7, 201) <= input(4);
output(7, 202) <= input(5);
output(7, 203) <= input(6);
output(7, 204) <= input(7);
output(7, 205) <= input(8);
output(7, 206) <= input(9);
output(7, 207) <= input(10);
output(7, 208) <= input(44);
output(7, 209) <= input(42);
output(7, 210) <= input(39);
output(7, 211) <= input(38);
output(7, 212) <= input(36);
output(7, 213) <= input(0);
output(7, 214) <= input(1);
output(7, 215) <= input(2);
output(7, 216) <= input(3);
output(7, 217) <= input(4);
output(7, 218) <= input(5);
output(7, 219) <= input(6);
output(7, 220) <= input(7);
output(7, 221) <= input(8);
output(7, 222) <= input(9);
output(7, 223) <= input(10);
output(7, 224) <= input(44);
output(7, 225) <= input(42);
output(7, 226) <= input(39);
output(7, 227) <= input(38);
output(7, 228) <= input(36);
output(7, 229) <= input(0);
output(7, 230) <= input(1);
output(7, 231) <= input(2);
output(7, 232) <= input(3);
output(7, 233) <= input(4);
output(7, 234) <= input(5);
output(7, 235) <= input(6);
output(7, 236) <= input(7);
output(7, 237) <= input(8);
output(7, 238) <= input(9);
output(7, 239) <= input(10);
output(7, 240) <= input(44);
output(7, 241) <= input(42);
output(7, 242) <= input(39);
output(7, 243) <= input(38);
output(7, 244) <= input(36);
output(7, 245) <= input(0);
output(7, 246) <= input(1);
output(7, 247) <= input(2);
output(7, 248) <= input(3);
output(7, 249) <= input(4);
output(7, 250) <= input(5);
output(7, 251) <= input(6);
output(7, 252) <= input(7);
output(7, 253) <= input(8);
output(7, 254) <= input(9);
output(7, 255) <= input(10);
when "0011" =>
output(0, 0) <= input(0);
output(0, 1) <= input(1);
output(0, 2) <= input(2);
output(0, 3) <= input(3);
output(0, 4) <= input(4);
output(0, 5) <= input(5);
output(0, 6) <= input(6);
output(0, 7) <= input(7);
output(0, 8) <= input(8);
output(0, 9) <= input(9);
output(0, 10) <= input(10);
output(0, 11) <= input(11);
output(0, 12) <= input(12);
output(0, 13) <= input(13);
output(0, 14) <= input(14);
output(0, 15) <= input(15);
output(0, 16) <= input(0);
output(0, 17) <= input(1);
output(0, 18) <= input(2);
output(0, 19) <= input(3);
output(0, 20) <= input(4);
output(0, 21) <= input(5);
output(0, 22) <= input(6);
output(0, 23) <= input(7);
output(0, 24) <= input(8);
output(0, 25) <= input(9);
output(0, 26) <= input(10);
output(0, 27) <= input(11);
output(0, 28) <= input(12);
output(0, 29) <= input(13);
output(0, 30) <= input(14);
output(0, 31) <= input(15);
output(0, 32) <= input(0);
output(0, 33) <= input(1);
output(0, 34) <= input(2);
output(0, 35) <= input(3);
output(0, 36) <= input(4);
output(0, 37) <= input(5);
output(0, 38) <= input(6);
output(0, 39) <= input(7);
output(0, 40) <= input(8);
output(0, 41) <= input(9);
output(0, 42) <= input(10);
output(0, 43) <= input(11);
output(0, 44) <= input(12);
output(0, 45) <= input(13);
output(0, 46) <= input(14);
output(0, 47) <= input(15);
output(0, 48) <= input(0);
output(0, 49) <= input(1);
output(0, 50) <= input(2);
output(0, 51) <= input(3);
output(0, 52) <= input(4);
output(0, 53) <= input(5);
output(0, 54) <= input(6);
output(0, 55) <= input(7);
output(0, 56) <= input(8);
output(0, 57) <= input(9);
output(0, 58) <= input(10);
output(0, 59) <= input(11);
output(0, 60) <= input(12);
output(0, 61) <= input(13);
output(0, 62) <= input(14);
output(0, 63) <= input(15);
output(0, 64) <= input(16);
output(0, 65) <= input(17);
output(0, 66) <= input(18);
output(0, 67) <= input(19);
output(0, 68) <= input(20);
output(0, 69) <= input(21);
output(0, 70) <= input(22);
output(0, 71) <= input(23);
output(0, 72) <= input(24);
output(0, 73) <= input(25);
output(0, 74) <= input(26);
output(0, 75) <= input(27);
output(0, 76) <= input(28);
output(0, 77) <= input(29);
output(0, 78) <= input(30);
output(0, 79) <= input(31);
output(0, 80) <= input(16);
output(0, 81) <= input(17);
output(0, 82) <= input(18);
output(0, 83) <= input(19);
output(0, 84) <= input(20);
output(0, 85) <= input(21);
output(0, 86) <= input(22);
output(0, 87) <= input(23);
output(0, 88) <= input(24);
output(0, 89) <= input(25);
output(0, 90) <= input(26);
output(0, 91) <= input(27);
output(0, 92) <= input(28);
output(0, 93) <= input(29);
output(0, 94) <= input(30);
output(0, 95) <= input(31);
output(0, 96) <= input(16);
output(0, 97) <= input(17);
output(0, 98) <= input(18);
output(0, 99) <= input(19);
output(0, 100) <= input(20);
output(0, 101) <= input(21);
output(0, 102) <= input(22);
output(0, 103) <= input(23);
output(0, 104) <= input(24);
output(0, 105) <= input(25);
output(0, 106) <= input(26);
output(0, 107) <= input(27);
output(0, 108) <= input(28);
output(0, 109) <= input(29);
output(0, 110) <= input(30);
output(0, 111) <= input(31);
output(0, 112) <= input(16);
output(0, 113) <= input(17);
output(0, 114) <= input(18);
output(0, 115) <= input(19);
output(0, 116) <= input(20);
output(0, 117) <= input(21);
output(0, 118) <= input(22);
output(0, 119) <= input(23);
output(0, 120) <= input(24);
output(0, 121) <= input(25);
output(0, 122) <= input(26);
output(0, 123) <= input(27);
output(0, 124) <= input(28);
output(0, 125) <= input(29);
output(0, 126) <= input(30);
output(0, 127) <= input(31);
output(0, 128) <= input(32);
output(0, 129) <= input(0);
output(0, 130) <= input(1);
output(0, 131) <= input(2);
output(0, 132) <= input(3);
output(0, 133) <= input(4);
output(0, 134) <= input(5);
output(0, 135) <= input(6);
output(0, 136) <= input(7);
output(0, 137) <= input(8);
output(0, 138) <= input(9);
output(0, 139) <= input(10);
output(0, 140) <= input(11);
output(0, 141) <= input(12);
output(0, 142) <= input(13);
output(0, 143) <= input(14);
output(0, 144) <= input(32);
output(0, 145) <= input(0);
output(0, 146) <= input(1);
output(0, 147) <= input(2);
output(0, 148) <= input(3);
output(0, 149) <= input(4);
output(0, 150) <= input(5);
output(0, 151) <= input(6);
output(0, 152) <= input(7);
output(0, 153) <= input(8);
output(0, 154) <= input(9);
output(0, 155) <= input(10);
output(0, 156) <= input(11);
output(0, 157) <= input(12);
output(0, 158) <= input(13);
output(0, 159) <= input(14);
output(0, 160) <= input(32);
output(0, 161) <= input(0);
output(0, 162) <= input(1);
output(0, 163) <= input(2);
output(0, 164) <= input(3);
output(0, 165) <= input(4);
output(0, 166) <= input(5);
output(0, 167) <= input(6);
output(0, 168) <= input(7);
output(0, 169) <= input(8);
output(0, 170) <= input(9);
output(0, 171) <= input(10);
output(0, 172) <= input(11);
output(0, 173) <= input(12);
output(0, 174) <= input(13);
output(0, 175) <= input(14);
output(0, 176) <= input(32);
output(0, 177) <= input(0);
output(0, 178) <= input(1);
output(0, 179) <= input(2);
output(0, 180) <= input(3);
output(0, 181) <= input(4);
output(0, 182) <= input(5);
output(0, 183) <= input(6);
output(0, 184) <= input(7);
output(0, 185) <= input(8);
output(0, 186) <= input(9);
output(0, 187) <= input(10);
output(0, 188) <= input(11);
output(0, 189) <= input(12);
output(0, 190) <= input(13);
output(0, 191) <= input(14);
output(0, 192) <= input(33);
output(0, 193) <= input(16);
output(0, 194) <= input(17);
output(0, 195) <= input(18);
output(0, 196) <= input(19);
output(0, 197) <= input(20);
output(0, 198) <= input(21);
output(0, 199) <= input(22);
output(0, 200) <= input(23);
output(0, 201) <= input(24);
output(0, 202) <= input(25);
output(0, 203) <= input(26);
output(0, 204) <= input(27);
output(0, 205) <= input(28);
output(0, 206) <= input(29);
output(0, 207) <= input(30);
output(0, 208) <= input(33);
output(0, 209) <= input(16);
output(0, 210) <= input(17);
output(0, 211) <= input(18);
output(0, 212) <= input(19);
output(0, 213) <= input(20);
output(0, 214) <= input(21);
output(0, 215) <= input(22);
output(0, 216) <= input(23);
output(0, 217) <= input(24);
output(0, 218) <= input(25);
output(0, 219) <= input(26);
output(0, 220) <= input(27);
output(0, 221) <= input(28);
output(0, 222) <= input(29);
output(0, 223) <= input(30);
output(0, 224) <= input(33);
output(0, 225) <= input(16);
output(0, 226) <= input(17);
output(0, 227) <= input(18);
output(0, 228) <= input(19);
output(0, 229) <= input(20);
output(0, 230) <= input(21);
output(0, 231) <= input(22);
output(0, 232) <= input(23);
output(0, 233) <= input(24);
output(0, 234) <= input(25);
output(0, 235) <= input(26);
output(0, 236) <= input(27);
output(0, 237) <= input(28);
output(0, 238) <= input(29);
output(0, 239) <= input(30);
output(0, 240) <= input(33);
output(0, 241) <= input(16);
output(0, 242) <= input(17);
output(0, 243) <= input(18);
output(0, 244) <= input(19);
output(0, 245) <= input(20);
output(0, 246) <= input(21);
output(0, 247) <= input(22);
output(0, 248) <= input(23);
output(0, 249) <= input(24);
output(0, 250) <= input(25);
output(0, 251) <= input(26);
output(0, 252) <= input(27);
output(0, 253) <= input(28);
output(0, 254) <= input(29);
output(0, 255) <= input(30);
output(1, 0) <= input(32);
output(1, 1) <= input(0);
output(1, 2) <= input(1);
output(1, 3) <= input(2);
output(1, 4) <= input(3);
output(1, 5) <= input(4);
output(1, 6) <= input(5);
output(1, 7) <= input(6);
output(1, 8) <= input(7);
output(1, 9) <= input(8);
output(1, 10) <= input(9);
output(1, 11) <= input(10);
output(1, 12) <= input(11);
output(1, 13) <= input(12);
output(1, 14) <= input(13);
output(1, 15) <= input(14);
output(1, 16) <= input(32);
output(1, 17) <= input(0);
output(1, 18) <= input(1);
output(1, 19) <= input(2);
output(1, 20) <= input(3);
output(1, 21) <= input(4);
output(1, 22) <= input(5);
output(1, 23) <= input(6);
output(1, 24) <= input(7);
output(1, 25) <= input(8);
output(1, 26) <= input(9);
output(1, 27) <= input(10);
output(1, 28) <= input(11);
output(1, 29) <= input(12);
output(1, 30) <= input(13);
output(1, 31) <= input(14);
output(1, 32) <= input(33);
output(1, 33) <= input(16);
output(1, 34) <= input(17);
output(1, 35) <= input(18);
output(1, 36) <= input(19);
output(1, 37) <= input(20);
output(1, 38) <= input(21);
output(1, 39) <= input(22);
output(1, 40) <= input(23);
output(1, 41) <= input(24);
output(1, 42) <= input(25);
output(1, 43) <= input(26);
output(1, 44) <= input(27);
output(1, 45) <= input(28);
output(1, 46) <= input(29);
output(1, 47) <= input(30);
output(1, 48) <= input(33);
output(1, 49) <= input(16);
output(1, 50) <= input(17);
output(1, 51) <= input(18);
output(1, 52) <= input(19);
output(1, 53) <= input(20);
output(1, 54) <= input(21);
output(1, 55) <= input(22);
output(1, 56) <= input(23);
output(1, 57) <= input(24);
output(1, 58) <= input(25);
output(1, 59) <= input(26);
output(1, 60) <= input(27);
output(1, 61) <= input(28);
output(1, 62) <= input(29);
output(1, 63) <= input(30);
output(1, 64) <= input(33);
output(1, 65) <= input(16);
output(1, 66) <= input(17);
output(1, 67) <= input(18);
output(1, 68) <= input(19);
output(1, 69) <= input(20);
output(1, 70) <= input(21);
output(1, 71) <= input(22);
output(1, 72) <= input(23);
output(1, 73) <= input(24);
output(1, 74) <= input(25);
output(1, 75) <= input(26);
output(1, 76) <= input(27);
output(1, 77) <= input(28);
output(1, 78) <= input(29);
output(1, 79) <= input(30);
output(1, 80) <= input(34);
output(1, 81) <= input(32);
output(1, 82) <= input(0);
output(1, 83) <= input(1);
output(1, 84) <= input(2);
output(1, 85) <= input(3);
output(1, 86) <= input(4);
output(1, 87) <= input(5);
output(1, 88) <= input(6);
output(1, 89) <= input(7);
output(1, 90) <= input(8);
output(1, 91) <= input(9);
output(1, 92) <= input(10);
output(1, 93) <= input(11);
output(1, 94) <= input(12);
output(1, 95) <= input(13);
output(1, 96) <= input(34);
output(1, 97) <= input(32);
output(1, 98) <= input(0);
output(1, 99) <= input(1);
output(1, 100) <= input(2);
output(1, 101) <= input(3);
output(1, 102) <= input(4);
output(1, 103) <= input(5);
output(1, 104) <= input(6);
output(1, 105) <= input(7);
output(1, 106) <= input(8);
output(1, 107) <= input(9);
output(1, 108) <= input(10);
output(1, 109) <= input(11);
output(1, 110) <= input(12);
output(1, 111) <= input(13);
output(1, 112) <= input(34);
output(1, 113) <= input(32);
output(1, 114) <= input(0);
output(1, 115) <= input(1);
output(1, 116) <= input(2);
output(1, 117) <= input(3);
output(1, 118) <= input(4);
output(1, 119) <= input(5);
output(1, 120) <= input(6);
output(1, 121) <= input(7);
output(1, 122) <= input(8);
output(1, 123) <= input(9);
output(1, 124) <= input(10);
output(1, 125) <= input(11);
output(1, 126) <= input(12);
output(1, 127) <= input(13);
output(1, 128) <= input(35);
output(1, 129) <= input(33);
output(1, 130) <= input(16);
output(1, 131) <= input(17);
output(1, 132) <= input(18);
output(1, 133) <= input(19);
output(1, 134) <= input(20);
output(1, 135) <= input(21);
output(1, 136) <= input(22);
output(1, 137) <= input(23);
output(1, 138) <= input(24);
output(1, 139) <= input(25);
output(1, 140) <= input(26);
output(1, 141) <= input(27);
output(1, 142) <= input(28);
output(1, 143) <= input(29);
output(1, 144) <= input(35);
output(1, 145) <= input(33);
output(1, 146) <= input(16);
output(1, 147) <= input(17);
output(1, 148) <= input(18);
output(1, 149) <= input(19);
output(1, 150) <= input(20);
output(1, 151) <= input(21);
output(1, 152) <= input(22);
output(1, 153) <= input(23);
output(1, 154) <= input(24);
output(1, 155) <= input(25);
output(1, 156) <= input(26);
output(1, 157) <= input(27);
output(1, 158) <= input(28);
output(1, 159) <= input(29);
output(1, 160) <= input(36);
output(1, 161) <= input(34);
output(1, 162) <= input(32);
output(1, 163) <= input(0);
output(1, 164) <= input(1);
output(1, 165) <= input(2);
output(1, 166) <= input(3);
output(1, 167) <= input(4);
output(1, 168) <= input(5);
output(1, 169) <= input(6);
output(1, 170) <= input(7);
output(1, 171) <= input(8);
output(1, 172) <= input(9);
output(1, 173) <= input(10);
output(1, 174) <= input(11);
output(1, 175) <= input(12);
output(1, 176) <= input(36);
output(1, 177) <= input(34);
output(1, 178) <= input(32);
output(1, 179) <= input(0);
output(1, 180) <= input(1);
output(1, 181) <= input(2);
output(1, 182) <= input(3);
output(1, 183) <= input(4);
output(1, 184) <= input(5);
output(1, 185) <= input(6);
output(1, 186) <= input(7);
output(1, 187) <= input(8);
output(1, 188) <= input(9);
output(1, 189) <= input(10);
output(1, 190) <= input(11);
output(1, 191) <= input(12);
output(1, 192) <= input(36);
output(1, 193) <= input(34);
output(1, 194) <= input(32);
output(1, 195) <= input(0);
output(1, 196) <= input(1);
output(1, 197) <= input(2);
output(1, 198) <= input(3);
output(1, 199) <= input(4);
output(1, 200) <= input(5);
output(1, 201) <= input(6);
output(1, 202) <= input(7);
output(1, 203) <= input(8);
output(1, 204) <= input(9);
output(1, 205) <= input(10);
output(1, 206) <= input(11);
output(1, 207) <= input(12);
output(1, 208) <= input(37);
output(1, 209) <= input(35);
output(1, 210) <= input(33);
output(1, 211) <= input(16);
output(1, 212) <= input(17);
output(1, 213) <= input(18);
output(1, 214) <= input(19);
output(1, 215) <= input(20);
output(1, 216) <= input(21);
output(1, 217) <= input(22);
output(1, 218) <= input(23);
output(1, 219) <= input(24);
output(1, 220) <= input(25);
output(1, 221) <= input(26);
output(1, 222) <= input(27);
output(1, 223) <= input(28);
output(1, 224) <= input(37);
output(1, 225) <= input(35);
output(1, 226) <= input(33);
output(1, 227) <= input(16);
output(1, 228) <= input(17);
output(1, 229) <= input(18);
output(1, 230) <= input(19);
output(1, 231) <= input(20);
output(1, 232) <= input(21);
output(1, 233) <= input(22);
output(1, 234) <= input(23);
output(1, 235) <= input(24);
output(1, 236) <= input(25);
output(1, 237) <= input(26);
output(1, 238) <= input(27);
output(1, 239) <= input(28);
output(1, 240) <= input(37);
output(1, 241) <= input(35);
output(1, 242) <= input(33);
output(1, 243) <= input(16);
output(1, 244) <= input(17);
output(1, 245) <= input(18);
output(1, 246) <= input(19);
output(1, 247) <= input(20);
output(1, 248) <= input(21);
output(1, 249) <= input(22);
output(1, 250) <= input(23);
output(1, 251) <= input(24);
output(1, 252) <= input(25);
output(1, 253) <= input(26);
output(1, 254) <= input(27);
output(1, 255) <= input(28);
output(2, 0) <= input(34);
output(2, 1) <= input(32);
output(2, 2) <= input(0);
output(2, 3) <= input(1);
output(2, 4) <= input(2);
output(2, 5) <= input(3);
output(2, 6) <= input(4);
output(2, 7) <= input(5);
output(2, 8) <= input(6);
output(2, 9) <= input(7);
output(2, 10) <= input(8);
output(2, 11) <= input(9);
output(2, 12) <= input(10);
output(2, 13) <= input(11);
output(2, 14) <= input(12);
output(2, 15) <= input(13);
output(2, 16) <= input(34);
output(2, 17) <= input(32);
output(2, 18) <= input(0);
output(2, 19) <= input(1);
output(2, 20) <= input(2);
output(2, 21) <= input(3);
output(2, 22) <= input(4);
output(2, 23) <= input(5);
output(2, 24) <= input(6);
output(2, 25) <= input(7);
output(2, 26) <= input(8);
output(2, 27) <= input(9);
output(2, 28) <= input(10);
output(2, 29) <= input(11);
output(2, 30) <= input(12);
output(2, 31) <= input(13);
output(2, 32) <= input(35);
output(2, 33) <= input(33);
output(2, 34) <= input(16);
output(2, 35) <= input(17);
output(2, 36) <= input(18);
output(2, 37) <= input(19);
output(2, 38) <= input(20);
output(2, 39) <= input(21);
output(2, 40) <= input(22);
output(2, 41) <= input(23);
output(2, 42) <= input(24);
output(2, 43) <= input(25);
output(2, 44) <= input(26);
output(2, 45) <= input(27);
output(2, 46) <= input(28);
output(2, 47) <= input(29);
output(2, 48) <= input(35);
output(2, 49) <= input(33);
output(2, 50) <= input(16);
output(2, 51) <= input(17);
output(2, 52) <= input(18);
output(2, 53) <= input(19);
output(2, 54) <= input(20);
output(2, 55) <= input(21);
output(2, 56) <= input(22);
output(2, 57) <= input(23);
output(2, 58) <= input(24);
output(2, 59) <= input(25);
output(2, 60) <= input(26);
output(2, 61) <= input(27);
output(2, 62) <= input(28);
output(2, 63) <= input(29);
output(2, 64) <= input(36);
output(2, 65) <= input(34);
output(2, 66) <= input(32);
output(2, 67) <= input(0);
output(2, 68) <= input(1);
output(2, 69) <= input(2);
output(2, 70) <= input(3);
output(2, 71) <= input(4);
output(2, 72) <= input(5);
output(2, 73) <= input(6);
output(2, 74) <= input(7);
output(2, 75) <= input(8);
output(2, 76) <= input(9);
output(2, 77) <= input(10);
output(2, 78) <= input(11);
output(2, 79) <= input(12);
output(2, 80) <= input(36);
output(2, 81) <= input(34);
output(2, 82) <= input(32);
output(2, 83) <= input(0);
output(2, 84) <= input(1);
output(2, 85) <= input(2);
output(2, 86) <= input(3);
output(2, 87) <= input(4);
output(2, 88) <= input(5);
output(2, 89) <= input(6);
output(2, 90) <= input(7);
output(2, 91) <= input(8);
output(2, 92) <= input(9);
output(2, 93) <= input(10);
output(2, 94) <= input(11);
output(2, 95) <= input(12);
output(2, 96) <= input(37);
output(2, 97) <= input(35);
output(2, 98) <= input(33);
output(2, 99) <= input(16);
output(2, 100) <= input(17);
output(2, 101) <= input(18);
output(2, 102) <= input(19);
output(2, 103) <= input(20);
output(2, 104) <= input(21);
output(2, 105) <= input(22);
output(2, 106) <= input(23);
output(2, 107) <= input(24);
output(2, 108) <= input(25);
output(2, 109) <= input(26);
output(2, 110) <= input(27);
output(2, 111) <= input(28);
output(2, 112) <= input(37);
output(2, 113) <= input(35);
output(2, 114) <= input(33);
output(2, 115) <= input(16);
output(2, 116) <= input(17);
output(2, 117) <= input(18);
output(2, 118) <= input(19);
output(2, 119) <= input(20);
output(2, 120) <= input(21);
output(2, 121) <= input(22);
output(2, 122) <= input(23);
output(2, 123) <= input(24);
output(2, 124) <= input(25);
output(2, 125) <= input(26);
output(2, 126) <= input(27);
output(2, 127) <= input(28);
output(2, 128) <= input(38);
output(2, 129) <= input(36);
output(2, 130) <= input(34);
output(2, 131) <= input(32);
output(2, 132) <= input(0);
output(2, 133) <= input(1);
output(2, 134) <= input(2);
output(2, 135) <= input(3);
output(2, 136) <= input(4);
output(2, 137) <= input(5);
output(2, 138) <= input(6);
output(2, 139) <= input(7);
output(2, 140) <= input(8);
output(2, 141) <= input(9);
output(2, 142) <= input(10);
output(2, 143) <= input(11);
output(2, 144) <= input(38);
output(2, 145) <= input(36);
output(2, 146) <= input(34);
output(2, 147) <= input(32);
output(2, 148) <= input(0);
output(2, 149) <= input(1);
output(2, 150) <= input(2);
output(2, 151) <= input(3);
output(2, 152) <= input(4);
output(2, 153) <= input(5);
output(2, 154) <= input(6);
output(2, 155) <= input(7);
output(2, 156) <= input(8);
output(2, 157) <= input(9);
output(2, 158) <= input(10);
output(2, 159) <= input(11);
output(2, 160) <= input(39);
output(2, 161) <= input(37);
output(2, 162) <= input(35);
output(2, 163) <= input(33);
output(2, 164) <= input(16);
output(2, 165) <= input(17);
output(2, 166) <= input(18);
output(2, 167) <= input(19);
output(2, 168) <= input(20);
output(2, 169) <= input(21);
output(2, 170) <= input(22);
output(2, 171) <= input(23);
output(2, 172) <= input(24);
output(2, 173) <= input(25);
output(2, 174) <= input(26);
output(2, 175) <= input(27);
output(2, 176) <= input(39);
output(2, 177) <= input(37);
output(2, 178) <= input(35);
output(2, 179) <= input(33);
output(2, 180) <= input(16);
output(2, 181) <= input(17);
output(2, 182) <= input(18);
output(2, 183) <= input(19);
output(2, 184) <= input(20);
output(2, 185) <= input(21);
output(2, 186) <= input(22);
output(2, 187) <= input(23);
output(2, 188) <= input(24);
output(2, 189) <= input(25);
output(2, 190) <= input(26);
output(2, 191) <= input(27);
output(2, 192) <= input(40);
output(2, 193) <= input(38);
output(2, 194) <= input(36);
output(2, 195) <= input(34);
output(2, 196) <= input(32);
output(2, 197) <= input(0);
output(2, 198) <= input(1);
output(2, 199) <= input(2);
output(2, 200) <= input(3);
output(2, 201) <= input(4);
output(2, 202) <= input(5);
output(2, 203) <= input(6);
output(2, 204) <= input(7);
output(2, 205) <= input(8);
output(2, 206) <= input(9);
output(2, 207) <= input(10);
output(2, 208) <= input(40);
output(2, 209) <= input(38);
output(2, 210) <= input(36);
output(2, 211) <= input(34);
output(2, 212) <= input(32);
output(2, 213) <= input(0);
output(2, 214) <= input(1);
output(2, 215) <= input(2);
output(2, 216) <= input(3);
output(2, 217) <= input(4);
output(2, 218) <= input(5);
output(2, 219) <= input(6);
output(2, 220) <= input(7);
output(2, 221) <= input(8);
output(2, 222) <= input(9);
output(2, 223) <= input(10);
output(2, 224) <= input(41);
output(2, 225) <= input(39);
output(2, 226) <= input(37);
output(2, 227) <= input(35);
output(2, 228) <= input(33);
output(2, 229) <= input(16);
output(2, 230) <= input(17);
output(2, 231) <= input(18);
output(2, 232) <= input(19);
output(2, 233) <= input(20);
output(2, 234) <= input(21);
output(2, 235) <= input(22);
output(2, 236) <= input(23);
output(2, 237) <= input(24);
output(2, 238) <= input(25);
output(2, 239) <= input(26);
output(2, 240) <= input(41);
output(2, 241) <= input(39);
output(2, 242) <= input(37);
output(2, 243) <= input(35);
output(2, 244) <= input(33);
output(2, 245) <= input(16);
output(2, 246) <= input(17);
output(2, 247) <= input(18);
output(2, 248) <= input(19);
output(2, 249) <= input(20);
output(2, 250) <= input(21);
output(2, 251) <= input(22);
output(2, 252) <= input(23);
output(2, 253) <= input(24);
output(2, 254) <= input(25);
output(2, 255) <= input(26);
when "0100" =>
output(0, 0) <= input(0);
output(0, 1) <= input(1);
output(0, 2) <= input(2);
output(0, 3) <= input(3);
output(0, 4) <= input(4);
output(0, 5) <= input(5);
output(0, 6) <= input(6);
output(0, 7) <= input(7);
output(0, 8) <= input(8);
output(0, 9) <= input(9);
output(0, 10) <= input(10);
output(0, 11) <= input(11);
output(0, 12) <= input(12);
output(0, 13) <= input(13);
output(0, 14) <= input(14);
output(0, 15) <= input(15);
output(0, 16) <= input(16);
output(0, 17) <= input(17);
output(0, 18) <= input(18);
output(0, 19) <= input(19);
output(0, 20) <= input(20);
output(0, 21) <= input(21);
output(0, 22) <= input(22);
output(0, 23) <= input(23);
output(0, 24) <= input(24);
output(0, 25) <= input(25);
output(0, 26) <= input(26);
output(0, 27) <= input(27);
output(0, 28) <= input(28);
output(0, 29) <= input(29);
output(0, 30) <= input(30);
output(0, 31) <= input(31);
output(0, 32) <= input(16);
output(0, 33) <= input(17);
output(0, 34) <= input(18);
output(0, 35) <= input(19);
output(0, 36) <= input(20);
output(0, 37) <= input(21);
output(0, 38) <= input(22);
output(0, 39) <= input(23);
output(0, 40) <= input(24);
output(0, 41) <= input(25);
output(0, 42) <= input(26);
output(0, 43) <= input(27);
output(0, 44) <= input(28);
output(0, 45) <= input(29);
output(0, 46) <= input(30);
output(0, 47) <= input(31);
output(0, 48) <= input(32);
output(0, 49) <= input(0);
output(0, 50) <= input(1);
output(0, 51) <= input(2);
output(0, 52) <= input(3);
output(0, 53) <= input(4);
output(0, 54) <= input(5);
output(0, 55) <= input(6);
output(0, 56) <= input(7);
output(0, 57) <= input(8);
output(0, 58) <= input(9);
output(0, 59) <= input(10);
output(0, 60) <= input(11);
output(0, 61) <= input(12);
output(0, 62) <= input(13);
output(0, 63) <= input(14);
output(0, 64) <= input(33);
output(0, 65) <= input(16);
output(0, 66) <= input(17);
output(0, 67) <= input(18);
output(0, 68) <= input(19);
output(0, 69) <= input(20);
output(0, 70) <= input(21);
output(0, 71) <= input(22);
output(0, 72) <= input(23);
output(0, 73) <= input(24);
output(0, 74) <= input(25);
output(0, 75) <= input(26);
output(0, 76) <= input(27);
output(0, 77) <= input(28);
output(0, 78) <= input(29);
output(0, 79) <= input(30);
output(0, 80) <= input(33);
output(0, 81) <= input(16);
output(0, 82) <= input(17);
output(0, 83) <= input(18);
output(0, 84) <= input(19);
output(0, 85) <= input(20);
output(0, 86) <= input(21);
output(0, 87) <= input(22);
output(0, 88) <= input(23);
output(0, 89) <= input(24);
output(0, 90) <= input(25);
output(0, 91) <= input(26);
output(0, 92) <= input(27);
output(0, 93) <= input(28);
output(0, 94) <= input(29);
output(0, 95) <= input(30);
output(0, 96) <= input(34);
output(0, 97) <= input(32);
output(0, 98) <= input(0);
output(0, 99) <= input(1);
output(0, 100) <= input(2);
output(0, 101) <= input(3);
output(0, 102) <= input(4);
output(0, 103) <= input(5);
output(0, 104) <= input(6);
output(0, 105) <= input(7);
output(0, 106) <= input(8);
output(0, 107) <= input(9);
output(0, 108) <= input(10);
output(0, 109) <= input(11);
output(0, 110) <= input(12);
output(0, 111) <= input(13);
output(0, 112) <= input(34);
output(0, 113) <= input(32);
output(0, 114) <= input(0);
output(0, 115) <= input(1);
output(0, 116) <= input(2);
output(0, 117) <= input(3);
output(0, 118) <= input(4);
output(0, 119) <= input(5);
output(0, 120) <= input(6);
output(0, 121) <= input(7);
output(0, 122) <= input(8);
output(0, 123) <= input(9);
output(0, 124) <= input(10);
output(0, 125) <= input(11);
output(0, 126) <= input(12);
output(0, 127) <= input(13);
output(0, 128) <= input(35);
output(0, 129) <= input(33);
output(0, 130) <= input(16);
output(0, 131) <= input(17);
output(0, 132) <= input(18);
output(0, 133) <= input(19);
output(0, 134) <= input(20);
output(0, 135) <= input(21);
output(0, 136) <= input(22);
output(0, 137) <= input(23);
output(0, 138) <= input(24);
output(0, 139) <= input(25);
output(0, 140) <= input(26);
output(0, 141) <= input(27);
output(0, 142) <= input(28);
output(0, 143) <= input(29);
output(0, 144) <= input(36);
output(0, 145) <= input(34);
output(0, 146) <= input(32);
output(0, 147) <= input(0);
output(0, 148) <= input(1);
output(0, 149) <= input(2);
output(0, 150) <= input(3);
output(0, 151) <= input(4);
output(0, 152) <= input(5);
output(0, 153) <= input(6);
output(0, 154) <= input(7);
output(0, 155) <= input(8);
output(0, 156) <= input(9);
output(0, 157) <= input(10);
output(0, 158) <= input(11);
output(0, 159) <= input(12);
output(0, 160) <= input(36);
output(0, 161) <= input(34);
output(0, 162) <= input(32);
output(0, 163) <= input(0);
output(0, 164) <= input(1);
output(0, 165) <= input(2);
output(0, 166) <= input(3);
output(0, 167) <= input(4);
output(0, 168) <= input(5);
output(0, 169) <= input(6);
output(0, 170) <= input(7);
output(0, 171) <= input(8);
output(0, 172) <= input(9);
output(0, 173) <= input(10);
output(0, 174) <= input(11);
output(0, 175) <= input(12);
output(0, 176) <= input(37);
output(0, 177) <= input(35);
output(0, 178) <= input(33);
output(0, 179) <= input(16);
output(0, 180) <= input(17);
output(0, 181) <= input(18);
output(0, 182) <= input(19);
output(0, 183) <= input(20);
output(0, 184) <= input(21);
output(0, 185) <= input(22);
output(0, 186) <= input(23);
output(0, 187) <= input(24);
output(0, 188) <= input(25);
output(0, 189) <= input(26);
output(0, 190) <= input(27);
output(0, 191) <= input(28);
output(0, 192) <= input(38);
output(0, 193) <= input(36);
output(0, 194) <= input(34);
output(0, 195) <= input(32);
output(0, 196) <= input(0);
output(0, 197) <= input(1);
output(0, 198) <= input(2);
output(0, 199) <= input(3);
output(0, 200) <= input(4);
output(0, 201) <= input(5);
output(0, 202) <= input(6);
output(0, 203) <= input(7);
output(0, 204) <= input(8);
output(0, 205) <= input(9);
output(0, 206) <= input(10);
output(0, 207) <= input(11);
output(0, 208) <= input(38);
output(0, 209) <= input(36);
output(0, 210) <= input(34);
output(0, 211) <= input(32);
output(0, 212) <= input(0);
output(0, 213) <= input(1);
output(0, 214) <= input(2);
output(0, 215) <= input(3);
output(0, 216) <= input(4);
output(0, 217) <= input(5);
output(0, 218) <= input(6);
output(0, 219) <= input(7);
output(0, 220) <= input(8);
output(0, 221) <= input(9);
output(0, 222) <= input(10);
output(0, 223) <= input(11);
output(0, 224) <= input(39);
output(0, 225) <= input(37);
output(0, 226) <= input(35);
output(0, 227) <= input(33);
output(0, 228) <= input(16);
output(0, 229) <= input(17);
output(0, 230) <= input(18);
output(0, 231) <= input(19);
output(0, 232) <= input(20);
output(0, 233) <= input(21);
output(0, 234) <= input(22);
output(0, 235) <= input(23);
output(0, 236) <= input(24);
output(0, 237) <= input(25);
output(0, 238) <= input(26);
output(0, 239) <= input(27);
output(0, 240) <= input(39);
output(0, 241) <= input(37);
output(0, 242) <= input(35);
output(0, 243) <= input(33);
output(0, 244) <= input(16);
output(0, 245) <= input(17);
output(0, 246) <= input(18);
output(0, 247) <= input(19);
output(0, 248) <= input(20);
output(0, 249) <= input(21);
output(0, 250) <= input(22);
output(0, 251) <= input(23);
output(0, 252) <= input(24);
output(0, 253) <= input(25);
output(0, 254) <= input(26);
output(0, 255) <= input(27);
output(1, 0) <= input(32);
output(1, 1) <= input(0);
output(1, 2) <= input(1);
output(1, 3) <= input(2);
output(1, 4) <= input(3);
output(1, 5) <= input(4);
output(1, 6) <= input(5);
output(1, 7) <= input(6);
output(1, 8) <= input(7);
output(1, 9) <= input(8);
output(1, 10) <= input(9);
output(1, 11) <= input(10);
output(1, 12) <= input(11);
output(1, 13) <= input(12);
output(1, 14) <= input(13);
output(1, 15) <= input(14);
output(1, 16) <= input(33);
output(1, 17) <= input(16);
output(1, 18) <= input(17);
output(1, 19) <= input(18);
output(1, 20) <= input(19);
output(1, 21) <= input(20);
output(1, 22) <= input(21);
output(1, 23) <= input(22);
output(1, 24) <= input(23);
output(1, 25) <= input(24);
output(1, 26) <= input(25);
output(1, 27) <= input(26);
output(1, 28) <= input(27);
output(1, 29) <= input(28);
output(1, 30) <= input(29);
output(1, 31) <= input(30);
output(1, 32) <= input(34);
output(1, 33) <= input(32);
output(1, 34) <= input(0);
output(1, 35) <= input(1);
output(1, 36) <= input(2);
output(1, 37) <= input(3);
output(1, 38) <= input(4);
output(1, 39) <= input(5);
output(1, 40) <= input(6);
output(1, 41) <= input(7);
output(1, 42) <= input(8);
output(1, 43) <= input(9);
output(1, 44) <= input(10);
output(1, 45) <= input(11);
output(1, 46) <= input(12);
output(1, 47) <= input(13);
output(1, 48) <= input(34);
output(1, 49) <= input(32);
output(1, 50) <= input(0);
output(1, 51) <= input(1);
output(1, 52) <= input(2);
output(1, 53) <= input(3);
output(1, 54) <= input(4);
output(1, 55) <= input(5);
output(1, 56) <= input(6);
output(1, 57) <= input(7);
output(1, 58) <= input(8);
output(1, 59) <= input(9);
output(1, 60) <= input(10);
output(1, 61) <= input(11);
output(1, 62) <= input(12);
output(1, 63) <= input(13);
output(1, 64) <= input(35);
output(1, 65) <= input(33);
output(1, 66) <= input(16);
output(1, 67) <= input(17);
output(1, 68) <= input(18);
output(1, 69) <= input(19);
output(1, 70) <= input(20);
output(1, 71) <= input(21);
output(1, 72) <= input(22);
output(1, 73) <= input(23);
output(1, 74) <= input(24);
output(1, 75) <= input(25);
output(1, 76) <= input(26);
output(1, 77) <= input(27);
output(1, 78) <= input(28);
output(1, 79) <= input(29);
output(1, 80) <= input(36);
output(1, 81) <= input(34);
output(1, 82) <= input(32);
output(1, 83) <= input(0);
output(1, 84) <= input(1);
output(1, 85) <= input(2);
output(1, 86) <= input(3);
output(1, 87) <= input(4);
output(1, 88) <= input(5);
output(1, 89) <= input(6);
output(1, 90) <= input(7);
output(1, 91) <= input(8);
output(1, 92) <= input(9);
output(1, 93) <= input(10);
output(1, 94) <= input(11);
output(1, 95) <= input(12);
output(1, 96) <= input(37);
output(1, 97) <= input(35);
output(1, 98) <= input(33);
output(1, 99) <= input(16);
output(1, 100) <= input(17);
output(1, 101) <= input(18);
output(1, 102) <= input(19);
output(1, 103) <= input(20);
output(1, 104) <= input(21);
output(1, 105) <= input(22);
output(1, 106) <= input(23);
output(1, 107) <= input(24);
output(1, 108) <= input(25);
output(1, 109) <= input(26);
output(1, 110) <= input(27);
output(1, 111) <= input(28);
output(1, 112) <= input(37);
output(1, 113) <= input(35);
output(1, 114) <= input(33);
output(1, 115) <= input(16);
output(1, 116) <= input(17);
output(1, 117) <= input(18);
output(1, 118) <= input(19);
output(1, 119) <= input(20);
output(1, 120) <= input(21);
output(1, 121) <= input(22);
output(1, 122) <= input(23);
output(1, 123) <= input(24);
output(1, 124) <= input(25);
output(1, 125) <= input(26);
output(1, 126) <= input(27);
output(1, 127) <= input(28);
output(1, 128) <= input(38);
output(1, 129) <= input(36);
output(1, 130) <= input(34);
output(1, 131) <= input(32);
output(1, 132) <= input(0);
output(1, 133) <= input(1);
output(1, 134) <= input(2);
output(1, 135) <= input(3);
output(1, 136) <= input(4);
output(1, 137) <= input(5);
output(1, 138) <= input(6);
output(1, 139) <= input(7);
output(1, 140) <= input(8);
output(1, 141) <= input(9);
output(1, 142) <= input(10);
output(1, 143) <= input(11);
output(1, 144) <= input(39);
output(1, 145) <= input(37);
output(1, 146) <= input(35);
output(1, 147) <= input(33);
output(1, 148) <= input(16);
output(1, 149) <= input(17);
output(1, 150) <= input(18);
output(1, 151) <= input(19);
output(1, 152) <= input(20);
output(1, 153) <= input(21);
output(1, 154) <= input(22);
output(1, 155) <= input(23);
output(1, 156) <= input(24);
output(1, 157) <= input(25);
output(1, 158) <= input(26);
output(1, 159) <= input(27);
output(1, 160) <= input(40);
output(1, 161) <= input(38);
output(1, 162) <= input(36);
output(1, 163) <= input(34);
output(1, 164) <= input(32);
output(1, 165) <= input(0);
output(1, 166) <= input(1);
output(1, 167) <= input(2);
output(1, 168) <= input(3);
output(1, 169) <= input(4);
output(1, 170) <= input(5);
output(1, 171) <= input(6);
output(1, 172) <= input(7);
output(1, 173) <= input(8);
output(1, 174) <= input(9);
output(1, 175) <= input(10);
output(1, 176) <= input(40);
output(1, 177) <= input(38);
output(1, 178) <= input(36);
output(1, 179) <= input(34);
output(1, 180) <= input(32);
output(1, 181) <= input(0);
output(1, 182) <= input(1);
output(1, 183) <= input(2);
output(1, 184) <= input(3);
output(1, 185) <= input(4);
output(1, 186) <= input(5);
output(1, 187) <= input(6);
output(1, 188) <= input(7);
output(1, 189) <= input(8);
output(1, 190) <= input(9);
output(1, 191) <= input(10);
output(1, 192) <= input(41);
output(1, 193) <= input(39);
output(1, 194) <= input(37);
output(1, 195) <= input(35);
output(1, 196) <= input(33);
output(1, 197) <= input(16);
output(1, 198) <= input(17);
output(1, 199) <= input(18);
output(1, 200) <= input(19);
output(1, 201) <= input(20);
output(1, 202) <= input(21);
output(1, 203) <= input(22);
output(1, 204) <= input(23);
output(1, 205) <= input(24);
output(1, 206) <= input(25);
output(1, 207) <= input(26);
output(1, 208) <= input(42);
output(1, 209) <= input(40);
output(1, 210) <= input(38);
output(1, 211) <= input(36);
output(1, 212) <= input(34);
output(1, 213) <= input(32);
output(1, 214) <= input(0);
output(1, 215) <= input(1);
output(1, 216) <= input(2);
output(1, 217) <= input(3);
output(1, 218) <= input(4);
output(1, 219) <= input(5);
output(1, 220) <= input(6);
output(1, 221) <= input(7);
output(1, 222) <= input(8);
output(1, 223) <= input(9);
output(1, 224) <= input(43);
output(1, 225) <= input(41);
output(1, 226) <= input(39);
output(1, 227) <= input(37);
output(1, 228) <= input(35);
output(1, 229) <= input(33);
output(1, 230) <= input(16);
output(1, 231) <= input(17);
output(1, 232) <= input(18);
output(1, 233) <= input(19);
output(1, 234) <= input(20);
output(1, 235) <= input(21);
output(1, 236) <= input(22);
output(1, 237) <= input(23);
output(1, 238) <= input(24);
output(1, 239) <= input(25);
output(1, 240) <= input(43);
output(1, 241) <= input(41);
output(1, 242) <= input(39);
output(1, 243) <= input(37);
output(1, 244) <= input(35);
output(1, 245) <= input(33);
output(1, 246) <= input(16);
output(1, 247) <= input(17);
output(1, 248) <= input(18);
output(1, 249) <= input(19);
output(1, 250) <= input(20);
output(1, 251) <= input(21);
output(1, 252) <= input(22);
output(1, 253) <= input(23);
output(1, 254) <= input(24);
output(1, 255) <= input(25);
output(2, 0) <= input(34);
output(2, 1) <= input(32);
output(2, 2) <= input(0);
output(2, 3) <= input(1);
output(2, 4) <= input(2);
output(2, 5) <= input(3);
output(2, 6) <= input(4);
output(2, 7) <= input(5);
output(2, 8) <= input(6);
output(2, 9) <= input(7);
output(2, 10) <= input(8);
output(2, 11) <= input(9);
output(2, 12) <= input(10);
output(2, 13) <= input(11);
output(2, 14) <= input(12);
output(2, 15) <= input(13);
output(2, 16) <= input(35);
output(2, 17) <= input(33);
output(2, 18) <= input(16);
output(2, 19) <= input(17);
output(2, 20) <= input(18);
output(2, 21) <= input(19);
output(2, 22) <= input(20);
output(2, 23) <= input(21);
output(2, 24) <= input(22);
output(2, 25) <= input(23);
output(2, 26) <= input(24);
output(2, 27) <= input(25);
output(2, 28) <= input(26);
output(2, 29) <= input(27);
output(2, 30) <= input(28);
output(2, 31) <= input(29);
output(2, 32) <= input(36);
output(2, 33) <= input(34);
output(2, 34) <= input(32);
output(2, 35) <= input(0);
output(2, 36) <= input(1);
output(2, 37) <= input(2);
output(2, 38) <= input(3);
output(2, 39) <= input(4);
output(2, 40) <= input(5);
output(2, 41) <= input(6);
output(2, 42) <= input(7);
output(2, 43) <= input(8);
output(2, 44) <= input(9);
output(2, 45) <= input(10);
output(2, 46) <= input(11);
output(2, 47) <= input(12);
output(2, 48) <= input(37);
output(2, 49) <= input(35);
output(2, 50) <= input(33);
output(2, 51) <= input(16);
output(2, 52) <= input(17);
output(2, 53) <= input(18);
output(2, 54) <= input(19);
output(2, 55) <= input(20);
output(2, 56) <= input(21);
output(2, 57) <= input(22);
output(2, 58) <= input(23);
output(2, 59) <= input(24);
output(2, 60) <= input(25);
output(2, 61) <= input(26);
output(2, 62) <= input(27);
output(2, 63) <= input(28);
output(2, 64) <= input(38);
output(2, 65) <= input(36);
output(2, 66) <= input(34);
output(2, 67) <= input(32);
output(2, 68) <= input(0);
output(2, 69) <= input(1);
output(2, 70) <= input(2);
output(2, 71) <= input(3);
output(2, 72) <= input(4);
output(2, 73) <= input(5);
output(2, 74) <= input(6);
output(2, 75) <= input(7);
output(2, 76) <= input(8);
output(2, 77) <= input(9);
output(2, 78) <= input(10);
output(2, 79) <= input(11);
output(2, 80) <= input(39);
output(2, 81) <= input(37);
output(2, 82) <= input(35);
output(2, 83) <= input(33);
output(2, 84) <= input(16);
output(2, 85) <= input(17);
output(2, 86) <= input(18);
output(2, 87) <= input(19);
output(2, 88) <= input(20);
output(2, 89) <= input(21);
output(2, 90) <= input(22);
output(2, 91) <= input(23);
output(2, 92) <= input(24);
output(2, 93) <= input(25);
output(2, 94) <= input(26);
output(2, 95) <= input(27);
output(2, 96) <= input(40);
output(2, 97) <= input(38);
output(2, 98) <= input(36);
output(2, 99) <= input(34);
output(2, 100) <= input(32);
output(2, 101) <= input(0);
output(2, 102) <= input(1);
output(2, 103) <= input(2);
output(2, 104) <= input(3);
output(2, 105) <= input(4);
output(2, 106) <= input(5);
output(2, 107) <= input(6);
output(2, 108) <= input(7);
output(2, 109) <= input(8);
output(2, 110) <= input(9);
output(2, 111) <= input(10);
output(2, 112) <= input(40);
output(2, 113) <= input(38);
output(2, 114) <= input(36);
output(2, 115) <= input(34);
output(2, 116) <= input(32);
output(2, 117) <= input(0);
output(2, 118) <= input(1);
output(2, 119) <= input(2);
output(2, 120) <= input(3);
output(2, 121) <= input(4);
output(2, 122) <= input(5);
output(2, 123) <= input(6);
output(2, 124) <= input(7);
output(2, 125) <= input(8);
output(2, 126) <= input(9);
output(2, 127) <= input(10);
output(2, 128) <= input(41);
output(2, 129) <= input(39);
output(2, 130) <= input(37);
output(2, 131) <= input(35);
output(2, 132) <= input(33);
output(2, 133) <= input(16);
output(2, 134) <= input(17);
output(2, 135) <= input(18);
output(2, 136) <= input(19);
output(2, 137) <= input(20);
output(2, 138) <= input(21);
output(2, 139) <= input(22);
output(2, 140) <= input(23);
output(2, 141) <= input(24);
output(2, 142) <= input(25);
output(2, 143) <= input(26);
output(2, 144) <= input(42);
output(2, 145) <= input(40);
output(2, 146) <= input(38);
output(2, 147) <= input(36);
output(2, 148) <= input(34);
output(2, 149) <= input(32);
output(2, 150) <= input(0);
output(2, 151) <= input(1);
output(2, 152) <= input(2);
output(2, 153) <= input(3);
output(2, 154) <= input(4);
output(2, 155) <= input(5);
output(2, 156) <= input(6);
output(2, 157) <= input(7);
output(2, 158) <= input(8);
output(2, 159) <= input(9);
output(2, 160) <= input(43);
output(2, 161) <= input(41);
output(2, 162) <= input(39);
output(2, 163) <= input(37);
output(2, 164) <= input(35);
output(2, 165) <= input(33);
output(2, 166) <= input(16);
output(2, 167) <= input(17);
output(2, 168) <= input(18);
output(2, 169) <= input(19);
output(2, 170) <= input(20);
output(2, 171) <= input(21);
output(2, 172) <= input(22);
output(2, 173) <= input(23);
output(2, 174) <= input(24);
output(2, 175) <= input(25);
output(2, 176) <= input(44);
output(2, 177) <= input(42);
output(2, 178) <= input(40);
output(2, 179) <= input(38);
output(2, 180) <= input(36);
output(2, 181) <= input(34);
output(2, 182) <= input(32);
output(2, 183) <= input(0);
output(2, 184) <= input(1);
output(2, 185) <= input(2);
output(2, 186) <= input(3);
output(2, 187) <= input(4);
output(2, 188) <= input(5);
output(2, 189) <= input(6);
output(2, 190) <= input(7);
output(2, 191) <= input(8);
output(2, 192) <= input(45);
output(2, 193) <= input(43);
output(2, 194) <= input(41);
output(2, 195) <= input(39);
output(2, 196) <= input(37);
output(2, 197) <= input(35);
output(2, 198) <= input(33);
output(2, 199) <= input(16);
output(2, 200) <= input(17);
output(2, 201) <= input(18);
output(2, 202) <= input(19);
output(2, 203) <= input(20);
output(2, 204) <= input(21);
output(2, 205) <= input(22);
output(2, 206) <= input(23);
output(2, 207) <= input(24);
output(2, 208) <= input(46);
output(2, 209) <= input(44);
output(2, 210) <= input(42);
output(2, 211) <= input(40);
output(2, 212) <= input(38);
output(2, 213) <= input(36);
output(2, 214) <= input(34);
output(2, 215) <= input(32);
output(2, 216) <= input(0);
output(2, 217) <= input(1);
output(2, 218) <= input(2);
output(2, 219) <= input(3);
output(2, 220) <= input(4);
output(2, 221) <= input(5);
output(2, 222) <= input(6);
output(2, 223) <= input(7);
output(2, 224) <= input(47);
output(2, 225) <= input(45);
output(2, 226) <= input(43);
output(2, 227) <= input(41);
output(2, 228) <= input(39);
output(2, 229) <= input(37);
output(2, 230) <= input(35);
output(2, 231) <= input(33);
output(2, 232) <= input(16);
output(2, 233) <= input(17);
output(2, 234) <= input(18);
output(2, 235) <= input(19);
output(2, 236) <= input(20);
output(2, 237) <= input(21);
output(2, 238) <= input(22);
output(2, 239) <= input(23);
output(2, 240) <= input(47);
output(2, 241) <= input(45);
output(2, 242) <= input(43);
output(2, 243) <= input(41);
output(2, 244) <= input(39);
output(2, 245) <= input(37);
output(2, 246) <= input(35);
output(2, 247) <= input(33);
output(2, 248) <= input(16);
output(2, 249) <= input(17);
output(2, 250) <= input(18);
output(2, 251) <= input(19);
output(2, 252) <= input(20);
output(2, 253) <= input(21);
output(2, 254) <= input(22);
output(2, 255) <= input(23);
when "0101" =>
output(0, 0) <= input(0);
output(0, 1) <= input(1);
output(0, 2) <= input(2);
output(0, 3) <= input(3);
output(0, 4) <= input(4);
output(0, 5) <= input(5);
output(0, 6) <= input(6);
output(0, 7) <= input(7);
output(0, 8) <= input(8);
output(0, 9) <= input(9);
output(0, 10) <= input(10);
output(0, 11) <= input(11);
output(0, 12) <= input(12);
output(0, 13) <= input(13);
output(0, 14) <= input(14);
output(0, 15) <= input(15);
output(0, 16) <= input(16);
output(0, 17) <= input(17);
output(0, 18) <= input(18);
output(0, 19) <= input(19);
output(0, 20) <= input(20);
output(0, 21) <= input(21);
output(0, 22) <= input(22);
output(0, 23) <= input(23);
output(0, 24) <= input(24);
output(0, 25) <= input(25);
output(0, 26) <= input(26);
output(0, 27) <= input(27);
output(0, 28) <= input(28);
output(0, 29) <= input(29);
output(0, 30) <= input(30);
output(0, 31) <= input(31);
output(0, 32) <= input(32);
output(0, 33) <= input(0);
output(0, 34) <= input(1);
output(0, 35) <= input(2);
output(0, 36) <= input(3);
output(0, 37) <= input(4);
output(0, 38) <= input(5);
output(0, 39) <= input(6);
output(0, 40) <= input(7);
output(0, 41) <= input(8);
output(0, 42) <= input(9);
output(0, 43) <= input(10);
output(0, 44) <= input(11);
output(0, 45) <= input(12);
output(0, 46) <= input(13);
output(0, 47) <= input(14);
output(0, 48) <= input(33);
output(0, 49) <= input(16);
output(0, 50) <= input(17);
output(0, 51) <= input(18);
output(0, 52) <= input(19);
output(0, 53) <= input(20);
output(0, 54) <= input(21);
output(0, 55) <= input(22);
output(0, 56) <= input(23);
output(0, 57) <= input(24);
output(0, 58) <= input(25);
output(0, 59) <= input(26);
output(0, 60) <= input(27);
output(0, 61) <= input(28);
output(0, 62) <= input(29);
output(0, 63) <= input(30);
output(0, 64) <= input(34);
output(0, 65) <= input(32);
output(0, 66) <= input(0);
output(0, 67) <= input(1);
output(0, 68) <= input(2);
output(0, 69) <= input(3);
output(0, 70) <= input(4);
output(0, 71) <= input(5);
output(0, 72) <= input(6);
output(0, 73) <= input(7);
output(0, 74) <= input(8);
output(0, 75) <= input(9);
output(0, 76) <= input(10);
output(0, 77) <= input(11);
output(0, 78) <= input(12);
output(0, 79) <= input(13);
output(0, 80) <= input(35);
output(0, 81) <= input(33);
output(0, 82) <= input(16);
output(0, 83) <= input(17);
output(0, 84) <= input(18);
output(0, 85) <= input(19);
output(0, 86) <= input(20);
output(0, 87) <= input(21);
output(0, 88) <= input(22);
output(0, 89) <= input(23);
output(0, 90) <= input(24);
output(0, 91) <= input(25);
output(0, 92) <= input(26);
output(0, 93) <= input(27);
output(0, 94) <= input(28);
output(0, 95) <= input(29);
output(0, 96) <= input(36);
output(0, 97) <= input(34);
output(0, 98) <= input(32);
output(0, 99) <= input(0);
output(0, 100) <= input(1);
output(0, 101) <= input(2);
output(0, 102) <= input(3);
output(0, 103) <= input(4);
output(0, 104) <= input(5);
output(0, 105) <= input(6);
output(0, 106) <= input(7);
output(0, 107) <= input(8);
output(0, 108) <= input(9);
output(0, 109) <= input(10);
output(0, 110) <= input(11);
output(0, 111) <= input(12);
output(0, 112) <= input(37);
output(0, 113) <= input(35);
output(0, 114) <= input(33);
output(0, 115) <= input(16);
output(0, 116) <= input(17);
output(0, 117) <= input(18);
output(0, 118) <= input(19);
output(0, 119) <= input(20);
output(0, 120) <= input(21);
output(0, 121) <= input(22);
output(0, 122) <= input(23);
output(0, 123) <= input(24);
output(0, 124) <= input(25);
output(0, 125) <= input(26);
output(0, 126) <= input(27);
output(0, 127) <= input(28);
output(0, 128) <= input(38);
output(0, 129) <= input(36);
output(0, 130) <= input(34);
output(0, 131) <= input(32);
output(0, 132) <= input(0);
output(0, 133) <= input(1);
output(0, 134) <= input(2);
output(0, 135) <= input(3);
output(0, 136) <= input(4);
output(0, 137) <= input(5);
output(0, 138) <= input(6);
output(0, 139) <= input(7);
output(0, 140) <= input(8);
output(0, 141) <= input(9);
output(0, 142) <= input(10);
output(0, 143) <= input(11);
output(0, 144) <= input(39);
output(0, 145) <= input(37);
output(0, 146) <= input(35);
output(0, 147) <= input(33);
output(0, 148) <= input(16);
output(0, 149) <= input(17);
output(0, 150) <= input(18);
output(0, 151) <= input(19);
output(0, 152) <= input(20);
output(0, 153) <= input(21);
output(0, 154) <= input(22);
output(0, 155) <= input(23);
output(0, 156) <= input(24);
output(0, 157) <= input(25);
output(0, 158) <= input(26);
output(0, 159) <= input(27);
output(0, 160) <= input(40);
output(0, 161) <= input(38);
output(0, 162) <= input(36);
output(0, 163) <= input(34);
output(0, 164) <= input(32);
output(0, 165) <= input(0);
output(0, 166) <= input(1);
output(0, 167) <= input(2);
output(0, 168) <= input(3);
output(0, 169) <= input(4);
output(0, 170) <= input(5);
output(0, 171) <= input(6);
output(0, 172) <= input(7);
output(0, 173) <= input(8);
output(0, 174) <= input(9);
output(0, 175) <= input(10);
output(0, 176) <= input(41);
output(0, 177) <= input(39);
output(0, 178) <= input(37);
output(0, 179) <= input(35);
output(0, 180) <= input(33);
output(0, 181) <= input(16);
output(0, 182) <= input(17);
output(0, 183) <= input(18);
output(0, 184) <= input(19);
output(0, 185) <= input(20);
output(0, 186) <= input(21);
output(0, 187) <= input(22);
output(0, 188) <= input(23);
output(0, 189) <= input(24);
output(0, 190) <= input(25);
output(0, 191) <= input(26);
output(0, 192) <= input(42);
output(0, 193) <= input(40);
output(0, 194) <= input(38);
output(0, 195) <= input(36);
output(0, 196) <= input(34);
output(0, 197) <= input(32);
output(0, 198) <= input(0);
output(0, 199) <= input(1);
output(0, 200) <= input(2);
output(0, 201) <= input(3);
output(0, 202) <= input(4);
output(0, 203) <= input(5);
output(0, 204) <= input(6);
output(0, 205) <= input(7);
output(0, 206) <= input(8);
output(0, 207) <= input(9);
output(0, 208) <= input(43);
output(0, 209) <= input(41);
output(0, 210) <= input(39);
output(0, 211) <= input(37);
output(0, 212) <= input(35);
output(0, 213) <= input(33);
output(0, 214) <= input(16);
output(0, 215) <= input(17);
output(0, 216) <= input(18);
output(0, 217) <= input(19);
output(0, 218) <= input(20);
output(0, 219) <= input(21);
output(0, 220) <= input(22);
output(0, 221) <= input(23);
output(0, 222) <= input(24);
output(0, 223) <= input(25);
output(0, 224) <= input(44);
output(0, 225) <= input(42);
output(0, 226) <= input(40);
output(0, 227) <= input(38);
output(0, 228) <= input(36);
output(0, 229) <= input(34);
output(0, 230) <= input(32);
output(0, 231) <= input(0);
output(0, 232) <= input(1);
output(0, 233) <= input(2);
output(0, 234) <= input(3);
output(0, 235) <= input(4);
output(0, 236) <= input(5);
output(0, 237) <= input(6);
output(0, 238) <= input(7);
output(0, 239) <= input(8);
output(0, 240) <= input(45);
output(0, 241) <= input(43);
output(0, 242) <= input(41);
output(0, 243) <= input(39);
output(0, 244) <= input(37);
output(0, 245) <= input(35);
output(0, 246) <= input(33);
output(0, 247) <= input(16);
output(0, 248) <= input(17);
output(0, 249) <= input(18);
output(0, 250) <= input(19);
output(0, 251) <= input(20);
output(0, 252) <= input(21);
output(0, 253) <= input(22);
output(0, 254) <= input(23);
output(0, 255) <= input(24);
output(1, 0) <= input(33);
output(1, 1) <= input(16);
output(1, 2) <= input(17);
output(1, 3) <= input(18);
output(1, 4) <= input(19);
output(1, 5) <= input(20);
output(1, 6) <= input(21);
output(1, 7) <= input(22);
output(1, 8) <= input(23);
output(1, 9) <= input(24);
output(1, 10) <= input(25);
output(1, 11) <= input(26);
output(1, 12) <= input(27);
output(1, 13) <= input(28);
output(1, 14) <= input(29);
output(1, 15) <= input(30);
output(1, 16) <= input(34);
output(1, 17) <= input(32);
output(1, 18) <= input(0);
output(1, 19) <= input(1);
output(1, 20) <= input(2);
output(1, 21) <= input(3);
output(1, 22) <= input(4);
output(1, 23) <= input(5);
output(1, 24) <= input(6);
output(1, 25) <= input(7);
output(1, 26) <= input(8);
output(1, 27) <= input(9);
output(1, 28) <= input(10);
output(1, 29) <= input(11);
output(1, 30) <= input(12);
output(1, 31) <= input(13);
output(1, 32) <= input(35);
output(1, 33) <= input(33);
output(1, 34) <= input(16);
output(1, 35) <= input(17);
output(1, 36) <= input(18);
output(1, 37) <= input(19);
output(1, 38) <= input(20);
output(1, 39) <= input(21);
output(1, 40) <= input(22);
output(1, 41) <= input(23);
output(1, 42) <= input(24);
output(1, 43) <= input(25);
output(1, 44) <= input(26);
output(1, 45) <= input(27);
output(1, 46) <= input(28);
output(1, 47) <= input(29);
output(1, 48) <= input(36);
output(1, 49) <= input(34);
output(1, 50) <= input(32);
output(1, 51) <= input(0);
output(1, 52) <= input(1);
output(1, 53) <= input(2);
output(1, 54) <= input(3);
output(1, 55) <= input(4);
output(1, 56) <= input(5);
output(1, 57) <= input(6);
output(1, 58) <= input(7);
output(1, 59) <= input(8);
output(1, 60) <= input(9);
output(1, 61) <= input(10);
output(1, 62) <= input(11);
output(1, 63) <= input(12);
output(1, 64) <= input(37);
output(1, 65) <= input(35);
output(1, 66) <= input(33);
output(1, 67) <= input(16);
output(1, 68) <= input(17);
output(1, 69) <= input(18);
output(1, 70) <= input(19);
output(1, 71) <= input(20);
output(1, 72) <= input(21);
output(1, 73) <= input(22);
output(1, 74) <= input(23);
output(1, 75) <= input(24);
output(1, 76) <= input(25);
output(1, 77) <= input(26);
output(1, 78) <= input(27);
output(1, 79) <= input(28);
output(1, 80) <= input(38);
output(1, 81) <= input(36);
output(1, 82) <= input(34);
output(1, 83) <= input(32);
output(1, 84) <= input(0);
output(1, 85) <= input(1);
output(1, 86) <= input(2);
output(1, 87) <= input(3);
output(1, 88) <= input(4);
output(1, 89) <= input(5);
output(1, 90) <= input(6);
output(1, 91) <= input(7);
output(1, 92) <= input(8);
output(1, 93) <= input(9);
output(1, 94) <= input(10);
output(1, 95) <= input(11);
output(1, 96) <= input(39);
output(1, 97) <= input(37);
output(1, 98) <= input(35);
output(1, 99) <= input(33);
output(1, 100) <= input(16);
output(1, 101) <= input(17);
output(1, 102) <= input(18);
output(1, 103) <= input(19);
output(1, 104) <= input(20);
output(1, 105) <= input(21);
output(1, 106) <= input(22);
output(1, 107) <= input(23);
output(1, 108) <= input(24);
output(1, 109) <= input(25);
output(1, 110) <= input(26);
output(1, 111) <= input(27);
output(1, 112) <= input(40);
output(1, 113) <= input(38);
output(1, 114) <= input(36);
output(1, 115) <= input(34);
output(1, 116) <= input(32);
output(1, 117) <= input(0);
output(1, 118) <= input(1);
output(1, 119) <= input(2);
output(1, 120) <= input(3);
output(1, 121) <= input(4);
output(1, 122) <= input(5);
output(1, 123) <= input(6);
output(1, 124) <= input(7);
output(1, 125) <= input(8);
output(1, 126) <= input(9);
output(1, 127) <= input(10);
output(1, 128) <= input(42);
output(1, 129) <= input(40);
output(1, 130) <= input(38);
output(1, 131) <= input(36);
output(1, 132) <= input(34);
output(1, 133) <= input(32);
output(1, 134) <= input(0);
output(1, 135) <= input(1);
output(1, 136) <= input(2);
output(1, 137) <= input(3);
output(1, 138) <= input(4);
output(1, 139) <= input(5);
output(1, 140) <= input(6);
output(1, 141) <= input(7);
output(1, 142) <= input(8);
output(1, 143) <= input(9);
output(1, 144) <= input(43);
output(1, 145) <= input(41);
output(1, 146) <= input(39);
output(1, 147) <= input(37);
output(1, 148) <= input(35);
output(1, 149) <= input(33);
output(1, 150) <= input(16);
output(1, 151) <= input(17);
output(1, 152) <= input(18);
output(1, 153) <= input(19);
output(1, 154) <= input(20);
output(1, 155) <= input(21);
output(1, 156) <= input(22);
output(1, 157) <= input(23);
output(1, 158) <= input(24);
output(1, 159) <= input(25);
output(1, 160) <= input(44);
output(1, 161) <= input(42);
output(1, 162) <= input(40);
output(1, 163) <= input(38);
output(1, 164) <= input(36);
output(1, 165) <= input(34);
output(1, 166) <= input(32);
output(1, 167) <= input(0);
output(1, 168) <= input(1);
output(1, 169) <= input(2);
output(1, 170) <= input(3);
output(1, 171) <= input(4);
output(1, 172) <= input(5);
output(1, 173) <= input(6);
output(1, 174) <= input(7);
output(1, 175) <= input(8);
output(1, 176) <= input(45);
output(1, 177) <= input(43);
output(1, 178) <= input(41);
output(1, 179) <= input(39);
output(1, 180) <= input(37);
output(1, 181) <= input(35);
output(1, 182) <= input(33);
output(1, 183) <= input(16);
output(1, 184) <= input(17);
output(1, 185) <= input(18);
output(1, 186) <= input(19);
output(1, 187) <= input(20);
output(1, 188) <= input(21);
output(1, 189) <= input(22);
output(1, 190) <= input(23);
output(1, 191) <= input(24);
output(1, 192) <= input(46);
output(1, 193) <= input(44);
output(1, 194) <= input(42);
output(1, 195) <= input(40);
output(1, 196) <= input(38);
output(1, 197) <= input(36);
output(1, 198) <= input(34);
output(1, 199) <= input(32);
output(1, 200) <= input(0);
output(1, 201) <= input(1);
output(1, 202) <= input(2);
output(1, 203) <= input(3);
output(1, 204) <= input(4);
output(1, 205) <= input(5);
output(1, 206) <= input(6);
output(1, 207) <= input(7);
output(1, 208) <= input(47);
output(1, 209) <= input(45);
output(1, 210) <= input(43);
output(1, 211) <= input(41);
output(1, 212) <= input(39);
output(1, 213) <= input(37);
output(1, 214) <= input(35);
output(1, 215) <= input(33);
output(1, 216) <= input(16);
output(1, 217) <= input(17);
output(1, 218) <= input(18);
output(1, 219) <= input(19);
output(1, 220) <= input(20);
output(1, 221) <= input(21);
output(1, 222) <= input(22);
output(1, 223) <= input(23);
output(1, 224) <= input(48);
output(1, 225) <= input(46);
output(1, 226) <= input(44);
output(1, 227) <= input(42);
output(1, 228) <= input(40);
output(1, 229) <= input(38);
output(1, 230) <= input(36);
output(1, 231) <= input(34);
output(1, 232) <= input(32);
output(1, 233) <= input(0);
output(1, 234) <= input(1);
output(1, 235) <= input(2);
output(1, 236) <= input(3);
output(1, 237) <= input(4);
output(1, 238) <= input(5);
output(1, 239) <= input(6);
output(1, 240) <= input(49);
output(1, 241) <= input(47);
output(1, 242) <= input(45);
output(1, 243) <= input(43);
output(1, 244) <= input(41);
output(1, 245) <= input(39);
output(1, 246) <= input(37);
output(1, 247) <= input(35);
output(1, 248) <= input(33);
output(1, 249) <= input(16);
output(1, 250) <= input(17);
output(1, 251) <= input(18);
output(1, 252) <= input(19);
output(1, 253) <= input(20);
output(1, 254) <= input(21);
output(1, 255) <= input(22);
when "0110" =>
output(0, 0) <= input(0);
output(0, 1) <= input(1);
output(0, 2) <= input(2);
output(0, 3) <= input(3);
output(0, 4) <= input(4);
output(0, 5) <= input(5);
output(0, 6) <= input(6);
output(0, 7) <= input(7);
output(0, 8) <= input(8);
output(0, 9) <= input(9);
output(0, 10) <= input(10);
output(0, 11) <= input(11);
output(0, 12) <= input(12);
output(0, 13) <= input(13);
output(0, 14) <= input(14);
output(0, 15) <= input(15);
output(0, 16) <= input(16);
output(0, 17) <= input(17);
output(0, 18) <= input(18);
output(0, 19) <= input(19);
output(0, 20) <= input(20);
output(0, 21) <= input(21);
output(0, 22) <= input(22);
output(0, 23) <= input(23);
output(0, 24) <= input(24);
output(0, 25) <= input(25);
output(0, 26) <= input(26);
output(0, 27) <= input(27);
output(0, 28) <= input(28);
output(0, 29) <= input(29);
output(0, 30) <= input(30);
output(0, 31) <= input(31);
output(0, 32) <= input(32);
output(0, 33) <= input(0);
output(0, 34) <= input(1);
output(0, 35) <= input(2);
output(0, 36) <= input(3);
output(0, 37) <= input(4);
output(0, 38) <= input(5);
output(0, 39) <= input(6);
output(0, 40) <= input(7);
output(0, 41) <= input(8);
output(0, 42) <= input(9);
output(0, 43) <= input(10);
output(0, 44) <= input(11);
output(0, 45) <= input(12);
output(0, 46) <= input(13);
output(0, 47) <= input(14);
output(0, 48) <= input(33);
output(0, 49) <= input(16);
output(0, 50) <= input(17);
output(0, 51) <= input(18);
output(0, 52) <= input(19);
output(0, 53) <= input(20);
output(0, 54) <= input(21);
output(0, 55) <= input(22);
output(0, 56) <= input(23);
output(0, 57) <= input(24);
output(0, 58) <= input(25);
output(0, 59) <= input(26);
output(0, 60) <= input(27);
output(0, 61) <= input(28);
output(0, 62) <= input(29);
output(0, 63) <= input(30);
output(0, 64) <= input(34);
output(0, 65) <= input(33);
output(0, 66) <= input(16);
output(0, 67) <= input(17);
output(0, 68) <= input(18);
output(0, 69) <= input(19);
output(0, 70) <= input(20);
output(0, 71) <= input(21);
output(0, 72) <= input(22);
output(0, 73) <= input(23);
output(0, 74) <= input(24);
output(0, 75) <= input(25);
output(0, 76) <= input(26);
output(0, 77) <= input(27);
output(0, 78) <= input(28);
output(0, 79) <= input(29);
output(0, 80) <= input(35);
output(0, 81) <= input(36);
output(0, 82) <= input(32);
output(0, 83) <= input(0);
output(0, 84) <= input(1);
output(0, 85) <= input(2);
output(0, 86) <= input(3);
output(0, 87) <= input(4);
output(0, 88) <= input(5);
output(0, 89) <= input(6);
output(0, 90) <= input(7);
output(0, 91) <= input(8);
output(0, 92) <= input(9);
output(0, 93) <= input(10);
output(0, 94) <= input(11);
output(0, 95) <= input(12);
output(0, 96) <= input(37);
output(0, 97) <= input(34);
output(0, 98) <= input(33);
output(0, 99) <= input(16);
output(0, 100) <= input(17);
output(0, 101) <= input(18);
output(0, 102) <= input(19);
output(0, 103) <= input(20);
output(0, 104) <= input(21);
output(0, 105) <= input(22);
output(0, 106) <= input(23);
output(0, 107) <= input(24);
output(0, 108) <= input(25);
output(0, 109) <= input(26);
output(0, 110) <= input(27);
output(0, 111) <= input(28);
output(0, 112) <= input(38);
output(0, 113) <= input(35);
output(0, 114) <= input(36);
output(0, 115) <= input(32);
output(0, 116) <= input(0);
output(0, 117) <= input(1);
output(0, 118) <= input(2);
output(0, 119) <= input(3);
output(0, 120) <= input(4);
output(0, 121) <= input(5);
output(0, 122) <= input(6);
output(0, 123) <= input(7);
output(0, 124) <= input(8);
output(0, 125) <= input(9);
output(0, 126) <= input(10);
output(0, 127) <= input(11);
output(0, 128) <= input(39);
output(0, 129) <= input(38);
output(0, 130) <= input(35);
output(0, 131) <= input(36);
output(0, 132) <= input(32);
output(0, 133) <= input(0);
output(0, 134) <= input(1);
output(0, 135) <= input(2);
output(0, 136) <= input(3);
output(0, 137) <= input(4);
output(0, 138) <= input(5);
output(0, 139) <= input(6);
output(0, 140) <= input(7);
output(0, 141) <= input(8);
output(0, 142) <= input(9);
output(0, 143) <= input(10);
output(0, 144) <= input(40);
output(0, 145) <= input(41);
output(0, 146) <= input(37);
output(0, 147) <= input(34);
output(0, 148) <= input(33);
output(0, 149) <= input(16);
output(0, 150) <= input(17);
output(0, 151) <= input(18);
output(0, 152) <= input(19);
output(0, 153) <= input(20);
output(0, 154) <= input(21);
output(0, 155) <= input(22);
output(0, 156) <= input(23);
output(0, 157) <= input(24);
output(0, 158) <= input(25);
output(0, 159) <= input(26);
output(0, 160) <= input(42);
output(0, 161) <= input(39);
output(0, 162) <= input(38);
output(0, 163) <= input(35);
output(0, 164) <= input(36);
output(0, 165) <= input(32);
output(0, 166) <= input(0);
output(0, 167) <= input(1);
output(0, 168) <= input(2);
output(0, 169) <= input(3);
output(0, 170) <= input(4);
output(0, 171) <= input(5);
output(0, 172) <= input(6);
output(0, 173) <= input(7);
output(0, 174) <= input(8);
output(0, 175) <= input(9);
output(0, 176) <= input(43);
output(0, 177) <= input(40);
output(0, 178) <= input(41);
output(0, 179) <= input(37);
output(0, 180) <= input(34);
output(0, 181) <= input(33);
output(0, 182) <= input(16);
output(0, 183) <= input(17);
output(0, 184) <= input(18);
output(0, 185) <= input(19);
output(0, 186) <= input(20);
output(0, 187) <= input(21);
output(0, 188) <= input(22);
output(0, 189) <= input(23);
output(0, 190) <= input(24);
output(0, 191) <= input(25);
output(0, 192) <= input(44);
output(0, 193) <= input(43);
output(0, 194) <= input(40);
output(0, 195) <= input(41);
output(0, 196) <= input(37);
output(0, 197) <= input(34);
output(0, 198) <= input(33);
output(0, 199) <= input(16);
output(0, 200) <= input(17);
output(0, 201) <= input(18);
output(0, 202) <= input(19);
output(0, 203) <= input(20);
output(0, 204) <= input(21);
output(0, 205) <= input(22);
output(0, 206) <= input(23);
output(0, 207) <= input(24);
output(0, 208) <= input(45);
output(0, 209) <= input(46);
output(0, 210) <= input(42);
output(0, 211) <= input(39);
output(0, 212) <= input(38);
output(0, 213) <= input(35);
output(0, 214) <= input(36);
output(0, 215) <= input(32);
output(0, 216) <= input(0);
output(0, 217) <= input(1);
output(0, 218) <= input(2);
output(0, 219) <= input(3);
output(0, 220) <= input(4);
output(0, 221) <= input(5);
output(0, 222) <= input(6);
output(0, 223) <= input(7);
output(0, 224) <= input(47);
output(0, 225) <= input(44);
output(0, 226) <= input(43);
output(0, 227) <= input(40);
output(0, 228) <= input(41);
output(0, 229) <= input(37);
output(0, 230) <= input(34);
output(0, 231) <= input(33);
output(0, 232) <= input(16);
output(0, 233) <= input(17);
output(0, 234) <= input(18);
output(0, 235) <= input(19);
output(0, 236) <= input(20);
output(0, 237) <= input(21);
output(0, 238) <= input(22);
output(0, 239) <= input(23);
output(0, 240) <= input(48);
output(0, 241) <= input(45);
output(0, 242) <= input(46);
output(0, 243) <= input(42);
output(0, 244) <= input(39);
output(0, 245) <= input(38);
output(0, 246) <= input(35);
output(0, 247) <= input(36);
output(0, 248) <= input(32);
output(0, 249) <= input(0);
output(0, 250) <= input(1);
output(0, 251) <= input(2);
output(0, 252) <= input(3);
output(0, 253) <= input(4);
output(0, 254) <= input(5);
output(0, 255) <= input(6);
output(1, 0) <= input(33);
output(1, 1) <= input(16);
output(1, 2) <= input(17);
output(1, 3) <= input(18);
output(1, 4) <= input(19);
output(1, 5) <= input(20);
output(1, 6) <= input(21);
output(1, 7) <= input(22);
output(1, 8) <= input(23);
output(1, 9) <= input(24);
output(1, 10) <= input(25);
output(1, 11) <= input(26);
output(1, 12) <= input(27);
output(1, 13) <= input(28);
output(1, 14) <= input(29);
output(1, 15) <= input(30);
output(1, 16) <= input(36);
output(1, 17) <= input(32);
output(1, 18) <= input(0);
output(1, 19) <= input(1);
output(1, 20) <= input(2);
output(1, 21) <= input(3);
output(1, 22) <= input(4);
output(1, 23) <= input(5);
output(1, 24) <= input(6);
output(1, 25) <= input(7);
output(1, 26) <= input(8);
output(1, 27) <= input(9);
output(1, 28) <= input(10);
output(1, 29) <= input(11);
output(1, 30) <= input(12);
output(1, 31) <= input(13);
output(1, 32) <= input(35);
output(1, 33) <= input(36);
output(1, 34) <= input(32);
output(1, 35) <= input(0);
output(1, 36) <= input(1);
output(1, 37) <= input(2);
output(1, 38) <= input(3);
output(1, 39) <= input(4);
output(1, 40) <= input(5);
output(1, 41) <= input(6);
output(1, 42) <= input(7);
output(1, 43) <= input(8);
output(1, 44) <= input(9);
output(1, 45) <= input(10);
output(1, 46) <= input(11);
output(1, 47) <= input(12);
output(1, 48) <= input(37);
output(1, 49) <= input(34);
output(1, 50) <= input(33);
output(1, 51) <= input(16);
output(1, 52) <= input(17);
output(1, 53) <= input(18);
output(1, 54) <= input(19);
output(1, 55) <= input(20);
output(1, 56) <= input(21);
output(1, 57) <= input(22);
output(1, 58) <= input(23);
output(1, 59) <= input(24);
output(1, 60) <= input(25);
output(1, 61) <= input(26);
output(1, 62) <= input(27);
output(1, 63) <= input(28);
output(1, 64) <= input(41);
output(1, 65) <= input(37);
output(1, 66) <= input(34);
output(1, 67) <= input(33);
output(1, 68) <= input(16);
output(1, 69) <= input(17);
output(1, 70) <= input(18);
output(1, 71) <= input(19);
output(1, 72) <= input(20);
output(1, 73) <= input(21);
output(1, 74) <= input(22);
output(1, 75) <= input(23);
output(1, 76) <= input(24);
output(1, 77) <= input(25);
output(1, 78) <= input(26);
output(1, 79) <= input(27);
output(1, 80) <= input(39);
output(1, 81) <= input(38);
output(1, 82) <= input(35);
output(1, 83) <= input(36);
output(1, 84) <= input(32);
output(1, 85) <= input(0);
output(1, 86) <= input(1);
output(1, 87) <= input(2);
output(1, 88) <= input(3);
output(1, 89) <= input(4);
output(1, 90) <= input(5);
output(1, 91) <= input(6);
output(1, 92) <= input(7);
output(1, 93) <= input(8);
output(1, 94) <= input(9);
output(1, 95) <= input(10);
output(1, 96) <= input(42);
output(1, 97) <= input(39);
output(1, 98) <= input(38);
output(1, 99) <= input(35);
output(1, 100) <= input(36);
output(1, 101) <= input(32);
output(1, 102) <= input(0);
output(1, 103) <= input(1);
output(1, 104) <= input(2);
output(1, 105) <= input(3);
output(1, 106) <= input(4);
output(1, 107) <= input(5);
output(1, 108) <= input(6);
output(1, 109) <= input(7);
output(1, 110) <= input(8);
output(1, 111) <= input(9);
output(1, 112) <= input(43);
output(1, 113) <= input(40);
output(1, 114) <= input(41);
output(1, 115) <= input(37);
output(1, 116) <= input(34);
output(1, 117) <= input(33);
output(1, 118) <= input(16);
output(1, 119) <= input(17);
output(1, 120) <= input(18);
output(1, 121) <= input(19);
output(1, 122) <= input(20);
output(1, 123) <= input(21);
output(1, 124) <= input(22);
output(1, 125) <= input(23);
output(1, 126) <= input(24);
output(1, 127) <= input(25);
output(1, 128) <= input(46);
output(1, 129) <= input(42);
output(1, 130) <= input(39);
output(1, 131) <= input(38);
output(1, 132) <= input(35);
output(1, 133) <= input(36);
output(1, 134) <= input(32);
output(1, 135) <= input(0);
output(1, 136) <= input(1);
output(1, 137) <= input(2);
output(1, 138) <= input(3);
output(1, 139) <= input(4);
output(1, 140) <= input(5);
output(1, 141) <= input(6);
output(1, 142) <= input(7);
output(1, 143) <= input(8);
output(1, 144) <= input(45);
output(1, 145) <= input(46);
output(1, 146) <= input(42);
output(1, 147) <= input(39);
output(1, 148) <= input(38);
output(1, 149) <= input(35);
output(1, 150) <= input(36);
output(1, 151) <= input(32);
output(1, 152) <= input(0);
output(1, 153) <= input(1);
output(1, 154) <= input(2);
output(1, 155) <= input(3);
output(1, 156) <= input(4);
output(1, 157) <= input(5);
output(1, 158) <= input(6);
output(1, 159) <= input(7);
output(1, 160) <= input(47);
output(1, 161) <= input(44);
output(1, 162) <= input(43);
output(1, 163) <= input(40);
output(1, 164) <= input(41);
output(1, 165) <= input(37);
output(1, 166) <= input(34);
output(1, 167) <= input(33);
output(1, 168) <= input(16);
output(1, 169) <= input(17);
output(1, 170) <= input(18);
output(1, 171) <= input(19);
output(1, 172) <= input(20);
output(1, 173) <= input(21);
output(1, 174) <= input(22);
output(1, 175) <= input(23);
output(1, 176) <= input(49);
output(1, 177) <= input(47);
output(1, 178) <= input(44);
output(1, 179) <= input(43);
output(1, 180) <= input(40);
output(1, 181) <= input(41);
output(1, 182) <= input(37);
output(1, 183) <= input(34);
output(1, 184) <= input(33);
output(1, 185) <= input(16);
output(1, 186) <= input(17);
output(1, 187) <= input(18);
output(1, 188) <= input(19);
output(1, 189) <= input(20);
output(1, 190) <= input(21);
output(1, 191) <= input(22);
output(1, 192) <= input(50);
output(1, 193) <= input(48);
output(1, 194) <= input(45);
output(1, 195) <= input(46);
output(1, 196) <= input(42);
output(1, 197) <= input(39);
output(1, 198) <= input(38);
output(1, 199) <= input(35);
output(1, 200) <= input(36);
output(1, 201) <= input(32);
output(1, 202) <= input(0);
output(1, 203) <= input(1);
output(1, 204) <= input(2);
output(1, 205) <= input(3);
output(1, 206) <= input(4);
output(1, 207) <= input(5);
output(1, 208) <= input(51);
output(1, 209) <= input(50);
output(1, 210) <= input(48);
output(1, 211) <= input(45);
output(1, 212) <= input(46);
output(1, 213) <= input(42);
output(1, 214) <= input(39);
output(1, 215) <= input(38);
output(1, 216) <= input(35);
output(1, 217) <= input(36);
output(1, 218) <= input(32);
output(1, 219) <= input(0);
output(1, 220) <= input(1);
output(1, 221) <= input(2);
output(1, 222) <= input(3);
output(1, 223) <= input(4);
output(1, 224) <= input(52);
output(1, 225) <= input(53);
output(1, 226) <= input(49);
output(1, 227) <= input(47);
output(1, 228) <= input(44);
output(1, 229) <= input(43);
output(1, 230) <= input(40);
output(1, 231) <= input(41);
output(1, 232) <= input(37);
output(1, 233) <= input(34);
output(1, 234) <= input(33);
output(1, 235) <= input(16);
output(1, 236) <= input(17);
output(1, 237) <= input(18);
output(1, 238) <= input(19);
output(1, 239) <= input(20);
output(1, 240) <= input(54);
output(1, 241) <= input(51);
output(1, 242) <= input(50);
output(1, 243) <= input(48);
output(1, 244) <= input(45);
output(1, 245) <= input(46);
output(1, 246) <= input(42);
output(1, 247) <= input(39);
output(1, 248) <= input(38);
output(1, 249) <= input(35);
output(1, 250) <= input(36);
output(1, 251) <= input(32);
output(1, 252) <= input(0);
output(1, 253) <= input(1);
output(1, 254) <= input(2);
output(1, 255) <= input(3);
output(2, 0) <= input(35);
output(2, 1) <= input(36);
output(2, 2) <= input(32);
output(2, 3) <= input(0);
output(2, 4) <= input(1);
output(2, 5) <= input(2);
output(2, 6) <= input(3);
output(2, 7) <= input(4);
output(2, 8) <= input(5);
output(2, 9) <= input(6);
output(2, 10) <= input(7);
output(2, 11) <= input(8);
output(2, 12) <= input(9);
output(2, 13) <= input(10);
output(2, 14) <= input(11);
output(2, 15) <= input(12);
output(2, 16) <= input(38);
output(2, 17) <= input(35);
output(2, 18) <= input(36);
output(2, 19) <= input(32);
output(2, 20) <= input(0);
output(2, 21) <= input(1);
output(2, 22) <= input(2);
output(2, 23) <= input(3);
output(2, 24) <= input(4);
output(2, 25) <= input(5);
output(2, 26) <= input(6);
output(2, 27) <= input(7);
output(2, 28) <= input(8);
output(2, 29) <= input(9);
output(2, 30) <= input(10);
output(2, 31) <= input(11);
output(2, 32) <= input(41);
output(2, 33) <= input(37);
output(2, 34) <= input(34);
output(2, 35) <= input(33);
output(2, 36) <= input(16);
output(2, 37) <= input(17);
output(2, 38) <= input(18);
output(2, 39) <= input(19);
output(2, 40) <= input(20);
output(2, 41) <= input(21);
output(2, 42) <= input(22);
output(2, 43) <= input(23);
output(2, 44) <= input(24);
output(2, 45) <= input(25);
output(2, 46) <= input(26);
output(2, 47) <= input(27);
output(2, 48) <= input(40);
output(2, 49) <= input(41);
output(2, 50) <= input(37);
output(2, 51) <= input(34);
output(2, 52) <= input(33);
output(2, 53) <= input(16);
output(2, 54) <= input(17);
output(2, 55) <= input(18);
output(2, 56) <= input(19);
output(2, 57) <= input(20);
output(2, 58) <= input(21);
output(2, 59) <= input(22);
output(2, 60) <= input(23);
output(2, 61) <= input(24);
output(2, 62) <= input(25);
output(2, 63) <= input(26);
output(2, 64) <= input(43);
output(2, 65) <= input(40);
output(2, 66) <= input(41);
output(2, 67) <= input(37);
output(2, 68) <= input(34);
output(2, 69) <= input(33);
output(2, 70) <= input(16);
output(2, 71) <= input(17);
output(2, 72) <= input(18);
output(2, 73) <= input(19);
output(2, 74) <= input(20);
output(2, 75) <= input(21);
output(2, 76) <= input(22);
output(2, 77) <= input(23);
output(2, 78) <= input(24);
output(2, 79) <= input(25);
output(2, 80) <= input(46);
output(2, 81) <= input(42);
output(2, 82) <= input(39);
output(2, 83) <= input(38);
output(2, 84) <= input(35);
output(2, 85) <= input(36);
output(2, 86) <= input(32);
output(2, 87) <= input(0);
output(2, 88) <= input(1);
output(2, 89) <= input(2);
output(2, 90) <= input(3);
output(2, 91) <= input(4);
output(2, 92) <= input(5);
output(2, 93) <= input(6);
output(2, 94) <= input(7);
output(2, 95) <= input(8);
output(2, 96) <= input(45);
output(2, 97) <= input(46);
output(2, 98) <= input(42);
output(2, 99) <= input(39);
output(2, 100) <= input(38);
output(2, 101) <= input(35);
output(2, 102) <= input(36);
output(2, 103) <= input(32);
output(2, 104) <= input(0);
output(2, 105) <= input(1);
output(2, 106) <= input(2);
output(2, 107) <= input(3);
output(2, 108) <= input(4);
output(2, 109) <= input(5);
output(2, 110) <= input(6);
output(2, 111) <= input(7);
output(2, 112) <= input(47);
output(2, 113) <= input(44);
output(2, 114) <= input(43);
output(2, 115) <= input(40);
output(2, 116) <= input(41);
output(2, 117) <= input(37);
output(2, 118) <= input(34);
output(2, 119) <= input(33);
output(2, 120) <= input(16);
output(2, 121) <= input(17);
output(2, 122) <= input(18);
output(2, 123) <= input(19);
output(2, 124) <= input(20);
output(2, 125) <= input(21);
output(2, 126) <= input(22);
output(2, 127) <= input(23);
output(2, 128) <= input(49);
output(2, 129) <= input(47);
output(2, 130) <= input(44);
output(2, 131) <= input(43);
output(2, 132) <= input(40);
output(2, 133) <= input(41);
output(2, 134) <= input(37);
output(2, 135) <= input(34);
output(2, 136) <= input(33);
output(2, 137) <= input(16);
output(2, 138) <= input(17);
output(2, 139) <= input(18);
output(2, 140) <= input(19);
output(2, 141) <= input(20);
output(2, 142) <= input(21);
output(2, 143) <= input(22);
output(2, 144) <= input(53);
output(2, 145) <= input(49);
output(2, 146) <= input(47);
output(2, 147) <= input(44);
output(2, 148) <= input(43);
output(2, 149) <= input(40);
output(2, 150) <= input(41);
output(2, 151) <= input(37);
output(2, 152) <= input(34);
output(2, 153) <= input(33);
output(2, 154) <= input(16);
output(2, 155) <= input(17);
output(2, 156) <= input(18);
output(2, 157) <= input(19);
output(2, 158) <= input(20);
output(2, 159) <= input(21);
output(2, 160) <= input(51);
output(2, 161) <= input(50);
output(2, 162) <= input(48);
output(2, 163) <= input(45);
output(2, 164) <= input(46);
output(2, 165) <= input(42);
output(2, 166) <= input(39);
output(2, 167) <= input(38);
output(2, 168) <= input(35);
output(2, 169) <= input(36);
output(2, 170) <= input(32);
output(2, 171) <= input(0);
output(2, 172) <= input(1);
output(2, 173) <= input(2);
output(2, 174) <= input(3);
output(2, 175) <= input(4);
output(2, 176) <= input(54);
output(2, 177) <= input(51);
output(2, 178) <= input(50);
output(2, 179) <= input(48);
output(2, 180) <= input(45);
output(2, 181) <= input(46);
output(2, 182) <= input(42);
output(2, 183) <= input(39);
output(2, 184) <= input(38);
output(2, 185) <= input(35);
output(2, 186) <= input(36);
output(2, 187) <= input(32);
output(2, 188) <= input(0);
output(2, 189) <= input(1);
output(2, 190) <= input(2);
output(2, 191) <= input(3);
output(2, 192) <= input(55);
output(2, 193) <= input(54);
output(2, 194) <= input(51);
output(2, 195) <= input(50);
output(2, 196) <= input(48);
output(2, 197) <= input(45);
output(2, 198) <= input(46);
output(2, 199) <= input(42);
output(2, 200) <= input(39);
output(2, 201) <= input(38);
output(2, 202) <= input(35);
output(2, 203) <= input(36);
output(2, 204) <= input(32);
output(2, 205) <= input(0);
output(2, 206) <= input(1);
output(2, 207) <= input(2);
output(2, 208) <= input(56);
output(2, 209) <= input(57);
output(2, 210) <= input(52);
output(2, 211) <= input(53);
output(2, 212) <= input(49);
output(2, 213) <= input(47);
output(2, 214) <= input(44);
output(2, 215) <= input(43);
output(2, 216) <= input(40);
output(2, 217) <= input(41);
output(2, 218) <= input(37);
output(2, 219) <= input(34);
output(2, 220) <= input(33);
output(2, 221) <= input(16);
output(2, 222) <= input(17);
output(2, 223) <= input(18);
output(2, 224) <= input(58);
output(2, 225) <= input(56);
output(2, 226) <= input(57);
output(2, 227) <= input(52);
output(2, 228) <= input(53);
output(2, 229) <= input(49);
output(2, 230) <= input(47);
output(2, 231) <= input(44);
output(2, 232) <= input(43);
output(2, 233) <= input(40);
output(2, 234) <= input(41);
output(2, 235) <= input(37);
output(2, 236) <= input(34);
output(2, 237) <= input(33);
output(2, 238) <= input(16);
output(2, 239) <= input(17);
output(2, 240) <= input(59);
output(2, 241) <= input(60);
output(2, 242) <= input(55);
output(2, 243) <= input(54);
output(2, 244) <= input(51);
output(2, 245) <= input(50);
output(2, 246) <= input(48);
output(2, 247) <= input(45);
output(2, 248) <= input(46);
output(2, 249) <= input(42);
output(2, 250) <= input(39);
output(2, 251) <= input(38);
output(2, 252) <= input(35);
output(2, 253) <= input(36);
output(2, 254) <= input(32);
output(2, 255) <= input(0);
when "0111" =>
output(0, 0) <= input(0);
output(0, 1) <= input(1);
output(0, 2) <= input(2);
output(0, 3) <= input(3);
output(0, 4) <= input(4);
output(0, 5) <= input(5);
output(0, 6) <= input(6);
output(0, 7) <= input(7);
output(0, 8) <= input(8);
output(0, 9) <= input(9);
output(0, 10) <= input(10);
output(0, 11) <= input(11);
output(0, 12) <= input(12);
output(0, 13) <= input(13);
output(0, 14) <= input(14);
output(0, 15) <= input(15);
output(0, 16) <= input(16);
output(0, 17) <= input(0);
output(0, 18) <= input(1);
output(0, 19) <= input(2);
output(0, 20) <= input(3);
output(0, 21) <= input(4);
output(0, 22) <= input(5);
output(0, 23) <= input(6);
output(0, 24) <= input(7);
output(0, 25) <= input(8);
output(0, 26) <= input(9);
output(0, 27) <= input(10);
output(0, 28) <= input(11);
output(0, 29) <= input(12);
output(0, 30) <= input(13);
output(0, 31) <= input(14);
output(0, 32) <= input(17);
output(0, 33) <= input(16);
output(0, 34) <= input(0);
output(0, 35) <= input(1);
output(0, 36) <= input(2);
output(0, 37) <= input(3);
output(0, 38) <= input(4);
output(0, 39) <= input(5);
output(0, 40) <= input(6);
output(0, 41) <= input(7);
output(0, 42) <= input(8);
output(0, 43) <= input(9);
output(0, 44) <= input(10);
output(0, 45) <= input(11);
output(0, 46) <= input(12);
output(0, 47) <= input(13);
output(0, 48) <= input(18);
output(0, 49) <= input(17);
output(0, 50) <= input(16);
output(0, 51) <= input(0);
output(0, 52) <= input(1);
output(0, 53) <= input(2);
output(0, 54) <= input(3);
output(0, 55) <= input(4);
output(0, 56) <= input(5);
output(0, 57) <= input(6);
output(0, 58) <= input(7);
output(0, 59) <= input(8);
output(0, 60) <= input(9);
output(0, 61) <= input(10);
output(0, 62) <= input(11);
output(0, 63) <= input(12);
output(0, 64) <= input(19);
output(0, 65) <= input(18);
output(0, 66) <= input(17);
output(0, 67) <= input(16);
output(0, 68) <= input(0);
output(0, 69) <= input(1);
output(0, 70) <= input(2);
output(0, 71) <= input(3);
output(0, 72) <= input(4);
output(0, 73) <= input(5);
output(0, 74) <= input(6);
output(0, 75) <= input(7);
output(0, 76) <= input(8);
output(0, 77) <= input(9);
output(0, 78) <= input(10);
output(0, 79) <= input(11);
output(0, 80) <= input(20);
output(0, 81) <= input(21);
output(0, 82) <= input(22);
output(0, 83) <= input(23);
output(0, 84) <= input(24);
output(0, 85) <= input(25);
output(0, 86) <= input(26);
output(0, 87) <= input(27);
output(0, 88) <= input(28);
output(0, 89) <= input(29);
output(0, 90) <= input(30);
output(0, 91) <= input(31);
output(0, 92) <= input(32);
output(0, 93) <= input(33);
output(0, 94) <= input(34);
output(0, 95) <= input(35);
output(0, 96) <= input(36);
output(0, 97) <= input(20);
output(0, 98) <= input(21);
output(0, 99) <= input(22);
output(0, 100) <= input(23);
output(0, 101) <= input(24);
output(0, 102) <= input(25);
output(0, 103) <= input(26);
output(0, 104) <= input(27);
output(0, 105) <= input(28);
output(0, 106) <= input(29);
output(0, 107) <= input(30);
output(0, 108) <= input(31);
output(0, 109) <= input(32);
output(0, 110) <= input(33);
output(0, 111) <= input(34);
output(0, 112) <= input(37);
output(0, 113) <= input(36);
output(0, 114) <= input(20);
output(0, 115) <= input(21);
output(0, 116) <= input(22);
output(0, 117) <= input(23);
output(0, 118) <= input(24);
output(0, 119) <= input(25);
output(0, 120) <= input(26);
output(0, 121) <= input(27);
output(0, 122) <= input(28);
output(0, 123) <= input(29);
output(0, 124) <= input(30);
output(0, 125) <= input(31);
output(0, 126) <= input(32);
output(0, 127) <= input(33);
output(0, 128) <= input(38);
output(0, 129) <= input(37);
output(0, 130) <= input(36);
output(0, 131) <= input(20);
output(0, 132) <= input(21);
output(0, 133) <= input(22);
output(0, 134) <= input(23);
output(0, 135) <= input(24);
output(0, 136) <= input(25);
output(0, 137) <= input(26);
output(0, 138) <= input(27);
output(0, 139) <= input(28);
output(0, 140) <= input(29);
output(0, 141) <= input(30);
output(0, 142) <= input(31);
output(0, 143) <= input(32);
output(0, 144) <= input(39);
output(0, 145) <= input(38);
output(0, 146) <= input(37);
output(0, 147) <= input(36);
output(0, 148) <= input(20);
output(0, 149) <= input(21);
output(0, 150) <= input(22);
output(0, 151) <= input(23);
output(0, 152) <= input(24);
output(0, 153) <= input(25);
output(0, 154) <= input(26);
output(0, 155) <= input(27);
output(0, 156) <= input(28);
output(0, 157) <= input(29);
output(0, 158) <= input(30);
output(0, 159) <= input(31);
output(0, 160) <= input(40);
output(0, 161) <= input(41);
output(0, 162) <= input(42);
output(0, 163) <= input(43);
output(0, 164) <= input(44);
output(0, 165) <= input(19);
output(0, 166) <= input(18);
output(0, 167) <= input(17);
output(0, 168) <= input(16);
output(0, 169) <= input(0);
output(0, 170) <= input(1);
output(0, 171) <= input(2);
output(0, 172) <= input(3);
output(0, 173) <= input(4);
output(0, 174) <= input(5);
output(0, 175) <= input(6);
output(0, 176) <= input(45);
output(0, 177) <= input(40);
output(0, 178) <= input(41);
output(0, 179) <= input(42);
output(0, 180) <= input(43);
output(0, 181) <= input(44);
output(0, 182) <= input(19);
output(0, 183) <= input(18);
output(0, 184) <= input(17);
output(0, 185) <= input(16);
output(0, 186) <= input(0);
output(0, 187) <= input(1);
output(0, 188) <= input(2);
output(0, 189) <= input(3);
output(0, 190) <= input(4);
output(0, 191) <= input(5);
output(0, 192) <= input(46);
output(0, 193) <= input(45);
output(0, 194) <= input(40);
output(0, 195) <= input(41);
output(0, 196) <= input(42);
output(0, 197) <= input(43);
output(0, 198) <= input(44);
output(0, 199) <= input(19);
output(0, 200) <= input(18);
output(0, 201) <= input(17);
output(0, 202) <= input(16);
output(0, 203) <= input(0);
output(0, 204) <= input(1);
output(0, 205) <= input(2);
output(0, 206) <= input(3);
output(0, 207) <= input(4);
output(0, 208) <= input(47);
output(0, 209) <= input(46);
output(0, 210) <= input(45);
output(0, 211) <= input(40);
output(0, 212) <= input(41);
output(0, 213) <= input(42);
output(0, 214) <= input(43);
output(0, 215) <= input(44);
output(0, 216) <= input(19);
output(0, 217) <= input(18);
output(0, 218) <= input(17);
output(0, 219) <= input(16);
output(0, 220) <= input(0);
output(0, 221) <= input(1);
output(0, 222) <= input(2);
output(0, 223) <= input(3);
output(0, 224) <= input(48);
output(0, 225) <= input(47);
output(0, 226) <= input(46);
output(0, 227) <= input(45);
output(0, 228) <= input(40);
output(0, 229) <= input(41);
output(0, 230) <= input(42);
output(0, 231) <= input(43);
output(0, 232) <= input(44);
output(0, 233) <= input(19);
output(0, 234) <= input(18);
output(0, 235) <= input(17);
output(0, 236) <= input(16);
output(0, 237) <= input(0);
output(0, 238) <= input(1);
output(0, 239) <= input(2);
output(0, 240) <= input(49);
output(0, 241) <= input(50);
output(0, 242) <= input(51);
output(0, 243) <= input(52);
output(0, 244) <= input(53);
output(0, 245) <= input(39);
output(0, 246) <= input(38);
output(0, 247) <= input(37);
output(0, 248) <= input(36);
output(0, 249) <= input(20);
output(0, 250) <= input(21);
output(0, 251) <= input(22);
output(0, 252) <= input(23);
output(0, 253) <= input(24);
output(0, 254) <= input(25);
output(0, 255) <= input(26);
output(1, 0) <= input(54);
output(1, 1) <= input(55);
output(1, 2) <= input(56);
output(1, 3) <= input(57);
output(1, 4) <= input(58);
output(1, 5) <= input(59);
output(1, 6) <= input(60);
output(1, 7) <= input(61);
output(1, 8) <= input(62);
output(1, 9) <= input(63);
output(1, 10) <= input(64);
output(1, 11) <= input(65);
output(1, 12) <= input(66);
output(1, 13) <= input(67);
output(1, 14) <= input(68);
output(1, 15) <= input(69);
output(1, 16) <= input(70);
output(1, 17) <= input(54);
output(1, 18) <= input(55);
output(1, 19) <= input(56);
output(1, 20) <= input(57);
output(1, 21) <= input(58);
output(1, 22) <= input(59);
output(1, 23) <= input(60);
output(1, 24) <= input(61);
output(1, 25) <= input(62);
output(1, 26) <= input(63);
output(1, 27) <= input(64);
output(1, 28) <= input(65);
output(1, 29) <= input(66);
output(1, 30) <= input(67);
output(1, 31) <= input(68);
output(1, 32) <= input(71);
output(1, 33) <= input(70);
output(1, 34) <= input(54);
output(1, 35) <= input(55);
output(1, 36) <= input(56);
output(1, 37) <= input(57);
output(1, 38) <= input(58);
output(1, 39) <= input(59);
output(1, 40) <= input(60);
output(1, 41) <= input(61);
output(1, 42) <= input(62);
output(1, 43) <= input(63);
output(1, 44) <= input(64);
output(1, 45) <= input(65);
output(1, 46) <= input(66);
output(1, 47) <= input(67);
output(1, 48) <= input(72);
output(1, 49) <= input(71);
output(1, 50) <= input(70);
output(1, 51) <= input(54);
output(1, 52) <= input(55);
output(1, 53) <= input(56);
output(1, 54) <= input(57);
output(1, 55) <= input(58);
output(1, 56) <= input(59);
output(1, 57) <= input(60);
output(1, 58) <= input(61);
output(1, 59) <= input(62);
output(1, 60) <= input(63);
output(1, 61) <= input(64);
output(1, 62) <= input(65);
output(1, 63) <= input(66);
output(1, 64) <= input(73);
output(1, 65) <= input(72);
output(1, 66) <= input(71);
output(1, 67) <= input(70);
output(1, 68) <= input(54);
output(1, 69) <= input(55);
output(1, 70) <= input(56);
output(1, 71) <= input(57);
output(1, 72) <= input(58);
output(1, 73) <= input(59);
output(1, 74) <= input(60);
output(1, 75) <= input(61);
output(1, 76) <= input(62);
output(1, 77) <= input(63);
output(1, 78) <= input(64);
output(1, 79) <= input(65);
output(1, 80) <= input(74);
output(1, 81) <= input(73);
output(1, 82) <= input(72);
output(1, 83) <= input(71);
output(1, 84) <= input(70);
output(1, 85) <= input(54);
output(1, 86) <= input(55);
output(1, 87) <= input(56);
output(1, 88) <= input(57);
output(1, 89) <= input(58);
output(1, 90) <= input(59);
output(1, 91) <= input(60);
output(1, 92) <= input(61);
output(1, 93) <= input(62);
output(1, 94) <= input(63);
output(1, 95) <= input(64);
output(1, 96) <= input(75);
output(1, 97) <= input(74);
output(1, 98) <= input(73);
output(1, 99) <= input(72);
output(1, 100) <= input(71);
output(1, 101) <= input(70);
output(1, 102) <= input(54);
output(1, 103) <= input(55);
output(1, 104) <= input(56);
output(1, 105) <= input(57);
output(1, 106) <= input(58);
output(1, 107) <= input(59);
output(1, 108) <= input(60);
output(1, 109) <= input(61);
output(1, 110) <= input(62);
output(1, 111) <= input(63);
output(1, 112) <= input(76);
output(1, 113) <= input(75);
output(1, 114) <= input(74);
output(1, 115) <= input(73);
output(1, 116) <= input(72);
output(1, 117) <= input(71);
output(1, 118) <= input(70);
output(1, 119) <= input(54);
output(1, 120) <= input(55);
output(1, 121) <= input(56);
output(1, 122) <= input(57);
output(1, 123) <= input(58);
output(1, 124) <= input(59);
output(1, 125) <= input(60);
output(1, 126) <= input(61);
output(1, 127) <= input(62);
output(1, 128) <= input(77);
output(1, 129) <= input(76);
output(1, 130) <= input(75);
output(1, 131) <= input(74);
output(1, 132) <= input(73);
output(1, 133) <= input(72);
output(1, 134) <= input(71);
output(1, 135) <= input(70);
output(1, 136) <= input(54);
output(1, 137) <= input(55);
output(1, 138) <= input(56);
output(1, 139) <= input(57);
output(1, 140) <= input(58);
output(1, 141) <= input(59);
output(1, 142) <= input(60);
output(1, 143) <= input(61);
output(1, 144) <= input(78);
output(1, 145) <= input(77);
output(1, 146) <= input(76);
output(1, 147) <= input(75);
output(1, 148) <= input(74);
output(1, 149) <= input(73);
output(1, 150) <= input(72);
output(1, 151) <= input(71);
output(1, 152) <= input(70);
output(1, 153) <= input(54);
output(1, 154) <= input(55);
output(1, 155) <= input(56);
output(1, 156) <= input(57);
output(1, 157) <= input(58);
output(1, 158) <= input(59);
output(1, 159) <= input(60);
output(1, 160) <= input(79);
output(1, 161) <= input(78);
output(1, 162) <= input(77);
output(1, 163) <= input(76);
output(1, 164) <= input(75);
output(1, 165) <= input(74);
output(1, 166) <= input(73);
output(1, 167) <= input(72);
output(1, 168) <= input(71);
output(1, 169) <= input(70);
output(1, 170) <= input(54);
output(1, 171) <= input(55);
output(1, 172) <= input(56);
output(1, 173) <= input(57);
output(1, 174) <= input(58);
output(1, 175) <= input(59);
output(1, 176) <= input(80);
output(1, 177) <= input(79);
output(1, 178) <= input(78);
output(1, 179) <= input(77);
output(1, 180) <= input(76);
output(1, 181) <= input(75);
output(1, 182) <= input(74);
output(1, 183) <= input(73);
output(1, 184) <= input(72);
output(1, 185) <= input(71);
output(1, 186) <= input(70);
output(1, 187) <= input(54);
output(1, 188) <= input(55);
output(1, 189) <= input(56);
output(1, 190) <= input(57);
output(1, 191) <= input(58);
output(1, 192) <= input(81);
output(1, 193) <= input(80);
output(1, 194) <= input(79);
output(1, 195) <= input(78);
output(1, 196) <= input(77);
output(1, 197) <= input(76);
output(1, 198) <= input(75);
output(1, 199) <= input(74);
output(1, 200) <= input(73);
output(1, 201) <= input(72);
output(1, 202) <= input(71);
output(1, 203) <= input(70);
output(1, 204) <= input(54);
output(1, 205) <= input(55);
output(1, 206) <= input(56);
output(1, 207) <= input(57);
output(1, 208) <= input(82);
output(1, 209) <= input(81);
output(1, 210) <= input(80);
output(1, 211) <= input(79);
output(1, 212) <= input(78);
output(1, 213) <= input(77);
output(1, 214) <= input(76);
output(1, 215) <= input(75);
output(1, 216) <= input(74);
output(1, 217) <= input(73);
output(1, 218) <= input(72);
output(1, 219) <= input(71);
output(1, 220) <= input(70);
output(1, 221) <= input(54);
output(1, 222) <= input(55);
output(1, 223) <= input(56);
output(1, 224) <= input(83);
output(1, 225) <= input(82);
output(1, 226) <= input(81);
output(1, 227) <= input(80);
output(1, 228) <= input(79);
output(1, 229) <= input(78);
output(1, 230) <= input(77);
output(1, 231) <= input(76);
output(1, 232) <= input(75);
output(1, 233) <= input(74);
output(1, 234) <= input(73);
output(1, 235) <= input(72);
output(1, 236) <= input(71);
output(1, 237) <= input(70);
output(1, 238) <= input(54);
output(1, 239) <= input(55);
output(1, 240) <= input(84);
output(1, 241) <= input(83);
output(1, 242) <= input(82);
output(1, 243) <= input(81);
output(1, 244) <= input(80);
output(1, 245) <= input(79);
output(1, 246) <= input(78);
output(1, 247) <= input(77);
output(1, 248) <= input(76);
output(1, 249) <= input(75);
output(1, 250) <= input(74);
output(1, 251) <= input(73);
output(1, 252) <= input(72);
output(1, 253) <= input(71);
output(1, 254) <= input(70);
output(1, 255) <= input(54);
when "1000" =>
output(0, 0) <= input(0);
output(0, 1) <= input(1);
output(0, 2) <= input(2);
output(0, 3) <= input(3);
output(0, 4) <= input(4);
output(0, 5) <= input(5);
output(0, 6) <= input(6);
output(0, 7) <= input(7);
output(0, 8) <= input(8);
output(0, 9) <= input(9);
output(0, 10) <= input(10);
output(0, 11) <= input(11);
output(0, 12) <= input(12);
output(0, 13) <= input(13);
output(0, 14) <= input(14);
output(0, 15) <= input(15);
output(0, 16) <= input(16);
output(0, 17) <= input(0);
output(0, 18) <= input(1);
output(0, 19) <= input(2);
output(0, 20) <= input(3);
output(0, 21) <= input(4);
output(0, 22) <= input(5);
output(0, 23) <= input(6);
output(0, 24) <= input(7);
output(0, 25) <= input(8);
output(0, 26) <= input(9);
output(0, 27) <= input(10);
output(0, 28) <= input(11);
output(0, 29) <= input(12);
output(0, 30) <= input(13);
output(0, 31) <= input(14);
output(0, 32) <= input(17);
output(0, 33) <= input(16);
output(0, 34) <= input(0);
output(0, 35) <= input(1);
output(0, 36) <= input(2);
output(0, 37) <= input(3);
output(0, 38) <= input(4);
output(0, 39) <= input(5);
output(0, 40) <= input(6);
output(0, 41) <= input(7);
output(0, 42) <= input(8);
output(0, 43) <= input(9);
output(0, 44) <= input(10);
output(0, 45) <= input(11);
output(0, 46) <= input(12);
output(0, 47) <= input(13);
output(0, 48) <= input(18);
output(0, 49) <= input(17);
output(0, 50) <= input(16);
output(0, 51) <= input(0);
output(0, 52) <= input(1);
output(0, 53) <= input(2);
output(0, 54) <= input(3);
output(0, 55) <= input(4);
output(0, 56) <= input(5);
output(0, 57) <= input(6);
output(0, 58) <= input(7);
output(0, 59) <= input(8);
output(0, 60) <= input(9);
output(0, 61) <= input(10);
output(0, 62) <= input(11);
output(0, 63) <= input(12);
output(0, 64) <= input(19);
output(0, 65) <= input(18);
output(0, 66) <= input(17);
output(0, 67) <= input(16);
output(0, 68) <= input(0);
output(0, 69) <= input(1);
output(0, 70) <= input(2);
output(0, 71) <= input(3);
output(0, 72) <= input(4);
output(0, 73) <= input(5);
output(0, 74) <= input(6);
output(0, 75) <= input(7);
output(0, 76) <= input(8);
output(0, 77) <= input(9);
output(0, 78) <= input(10);
output(0, 79) <= input(11);
output(0, 80) <= input(20);
output(0, 81) <= input(21);
output(0, 82) <= input(22);
output(0, 83) <= input(23);
output(0, 84) <= input(24);
output(0, 85) <= input(25);
output(0, 86) <= input(26);
output(0, 87) <= input(27);
output(0, 88) <= input(28);
output(0, 89) <= input(29);
output(0, 90) <= input(30);
output(0, 91) <= input(31);
output(0, 92) <= input(32);
output(0, 93) <= input(33);
output(0, 94) <= input(34);
output(0, 95) <= input(35);
output(0, 96) <= input(36);
output(0, 97) <= input(20);
output(0, 98) <= input(21);
output(0, 99) <= input(22);
output(0, 100) <= input(23);
output(0, 101) <= input(24);
output(0, 102) <= input(25);
output(0, 103) <= input(26);
output(0, 104) <= input(27);
output(0, 105) <= input(28);
output(0, 106) <= input(29);
output(0, 107) <= input(30);
output(0, 108) <= input(31);
output(0, 109) <= input(32);
output(0, 110) <= input(33);
output(0, 111) <= input(34);
output(0, 112) <= input(37);
output(0, 113) <= input(36);
output(0, 114) <= input(20);
output(0, 115) <= input(21);
output(0, 116) <= input(22);
output(0, 117) <= input(23);
output(0, 118) <= input(24);
output(0, 119) <= input(25);
output(0, 120) <= input(26);
output(0, 121) <= input(27);
output(0, 122) <= input(28);
output(0, 123) <= input(29);
output(0, 124) <= input(30);
output(0, 125) <= input(31);
output(0, 126) <= input(32);
output(0, 127) <= input(33);
output(0, 128) <= input(38);
output(0, 129) <= input(37);
output(0, 130) <= input(36);
output(0, 131) <= input(20);
output(0, 132) <= input(21);
output(0, 133) <= input(22);
output(0, 134) <= input(23);
output(0, 135) <= input(24);
output(0, 136) <= input(25);
output(0, 137) <= input(26);
output(0, 138) <= input(27);
output(0, 139) <= input(28);
output(0, 140) <= input(29);
output(0, 141) <= input(30);
output(0, 142) <= input(31);
output(0, 143) <= input(32);
output(0, 144) <= input(39);
output(0, 145) <= input(38);
output(0, 146) <= input(37);
output(0, 147) <= input(36);
output(0, 148) <= input(20);
output(0, 149) <= input(21);
output(0, 150) <= input(22);
output(0, 151) <= input(23);
output(0, 152) <= input(24);
output(0, 153) <= input(25);
output(0, 154) <= input(26);
output(0, 155) <= input(27);
output(0, 156) <= input(28);
output(0, 157) <= input(29);
output(0, 158) <= input(30);
output(0, 159) <= input(31);
output(0, 160) <= input(40);
output(0, 161) <= input(41);
output(0, 162) <= input(42);
output(0, 163) <= input(43);
output(0, 164) <= input(44);
output(0, 165) <= input(19);
output(0, 166) <= input(18);
output(0, 167) <= input(17);
output(0, 168) <= input(16);
output(0, 169) <= input(0);
output(0, 170) <= input(1);
output(0, 171) <= input(2);
output(0, 172) <= input(3);
output(0, 173) <= input(4);
output(0, 174) <= input(5);
output(0, 175) <= input(6);
output(0, 176) <= input(45);
output(0, 177) <= input(40);
output(0, 178) <= input(41);
output(0, 179) <= input(42);
output(0, 180) <= input(43);
output(0, 181) <= input(44);
output(0, 182) <= input(19);
output(0, 183) <= input(18);
output(0, 184) <= input(17);
output(0, 185) <= input(16);
output(0, 186) <= input(0);
output(0, 187) <= input(1);
output(0, 188) <= input(2);
output(0, 189) <= input(3);
output(0, 190) <= input(4);
output(0, 191) <= input(5);
output(0, 192) <= input(46);
output(0, 193) <= input(45);
output(0, 194) <= input(40);
output(0, 195) <= input(41);
output(0, 196) <= input(42);
output(0, 197) <= input(43);
output(0, 198) <= input(44);
output(0, 199) <= input(19);
output(0, 200) <= input(18);
output(0, 201) <= input(17);
output(0, 202) <= input(16);
output(0, 203) <= input(0);
output(0, 204) <= input(1);
output(0, 205) <= input(2);
output(0, 206) <= input(3);
output(0, 207) <= input(4);
output(0, 208) <= input(47);
output(0, 209) <= input(46);
output(0, 210) <= input(45);
output(0, 211) <= input(40);
output(0, 212) <= input(41);
output(0, 213) <= input(42);
output(0, 214) <= input(43);
output(0, 215) <= input(44);
output(0, 216) <= input(19);
output(0, 217) <= input(18);
output(0, 218) <= input(17);
output(0, 219) <= input(16);
output(0, 220) <= input(0);
output(0, 221) <= input(1);
output(0, 222) <= input(2);
output(0, 223) <= input(3);
output(0, 224) <= input(48);
output(0, 225) <= input(47);
output(0, 226) <= input(46);
output(0, 227) <= input(45);
output(0, 228) <= input(40);
output(0, 229) <= input(41);
output(0, 230) <= input(42);
output(0, 231) <= input(43);
output(0, 232) <= input(44);
output(0, 233) <= input(19);
output(0, 234) <= input(18);
output(0, 235) <= input(17);
output(0, 236) <= input(16);
output(0, 237) <= input(0);
output(0, 238) <= input(1);
output(0, 239) <= input(2);
output(0, 240) <= input(49);
output(0, 241) <= input(50);
output(0, 242) <= input(51);
output(0, 243) <= input(52);
output(0, 244) <= input(53);
output(0, 245) <= input(39);
output(0, 246) <= input(38);
output(0, 247) <= input(37);
output(0, 248) <= input(36);
output(0, 249) <= input(20);
output(0, 250) <= input(21);
output(0, 251) <= input(22);
output(0, 252) <= input(23);
output(0, 253) <= input(24);
output(0, 254) <= input(25);
output(0, 255) <= input(26);
when "1001" =>
output(0, 0) <= input(0);
output(0, 1) <= input(1);
output(0, 2) <= input(2);
output(0, 3) <= input(3);
output(0, 4) <= input(4);
output(0, 5) <= input(5);
output(0, 6) <= input(6);
output(0, 7) <= input(7);
output(0, 8) <= input(8);
output(0, 9) <= input(9);
output(0, 10) <= input(10);
output(0, 11) <= input(11);
output(0, 12) <= input(12);
output(0, 13) <= input(13);
output(0, 14) <= input(14);
output(0, 15) <= input(15);
output(0, 16) <= input(16);
output(0, 17) <= input(0);
output(0, 18) <= input(1);
output(0, 19) <= input(2);
output(0, 20) <= input(3);
output(0, 21) <= input(4);
output(0, 22) <= input(5);
output(0, 23) <= input(6);
output(0, 24) <= input(7);
output(0, 25) <= input(8);
output(0, 26) <= input(9);
output(0, 27) <= input(10);
output(0, 28) <= input(11);
output(0, 29) <= input(12);
output(0, 30) <= input(13);
output(0, 31) <= input(14);
output(0, 32) <= input(17);
output(0, 33) <= input(18);
output(0, 34) <= input(19);
output(0, 35) <= input(20);
output(0, 36) <= input(21);
output(0, 37) <= input(22);
output(0, 38) <= input(23);
output(0, 39) <= input(24);
output(0, 40) <= input(25);
output(0, 41) <= input(26);
output(0, 42) <= input(27);
output(0, 43) <= input(28);
output(0, 44) <= input(29);
output(0, 45) <= input(30);
output(0, 46) <= input(31);
output(0, 47) <= input(32);
output(0, 48) <= input(33);
output(0, 49) <= input(17);
output(0, 50) <= input(18);
output(0, 51) <= input(19);
output(0, 52) <= input(20);
output(0, 53) <= input(21);
output(0, 54) <= input(22);
output(0, 55) <= input(23);
output(0, 56) <= input(24);
output(0, 57) <= input(25);
output(0, 58) <= input(26);
output(0, 59) <= input(27);
output(0, 60) <= input(28);
output(0, 61) <= input(29);
output(0, 62) <= input(30);
output(0, 63) <= input(31);
output(0, 64) <= input(34);
output(0, 65) <= input(33);
output(0, 66) <= input(17);
output(0, 67) <= input(18);
output(0, 68) <= input(19);
output(0, 69) <= input(20);
output(0, 70) <= input(21);
output(0, 71) <= input(22);
output(0, 72) <= input(23);
output(0, 73) <= input(24);
output(0, 74) <= input(25);
output(0, 75) <= input(26);
output(0, 76) <= input(27);
output(0, 77) <= input(28);
output(0, 78) <= input(29);
output(0, 79) <= input(30);
output(0, 80) <= input(35);
output(0, 81) <= input(36);
output(0, 82) <= input(37);
output(0, 83) <= input(16);
output(0, 84) <= input(0);
output(0, 85) <= input(1);
output(0, 86) <= input(2);
output(0, 87) <= input(3);
output(0, 88) <= input(4);
output(0, 89) <= input(5);
output(0, 90) <= input(6);
output(0, 91) <= input(7);
output(0, 92) <= input(8);
output(0, 93) <= input(9);
output(0, 94) <= input(10);
output(0, 95) <= input(11);
output(0, 96) <= input(38);
output(0, 97) <= input(35);
output(0, 98) <= input(36);
output(0, 99) <= input(37);
output(0, 100) <= input(16);
output(0, 101) <= input(0);
output(0, 102) <= input(1);
output(0, 103) <= input(2);
output(0, 104) <= input(3);
output(0, 105) <= input(4);
output(0, 106) <= input(5);
output(0, 107) <= input(6);
output(0, 108) <= input(7);
output(0, 109) <= input(8);
output(0, 110) <= input(9);
output(0, 111) <= input(10);
output(0, 112) <= input(39);
output(0, 113) <= input(40);
output(0, 114) <= input(34);
output(0, 115) <= input(33);
output(0, 116) <= input(17);
output(0, 117) <= input(18);
output(0, 118) <= input(19);
output(0, 119) <= input(20);
output(0, 120) <= input(21);
output(0, 121) <= input(22);
output(0, 122) <= input(23);
output(0, 123) <= input(24);
output(0, 124) <= input(25);
output(0, 125) <= input(26);
output(0, 126) <= input(27);
output(0, 127) <= input(28);
output(0, 128) <= input(41);
output(0, 129) <= input(39);
output(0, 130) <= input(40);
output(0, 131) <= input(34);
output(0, 132) <= input(33);
output(0, 133) <= input(17);
output(0, 134) <= input(18);
output(0, 135) <= input(19);
output(0, 136) <= input(20);
output(0, 137) <= input(21);
output(0, 138) <= input(22);
output(0, 139) <= input(23);
output(0, 140) <= input(24);
output(0, 141) <= input(25);
output(0, 142) <= input(26);
output(0, 143) <= input(27);
output(0, 144) <= input(42);
output(0, 145) <= input(41);
output(0, 146) <= input(39);
output(0, 147) <= input(40);
output(0, 148) <= input(34);
output(0, 149) <= input(33);
output(0, 150) <= input(17);
output(0, 151) <= input(18);
output(0, 152) <= input(19);
output(0, 153) <= input(20);
output(0, 154) <= input(21);
output(0, 155) <= input(22);
output(0, 156) <= input(23);
output(0, 157) <= input(24);
output(0, 158) <= input(25);
output(0, 159) <= input(26);
output(0, 160) <= input(43);
output(0, 161) <= input(44);
output(0, 162) <= input(45);
output(0, 163) <= input(38);
output(0, 164) <= input(35);
output(0, 165) <= input(36);
output(0, 166) <= input(37);
output(0, 167) <= input(16);
output(0, 168) <= input(0);
output(0, 169) <= input(1);
output(0, 170) <= input(2);
output(0, 171) <= input(3);
output(0, 172) <= input(4);
output(0, 173) <= input(5);
output(0, 174) <= input(6);
output(0, 175) <= input(7);
output(0, 176) <= input(46);
output(0, 177) <= input(43);
output(0, 178) <= input(44);
output(0, 179) <= input(45);
output(0, 180) <= input(38);
output(0, 181) <= input(35);
output(0, 182) <= input(36);
output(0, 183) <= input(37);
output(0, 184) <= input(16);
output(0, 185) <= input(0);
output(0, 186) <= input(1);
output(0, 187) <= input(2);
output(0, 188) <= input(3);
output(0, 189) <= input(4);
output(0, 190) <= input(5);
output(0, 191) <= input(6);
output(0, 192) <= input(47);
output(0, 193) <= input(46);
output(0, 194) <= input(43);
output(0, 195) <= input(44);
output(0, 196) <= input(45);
output(0, 197) <= input(38);
output(0, 198) <= input(35);
output(0, 199) <= input(36);
output(0, 200) <= input(37);
output(0, 201) <= input(16);
output(0, 202) <= input(0);
output(0, 203) <= input(1);
output(0, 204) <= input(2);
output(0, 205) <= input(3);
output(0, 206) <= input(4);
output(0, 207) <= input(5);
output(0, 208) <= input(48);
output(0, 209) <= input(49);
output(0, 210) <= input(50);
output(0, 211) <= input(42);
output(0, 212) <= input(41);
output(0, 213) <= input(39);
output(0, 214) <= input(40);
output(0, 215) <= input(34);
output(0, 216) <= input(33);
output(0, 217) <= input(17);
output(0, 218) <= input(18);
output(0, 219) <= input(19);
output(0, 220) <= input(20);
output(0, 221) <= input(21);
output(0, 222) <= input(22);
output(0, 223) <= input(23);
output(0, 224) <= input(51);
output(0, 225) <= input(48);
output(0, 226) <= input(49);
output(0, 227) <= input(50);
output(0, 228) <= input(42);
output(0, 229) <= input(41);
output(0, 230) <= input(39);
output(0, 231) <= input(40);
output(0, 232) <= input(34);
output(0, 233) <= input(33);
output(0, 234) <= input(17);
output(0, 235) <= input(18);
output(0, 236) <= input(19);
output(0, 237) <= input(20);
output(0, 238) <= input(21);
output(0, 239) <= input(22);
output(0, 240) <= input(52);
output(0, 241) <= input(53);
output(0, 242) <= input(47);
output(0, 243) <= input(46);
output(0, 244) <= input(43);
output(0, 245) <= input(44);
output(0, 246) <= input(45);
output(0, 247) <= input(38);
output(0, 248) <= input(35);
output(0, 249) <= input(36);
output(0, 250) <= input(37);
output(0, 251) <= input(16);
output(0, 252) <= input(0);
output(0, 253) <= input(1);
output(0, 254) <= input(2);
output(0, 255) <= input(3);
output(1, 0) <= input(20);
output(1, 1) <= input(21);
output(1, 2) <= input(22);
output(1, 3) <= input(23);
output(1, 4) <= input(24);
output(1, 5) <= input(25);
output(1, 6) <= input(26);
output(1, 7) <= input(27);
output(1, 8) <= input(28);
output(1, 9) <= input(29);
output(1, 10) <= input(30);
output(1, 11) <= input(31);
output(1, 12) <= input(32);
output(1, 13) <= input(54);
output(1, 14) <= input(55);
output(1, 15) <= input(56);
output(1, 16) <= input(1);
output(1, 17) <= input(2);
output(1, 18) <= input(3);
output(1, 19) <= input(4);
output(1, 20) <= input(5);
output(1, 21) <= input(6);
output(1, 22) <= input(7);
output(1, 23) <= input(8);
output(1, 24) <= input(9);
output(1, 25) <= input(10);
output(1, 26) <= input(11);
output(1, 27) <= input(12);
output(1, 28) <= input(13);
output(1, 29) <= input(14);
output(1, 30) <= input(15);
output(1, 31) <= input(57);
output(1, 32) <= input(0);
output(1, 33) <= input(1);
output(1, 34) <= input(2);
output(1, 35) <= input(3);
output(1, 36) <= input(4);
output(1, 37) <= input(5);
output(1, 38) <= input(6);
output(1, 39) <= input(7);
output(1, 40) <= input(8);
output(1, 41) <= input(9);
output(1, 42) <= input(10);
output(1, 43) <= input(11);
output(1, 44) <= input(12);
output(1, 45) <= input(13);
output(1, 46) <= input(14);
output(1, 47) <= input(15);
output(1, 48) <= input(18);
output(1, 49) <= input(19);
output(1, 50) <= input(20);
output(1, 51) <= input(21);
output(1, 52) <= input(22);
output(1, 53) <= input(23);
output(1, 54) <= input(24);
output(1, 55) <= input(25);
output(1, 56) <= input(26);
output(1, 57) <= input(27);
output(1, 58) <= input(28);
output(1, 59) <= input(29);
output(1, 60) <= input(30);
output(1, 61) <= input(31);
output(1, 62) <= input(32);
output(1, 63) <= input(54);
output(1, 64) <= input(17);
output(1, 65) <= input(18);
output(1, 66) <= input(19);
output(1, 67) <= input(20);
output(1, 68) <= input(21);
output(1, 69) <= input(22);
output(1, 70) <= input(23);
output(1, 71) <= input(24);
output(1, 72) <= input(25);
output(1, 73) <= input(26);
output(1, 74) <= input(27);
output(1, 75) <= input(28);
output(1, 76) <= input(29);
output(1, 77) <= input(30);
output(1, 78) <= input(31);
output(1, 79) <= input(32);
output(1, 80) <= input(37);
output(1, 81) <= input(16);
output(1, 82) <= input(0);
output(1, 83) <= input(1);
output(1, 84) <= input(2);
output(1, 85) <= input(3);
output(1, 86) <= input(4);
output(1, 87) <= input(5);
output(1, 88) <= input(6);
output(1, 89) <= input(7);
output(1, 90) <= input(8);
output(1, 91) <= input(9);
output(1, 92) <= input(10);
output(1, 93) <= input(11);
output(1, 94) <= input(12);
output(1, 95) <= input(13);
output(1, 96) <= input(36);
output(1, 97) <= input(37);
output(1, 98) <= input(16);
output(1, 99) <= input(0);
output(1, 100) <= input(1);
output(1, 101) <= input(2);
output(1, 102) <= input(3);
output(1, 103) <= input(4);
output(1, 104) <= input(5);
output(1, 105) <= input(6);
output(1, 106) <= input(7);
output(1, 107) <= input(8);
output(1, 108) <= input(9);
output(1, 109) <= input(10);
output(1, 110) <= input(11);
output(1, 111) <= input(12);
output(1, 112) <= input(34);
output(1, 113) <= input(33);
output(1, 114) <= input(17);
output(1, 115) <= input(18);
output(1, 116) <= input(19);
output(1, 117) <= input(20);
output(1, 118) <= input(21);
output(1, 119) <= input(22);
output(1, 120) <= input(23);
output(1, 121) <= input(24);
output(1, 122) <= input(25);
output(1, 123) <= input(26);
output(1, 124) <= input(27);
output(1, 125) <= input(28);
output(1, 126) <= input(29);
output(1, 127) <= input(30);
output(1, 128) <= input(35);
output(1, 129) <= input(36);
output(1, 130) <= input(37);
output(1, 131) <= input(16);
output(1, 132) <= input(0);
output(1, 133) <= input(1);
output(1, 134) <= input(2);
output(1, 135) <= input(3);
output(1, 136) <= input(4);
output(1, 137) <= input(5);
output(1, 138) <= input(6);
output(1, 139) <= input(7);
output(1, 140) <= input(8);
output(1, 141) <= input(9);
output(1, 142) <= input(10);
output(1, 143) <= input(11);
output(1, 144) <= input(38);
output(1, 145) <= input(35);
output(1, 146) <= input(36);
output(1, 147) <= input(37);
output(1, 148) <= input(16);
output(1, 149) <= input(0);
output(1, 150) <= input(1);
output(1, 151) <= input(2);
output(1, 152) <= input(3);
output(1, 153) <= input(4);
output(1, 154) <= input(5);
output(1, 155) <= input(6);
output(1, 156) <= input(7);
output(1, 157) <= input(8);
output(1, 158) <= input(9);
output(1, 159) <= input(10);
output(1, 160) <= input(39);
output(1, 161) <= input(40);
output(1, 162) <= input(34);
output(1, 163) <= input(33);
output(1, 164) <= input(17);
output(1, 165) <= input(18);
output(1, 166) <= input(19);
output(1, 167) <= input(20);
output(1, 168) <= input(21);
output(1, 169) <= input(22);
output(1, 170) <= input(23);
output(1, 171) <= input(24);
output(1, 172) <= input(25);
output(1, 173) <= input(26);
output(1, 174) <= input(27);
output(1, 175) <= input(28);
output(1, 176) <= input(41);
output(1, 177) <= input(39);
output(1, 178) <= input(40);
output(1, 179) <= input(34);
output(1, 180) <= input(33);
output(1, 181) <= input(17);
output(1, 182) <= input(18);
output(1, 183) <= input(19);
output(1, 184) <= input(20);
output(1, 185) <= input(21);
output(1, 186) <= input(22);
output(1, 187) <= input(23);
output(1, 188) <= input(24);
output(1, 189) <= input(25);
output(1, 190) <= input(26);
output(1, 191) <= input(27);
output(1, 192) <= input(44);
output(1, 193) <= input(45);
output(1, 194) <= input(38);
output(1, 195) <= input(35);
output(1, 196) <= input(36);
output(1, 197) <= input(37);
output(1, 198) <= input(16);
output(1, 199) <= input(0);
output(1, 200) <= input(1);
output(1, 201) <= input(2);
output(1, 202) <= input(3);
output(1, 203) <= input(4);
output(1, 204) <= input(5);
output(1, 205) <= input(6);
output(1, 206) <= input(7);
output(1, 207) <= input(8);
output(1, 208) <= input(43);
output(1, 209) <= input(44);
output(1, 210) <= input(45);
output(1, 211) <= input(38);
output(1, 212) <= input(35);
output(1, 213) <= input(36);
output(1, 214) <= input(37);
output(1, 215) <= input(16);
output(1, 216) <= input(0);
output(1, 217) <= input(1);
output(1, 218) <= input(2);
output(1, 219) <= input(3);
output(1, 220) <= input(4);
output(1, 221) <= input(5);
output(1, 222) <= input(6);
output(1, 223) <= input(7);
output(1, 224) <= input(50);
output(1, 225) <= input(42);
output(1, 226) <= input(41);
output(1, 227) <= input(39);
output(1, 228) <= input(40);
output(1, 229) <= input(34);
output(1, 230) <= input(33);
output(1, 231) <= input(17);
output(1, 232) <= input(18);
output(1, 233) <= input(19);
output(1, 234) <= input(20);
output(1, 235) <= input(21);
output(1, 236) <= input(22);
output(1, 237) <= input(23);
output(1, 238) <= input(24);
output(1, 239) <= input(25);
output(1, 240) <= input(46);
output(1, 241) <= input(43);
output(1, 242) <= input(44);
output(1, 243) <= input(45);
output(1, 244) <= input(38);
output(1, 245) <= input(35);
output(1, 246) <= input(36);
output(1, 247) <= input(37);
output(1, 248) <= input(16);
output(1, 249) <= input(0);
output(1, 250) <= input(1);
output(1, 251) <= input(2);
output(1, 252) <= input(3);
output(1, 253) <= input(4);
output(1, 254) <= input(5);
output(1, 255) <= input(6);
output(2, 0) <= input(3);
output(2, 1) <= input(4);
output(2, 2) <= input(5);
output(2, 3) <= input(6);
output(2, 4) <= input(7);
output(2, 5) <= input(8);
output(2, 6) <= input(9);
output(2, 7) <= input(10);
output(2, 8) <= input(11);
output(2, 9) <= input(12);
output(2, 10) <= input(13);
output(2, 11) <= input(14);
output(2, 12) <= input(15);
output(2, 13) <= input(57);
output(2, 14) <= input(58);
output(2, 15) <= input(59);
output(2, 16) <= input(21);
output(2, 17) <= input(22);
output(2, 18) <= input(23);
output(2, 19) <= input(24);
output(2, 20) <= input(25);
output(2, 21) <= input(26);
output(2, 22) <= input(27);
output(2, 23) <= input(28);
output(2, 24) <= input(29);
output(2, 25) <= input(30);
output(2, 26) <= input(31);
output(2, 27) <= input(32);
output(2, 28) <= input(54);
output(2, 29) <= input(55);
output(2, 30) <= input(56);
output(2, 31) <= input(60);
output(2, 32) <= input(2);
output(2, 33) <= input(3);
output(2, 34) <= input(4);
output(2, 35) <= input(5);
output(2, 36) <= input(6);
output(2, 37) <= input(7);
output(2, 38) <= input(8);
output(2, 39) <= input(9);
output(2, 40) <= input(10);
output(2, 41) <= input(11);
output(2, 42) <= input(12);
output(2, 43) <= input(13);
output(2, 44) <= input(14);
output(2, 45) <= input(15);
output(2, 46) <= input(57);
output(2, 47) <= input(58);
output(2, 48) <= input(20);
output(2, 49) <= input(21);
output(2, 50) <= input(22);
output(2, 51) <= input(23);
output(2, 52) <= input(24);
output(2, 53) <= input(25);
output(2, 54) <= input(26);
output(2, 55) <= input(27);
output(2, 56) <= input(28);
output(2, 57) <= input(29);
output(2, 58) <= input(30);
output(2, 59) <= input(31);
output(2, 60) <= input(32);
output(2, 61) <= input(54);
output(2, 62) <= input(55);
output(2, 63) <= input(56);
output(2, 64) <= input(19);
output(2, 65) <= input(20);
output(2, 66) <= input(21);
output(2, 67) <= input(22);
output(2, 68) <= input(23);
output(2, 69) <= input(24);
output(2, 70) <= input(25);
output(2, 71) <= input(26);
output(2, 72) <= input(27);
output(2, 73) <= input(28);
output(2, 74) <= input(29);
output(2, 75) <= input(30);
output(2, 76) <= input(31);
output(2, 77) <= input(32);
output(2, 78) <= input(54);
output(2, 79) <= input(55);
output(2, 80) <= input(0);
output(2, 81) <= input(1);
output(2, 82) <= input(2);
output(2, 83) <= input(3);
output(2, 84) <= input(4);
output(2, 85) <= input(5);
output(2, 86) <= input(6);
output(2, 87) <= input(7);
output(2, 88) <= input(8);
output(2, 89) <= input(9);
output(2, 90) <= input(10);
output(2, 91) <= input(11);
output(2, 92) <= input(12);
output(2, 93) <= input(13);
output(2, 94) <= input(14);
output(2, 95) <= input(15);
output(2, 96) <= input(18);
output(2, 97) <= input(19);
output(2, 98) <= input(20);
output(2, 99) <= input(21);
output(2, 100) <= input(22);
output(2, 101) <= input(23);
output(2, 102) <= input(24);
output(2, 103) <= input(25);
output(2, 104) <= input(26);
output(2, 105) <= input(27);
output(2, 106) <= input(28);
output(2, 107) <= input(29);
output(2, 108) <= input(30);
output(2, 109) <= input(31);
output(2, 110) <= input(32);
output(2, 111) <= input(54);
output(2, 112) <= input(16);
output(2, 113) <= input(0);
output(2, 114) <= input(1);
output(2, 115) <= input(2);
output(2, 116) <= input(3);
output(2, 117) <= input(4);
output(2, 118) <= input(5);
output(2, 119) <= input(6);
output(2, 120) <= input(7);
output(2, 121) <= input(8);
output(2, 122) <= input(9);
output(2, 123) <= input(10);
output(2, 124) <= input(11);
output(2, 125) <= input(12);
output(2, 126) <= input(13);
output(2, 127) <= input(14);
output(2, 128) <= input(37);
output(2, 129) <= input(16);
output(2, 130) <= input(0);
output(2, 131) <= input(1);
output(2, 132) <= input(2);
output(2, 133) <= input(3);
output(2, 134) <= input(4);
output(2, 135) <= input(5);
output(2, 136) <= input(6);
output(2, 137) <= input(7);
output(2, 138) <= input(8);
output(2, 139) <= input(9);
output(2, 140) <= input(10);
output(2, 141) <= input(11);
output(2, 142) <= input(12);
output(2, 143) <= input(13);
output(2, 144) <= input(33);
output(2, 145) <= input(17);
output(2, 146) <= input(18);
output(2, 147) <= input(19);
output(2, 148) <= input(20);
output(2, 149) <= input(21);
output(2, 150) <= input(22);
output(2, 151) <= input(23);
output(2, 152) <= input(24);
output(2, 153) <= input(25);
output(2, 154) <= input(26);
output(2, 155) <= input(27);
output(2, 156) <= input(28);
output(2, 157) <= input(29);
output(2, 158) <= input(30);
output(2, 159) <= input(31);
output(2, 160) <= input(36);
output(2, 161) <= input(37);
output(2, 162) <= input(16);
output(2, 163) <= input(0);
output(2, 164) <= input(1);
output(2, 165) <= input(2);
output(2, 166) <= input(3);
output(2, 167) <= input(4);
output(2, 168) <= input(5);
output(2, 169) <= input(6);
output(2, 170) <= input(7);
output(2, 171) <= input(8);
output(2, 172) <= input(9);
output(2, 173) <= input(10);
output(2, 174) <= input(11);
output(2, 175) <= input(12);
output(2, 176) <= input(34);
output(2, 177) <= input(33);
output(2, 178) <= input(17);
output(2, 179) <= input(18);
output(2, 180) <= input(19);
output(2, 181) <= input(20);
output(2, 182) <= input(21);
output(2, 183) <= input(22);
output(2, 184) <= input(23);
output(2, 185) <= input(24);
output(2, 186) <= input(25);
output(2, 187) <= input(26);
output(2, 188) <= input(27);
output(2, 189) <= input(28);
output(2, 190) <= input(29);
output(2, 191) <= input(30);
output(2, 192) <= input(40);
output(2, 193) <= input(34);
output(2, 194) <= input(33);
output(2, 195) <= input(17);
output(2, 196) <= input(18);
output(2, 197) <= input(19);
output(2, 198) <= input(20);
output(2, 199) <= input(21);
output(2, 200) <= input(22);
output(2, 201) <= input(23);
output(2, 202) <= input(24);
output(2, 203) <= input(25);
output(2, 204) <= input(26);
output(2, 205) <= input(27);
output(2, 206) <= input(28);
output(2, 207) <= input(29);
output(2, 208) <= input(38);
output(2, 209) <= input(35);
output(2, 210) <= input(36);
output(2, 211) <= input(37);
output(2, 212) <= input(16);
output(2, 213) <= input(0);
output(2, 214) <= input(1);
output(2, 215) <= input(2);
output(2, 216) <= input(3);
output(2, 217) <= input(4);
output(2, 218) <= input(5);
output(2, 219) <= input(6);
output(2, 220) <= input(7);
output(2, 221) <= input(8);
output(2, 222) <= input(9);
output(2, 223) <= input(10);
output(2, 224) <= input(39);
output(2, 225) <= input(40);
output(2, 226) <= input(34);
output(2, 227) <= input(33);
output(2, 228) <= input(17);
output(2, 229) <= input(18);
output(2, 230) <= input(19);
output(2, 231) <= input(20);
output(2, 232) <= input(21);
output(2, 233) <= input(22);
output(2, 234) <= input(23);
output(2, 235) <= input(24);
output(2, 236) <= input(25);
output(2, 237) <= input(26);
output(2, 238) <= input(27);
output(2, 239) <= input(28);
output(2, 240) <= input(45);
output(2, 241) <= input(38);
output(2, 242) <= input(35);
output(2, 243) <= input(36);
output(2, 244) <= input(37);
output(2, 245) <= input(16);
output(2, 246) <= input(0);
output(2, 247) <= input(1);
output(2, 248) <= input(2);
output(2, 249) <= input(3);
output(2, 250) <= input(4);
output(2, 251) <= input(5);
output(2, 252) <= input(6);
output(2, 253) <= input(7);
output(2, 254) <= input(8);
output(2, 255) <= input(9);
when "1010" =>
output(0, 0) <= input(0);
output(0, 1) <= input(1);
output(0, 2) <= input(2);
output(0, 3) <= input(3);
output(0, 4) <= input(4);
output(0, 5) <= input(5);
output(0, 6) <= input(6);
output(0, 7) <= input(7);
output(0, 8) <= input(8);
output(0, 9) <= input(9);
output(0, 10) <= input(10);
output(0, 11) <= input(11);
output(0, 12) <= input(12);
output(0, 13) <= input(13);
output(0, 14) <= input(14);
output(0, 15) <= input(15);
output(0, 16) <= input(16);
output(0, 17) <= input(17);
output(0, 18) <= input(18);
output(0, 19) <= input(19);
output(0, 20) <= input(20);
output(0, 21) <= input(21);
output(0, 22) <= input(22);
output(0, 23) <= input(23);
output(0, 24) <= input(24);
output(0, 25) <= input(25);
output(0, 26) <= input(26);
output(0, 27) <= input(27);
output(0, 28) <= input(28);
output(0, 29) <= input(29);
output(0, 30) <= input(30);
output(0, 31) <= input(31);
output(0, 32) <= input(32);
output(0, 33) <= input(0);
output(0, 34) <= input(1);
output(0, 35) <= input(2);
output(0, 36) <= input(3);
output(0, 37) <= input(4);
output(0, 38) <= input(5);
output(0, 39) <= input(6);
output(0, 40) <= input(7);
output(0, 41) <= input(8);
output(0, 42) <= input(9);
output(0, 43) <= input(10);
output(0, 44) <= input(11);
output(0, 45) <= input(12);
output(0, 46) <= input(13);
output(0, 47) <= input(14);
output(0, 48) <= input(33);
output(0, 49) <= input(16);
output(0, 50) <= input(17);
output(0, 51) <= input(18);
output(0, 52) <= input(19);
output(0, 53) <= input(20);
output(0, 54) <= input(21);
output(0, 55) <= input(22);
output(0, 56) <= input(23);
output(0, 57) <= input(24);
output(0, 58) <= input(25);
output(0, 59) <= input(26);
output(0, 60) <= input(27);
output(0, 61) <= input(28);
output(0, 62) <= input(29);
output(0, 63) <= input(30);
output(0, 64) <= input(34);
output(0, 65) <= input(32);
output(0, 66) <= input(0);
output(0, 67) <= input(1);
output(0, 68) <= input(2);
output(0, 69) <= input(3);
output(0, 70) <= input(4);
output(0, 71) <= input(5);
output(0, 72) <= input(6);
output(0, 73) <= input(7);
output(0, 74) <= input(8);
output(0, 75) <= input(9);
output(0, 76) <= input(10);
output(0, 77) <= input(11);
output(0, 78) <= input(12);
output(0, 79) <= input(13);
output(0, 80) <= input(35);
output(0, 81) <= input(33);
output(0, 82) <= input(16);
output(0, 83) <= input(17);
output(0, 84) <= input(18);
output(0, 85) <= input(19);
output(0, 86) <= input(20);
output(0, 87) <= input(21);
output(0, 88) <= input(22);
output(0, 89) <= input(23);
output(0, 90) <= input(24);
output(0, 91) <= input(25);
output(0, 92) <= input(26);
output(0, 93) <= input(27);
output(0, 94) <= input(28);
output(0, 95) <= input(29);
output(0, 96) <= input(36);
output(0, 97) <= input(34);
output(0, 98) <= input(32);
output(0, 99) <= input(0);
output(0, 100) <= input(1);
output(0, 101) <= input(2);
output(0, 102) <= input(3);
output(0, 103) <= input(4);
output(0, 104) <= input(5);
output(0, 105) <= input(6);
output(0, 106) <= input(7);
output(0, 107) <= input(8);
output(0, 108) <= input(9);
output(0, 109) <= input(10);
output(0, 110) <= input(11);
output(0, 111) <= input(12);
output(0, 112) <= input(37);
output(0, 113) <= input(35);
output(0, 114) <= input(33);
output(0, 115) <= input(16);
output(0, 116) <= input(17);
output(0, 117) <= input(18);
output(0, 118) <= input(19);
output(0, 119) <= input(20);
output(0, 120) <= input(21);
output(0, 121) <= input(22);
output(0, 122) <= input(23);
output(0, 123) <= input(24);
output(0, 124) <= input(25);
output(0, 125) <= input(26);
output(0, 126) <= input(27);
output(0, 127) <= input(28);
output(0, 128) <= input(38);
output(0, 129) <= input(37);
output(0, 130) <= input(35);
output(0, 131) <= input(33);
output(0, 132) <= input(16);
output(0, 133) <= input(17);
output(0, 134) <= input(18);
output(0, 135) <= input(19);
output(0, 136) <= input(20);
output(0, 137) <= input(21);
output(0, 138) <= input(22);
output(0, 139) <= input(23);
output(0, 140) <= input(24);
output(0, 141) <= input(25);
output(0, 142) <= input(26);
output(0, 143) <= input(27);
output(0, 144) <= input(39);
output(0, 145) <= input(40);
output(0, 146) <= input(36);
output(0, 147) <= input(34);
output(0, 148) <= input(32);
output(0, 149) <= input(0);
output(0, 150) <= input(1);
output(0, 151) <= input(2);
output(0, 152) <= input(3);
output(0, 153) <= input(4);
output(0, 154) <= input(5);
output(0, 155) <= input(6);
output(0, 156) <= input(7);
output(0, 157) <= input(8);
output(0, 158) <= input(9);
output(0, 159) <= input(10);
output(0, 160) <= input(41);
output(0, 161) <= input(38);
output(0, 162) <= input(37);
output(0, 163) <= input(35);
output(0, 164) <= input(33);
output(0, 165) <= input(16);
output(0, 166) <= input(17);
output(0, 167) <= input(18);
output(0, 168) <= input(19);
output(0, 169) <= input(20);
output(0, 170) <= input(21);
output(0, 171) <= input(22);
output(0, 172) <= input(23);
output(0, 173) <= input(24);
output(0, 174) <= input(25);
output(0, 175) <= input(26);
output(0, 176) <= input(42);
output(0, 177) <= input(39);
output(0, 178) <= input(40);
output(0, 179) <= input(36);
output(0, 180) <= input(34);
output(0, 181) <= input(32);
output(0, 182) <= input(0);
output(0, 183) <= input(1);
output(0, 184) <= input(2);
output(0, 185) <= input(3);
output(0, 186) <= input(4);
output(0, 187) <= input(5);
output(0, 188) <= input(6);
output(0, 189) <= input(7);
output(0, 190) <= input(8);
output(0, 191) <= input(9);
output(0, 192) <= input(43);
output(0, 193) <= input(41);
output(0, 194) <= input(38);
output(0, 195) <= input(37);
output(0, 196) <= input(35);
output(0, 197) <= input(33);
output(0, 198) <= input(16);
output(0, 199) <= input(17);
output(0, 200) <= input(18);
output(0, 201) <= input(19);
output(0, 202) <= input(20);
output(0, 203) <= input(21);
output(0, 204) <= input(22);
output(0, 205) <= input(23);
output(0, 206) <= input(24);
output(0, 207) <= input(25);
output(0, 208) <= input(44);
output(0, 209) <= input(42);
output(0, 210) <= input(39);
output(0, 211) <= input(40);
output(0, 212) <= input(36);
output(0, 213) <= input(34);
output(0, 214) <= input(32);
output(0, 215) <= input(0);
output(0, 216) <= input(1);
output(0, 217) <= input(2);
output(0, 218) <= input(3);
output(0, 219) <= input(4);
output(0, 220) <= input(5);
output(0, 221) <= input(6);
output(0, 222) <= input(7);
output(0, 223) <= input(8);
output(0, 224) <= input(45);
output(0, 225) <= input(43);
output(0, 226) <= input(41);
output(0, 227) <= input(38);
output(0, 228) <= input(37);
output(0, 229) <= input(35);
output(0, 230) <= input(33);
output(0, 231) <= input(16);
output(0, 232) <= input(17);
output(0, 233) <= input(18);
output(0, 234) <= input(19);
output(0, 235) <= input(20);
output(0, 236) <= input(21);
output(0, 237) <= input(22);
output(0, 238) <= input(23);
output(0, 239) <= input(24);
output(0, 240) <= input(46);
output(0, 241) <= input(44);
output(0, 242) <= input(42);
output(0, 243) <= input(39);
output(0, 244) <= input(40);
output(0, 245) <= input(36);
output(0, 246) <= input(34);
output(0, 247) <= input(32);
output(0, 248) <= input(0);
output(0, 249) <= input(1);
output(0, 250) <= input(2);
output(0, 251) <= input(3);
output(0, 252) <= input(4);
output(0, 253) <= input(5);
output(0, 254) <= input(6);
output(0, 255) <= input(7);
output(1, 0) <= input(18);
output(1, 1) <= input(19);
output(1, 2) <= input(20);
output(1, 3) <= input(21);
output(1, 4) <= input(22);
output(1, 5) <= input(23);
output(1, 6) <= input(24);
output(1, 7) <= input(25);
output(1, 8) <= input(26);
output(1, 9) <= input(27);
output(1, 10) <= input(28);
output(1, 11) <= input(29);
output(1, 12) <= input(30);
output(1, 13) <= input(31);
output(1, 14) <= input(47);
output(1, 15) <= input(48);
output(1, 16) <= input(1);
output(1, 17) <= input(2);
output(1, 18) <= input(3);
output(1, 19) <= input(4);
output(1, 20) <= input(5);
output(1, 21) <= input(6);
output(1, 22) <= input(7);
output(1, 23) <= input(8);
output(1, 24) <= input(9);
output(1, 25) <= input(10);
output(1, 26) <= input(11);
output(1, 27) <= input(12);
output(1, 28) <= input(13);
output(1, 29) <= input(14);
output(1, 30) <= input(15);
output(1, 31) <= input(49);
output(1, 32) <= input(17);
output(1, 33) <= input(18);
output(1, 34) <= input(19);
output(1, 35) <= input(20);
output(1, 36) <= input(21);
output(1, 37) <= input(22);
output(1, 38) <= input(23);
output(1, 39) <= input(24);
output(1, 40) <= input(25);
output(1, 41) <= input(26);
output(1, 42) <= input(27);
output(1, 43) <= input(28);
output(1, 44) <= input(29);
output(1, 45) <= input(30);
output(1, 46) <= input(31);
output(1, 47) <= input(47);
output(1, 48) <= input(0);
output(1, 49) <= input(1);
output(1, 50) <= input(2);
output(1, 51) <= input(3);
output(1, 52) <= input(4);
output(1, 53) <= input(5);
output(1, 54) <= input(6);
output(1, 55) <= input(7);
output(1, 56) <= input(8);
output(1, 57) <= input(9);
output(1, 58) <= input(10);
output(1, 59) <= input(11);
output(1, 60) <= input(12);
output(1, 61) <= input(13);
output(1, 62) <= input(14);
output(1, 63) <= input(15);
output(1, 64) <= input(16);
output(1, 65) <= input(17);
output(1, 66) <= input(18);
output(1, 67) <= input(19);
output(1, 68) <= input(20);
output(1, 69) <= input(21);
output(1, 70) <= input(22);
output(1, 71) <= input(23);
output(1, 72) <= input(24);
output(1, 73) <= input(25);
output(1, 74) <= input(26);
output(1, 75) <= input(27);
output(1, 76) <= input(28);
output(1, 77) <= input(29);
output(1, 78) <= input(30);
output(1, 79) <= input(31);
output(1, 80) <= input(32);
output(1, 81) <= input(0);
output(1, 82) <= input(1);
output(1, 83) <= input(2);
output(1, 84) <= input(3);
output(1, 85) <= input(4);
output(1, 86) <= input(5);
output(1, 87) <= input(6);
output(1, 88) <= input(7);
output(1, 89) <= input(8);
output(1, 90) <= input(9);
output(1, 91) <= input(10);
output(1, 92) <= input(11);
output(1, 93) <= input(12);
output(1, 94) <= input(13);
output(1, 95) <= input(14);
output(1, 96) <= input(33);
output(1, 97) <= input(16);
output(1, 98) <= input(17);
output(1, 99) <= input(18);
output(1, 100) <= input(19);
output(1, 101) <= input(20);
output(1, 102) <= input(21);
output(1, 103) <= input(22);
output(1, 104) <= input(23);
output(1, 105) <= input(24);
output(1, 106) <= input(25);
output(1, 107) <= input(26);
output(1, 108) <= input(27);
output(1, 109) <= input(28);
output(1, 110) <= input(29);
output(1, 111) <= input(30);
output(1, 112) <= input(34);
output(1, 113) <= input(32);
output(1, 114) <= input(0);
output(1, 115) <= input(1);
output(1, 116) <= input(2);
output(1, 117) <= input(3);
output(1, 118) <= input(4);
output(1, 119) <= input(5);
output(1, 120) <= input(6);
output(1, 121) <= input(7);
output(1, 122) <= input(8);
output(1, 123) <= input(9);
output(1, 124) <= input(10);
output(1, 125) <= input(11);
output(1, 126) <= input(12);
output(1, 127) <= input(13);
output(1, 128) <= input(35);
output(1, 129) <= input(33);
output(1, 130) <= input(16);
output(1, 131) <= input(17);
output(1, 132) <= input(18);
output(1, 133) <= input(19);
output(1, 134) <= input(20);
output(1, 135) <= input(21);
output(1, 136) <= input(22);
output(1, 137) <= input(23);
output(1, 138) <= input(24);
output(1, 139) <= input(25);
output(1, 140) <= input(26);
output(1, 141) <= input(27);
output(1, 142) <= input(28);
output(1, 143) <= input(29);
output(1, 144) <= input(36);
output(1, 145) <= input(34);
output(1, 146) <= input(32);
output(1, 147) <= input(0);
output(1, 148) <= input(1);
output(1, 149) <= input(2);
output(1, 150) <= input(3);
output(1, 151) <= input(4);
output(1, 152) <= input(5);
output(1, 153) <= input(6);
output(1, 154) <= input(7);
output(1, 155) <= input(8);
output(1, 156) <= input(9);
output(1, 157) <= input(10);
output(1, 158) <= input(11);
output(1, 159) <= input(12);
output(1, 160) <= input(37);
output(1, 161) <= input(35);
output(1, 162) <= input(33);
output(1, 163) <= input(16);
output(1, 164) <= input(17);
output(1, 165) <= input(18);
output(1, 166) <= input(19);
output(1, 167) <= input(20);
output(1, 168) <= input(21);
output(1, 169) <= input(22);
output(1, 170) <= input(23);
output(1, 171) <= input(24);
output(1, 172) <= input(25);
output(1, 173) <= input(26);
output(1, 174) <= input(27);
output(1, 175) <= input(28);
output(1, 176) <= input(40);
output(1, 177) <= input(36);
output(1, 178) <= input(34);
output(1, 179) <= input(32);
output(1, 180) <= input(0);
output(1, 181) <= input(1);
output(1, 182) <= input(2);
output(1, 183) <= input(3);
output(1, 184) <= input(4);
output(1, 185) <= input(5);
output(1, 186) <= input(6);
output(1, 187) <= input(7);
output(1, 188) <= input(8);
output(1, 189) <= input(9);
output(1, 190) <= input(10);
output(1, 191) <= input(11);
output(1, 192) <= input(38);
output(1, 193) <= input(37);
output(1, 194) <= input(35);
output(1, 195) <= input(33);
output(1, 196) <= input(16);
output(1, 197) <= input(17);
output(1, 198) <= input(18);
output(1, 199) <= input(19);
output(1, 200) <= input(20);
output(1, 201) <= input(21);
output(1, 202) <= input(22);
output(1, 203) <= input(23);
output(1, 204) <= input(24);
output(1, 205) <= input(25);
output(1, 206) <= input(26);
output(1, 207) <= input(27);
output(1, 208) <= input(39);
output(1, 209) <= input(40);
output(1, 210) <= input(36);
output(1, 211) <= input(34);
output(1, 212) <= input(32);
output(1, 213) <= input(0);
output(1, 214) <= input(1);
output(1, 215) <= input(2);
output(1, 216) <= input(3);
output(1, 217) <= input(4);
output(1, 218) <= input(5);
output(1, 219) <= input(6);
output(1, 220) <= input(7);
output(1, 221) <= input(8);
output(1, 222) <= input(9);
output(1, 223) <= input(10);
output(1, 224) <= input(41);
output(1, 225) <= input(38);
output(1, 226) <= input(37);
output(1, 227) <= input(35);
output(1, 228) <= input(33);
output(1, 229) <= input(16);
output(1, 230) <= input(17);
output(1, 231) <= input(18);
output(1, 232) <= input(19);
output(1, 233) <= input(20);
output(1, 234) <= input(21);
output(1, 235) <= input(22);
output(1, 236) <= input(23);
output(1, 237) <= input(24);
output(1, 238) <= input(25);
output(1, 239) <= input(26);
output(1, 240) <= input(42);
output(1, 241) <= input(39);
output(1, 242) <= input(40);
output(1, 243) <= input(36);
output(1, 244) <= input(34);
output(1, 245) <= input(32);
output(1, 246) <= input(0);
output(1, 247) <= input(1);
output(1, 248) <= input(2);
output(1, 249) <= input(3);
output(1, 250) <= input(4);
output(1, 251) <= input(5);
output(1, 252) <= input(6);
output(1, 253) <= input(7);
output(1, 254) <= input(8);
output(1, 255) <= input(9);
when "1011" =>
output(0, 0) <= input(0);
output(0, 1) <= input(1);
output(0, 2) <= input(2);
output(0, 3) <= input(3);
output(0, 4) <= input(4);
output(0, 5) <= input(5);
output(0, 6) <= input(6);
output(0, 7) <= input(7);
output(0, 8) <= input(8);
output(0, 9) <= input(9);
output(0, 10) <= input(10);
output(0, 11) <= input(11);
output(0, 12) <= input(12);
output(0, 13) <= input(13);
output(0, 14) <= input(14);
output(0, 15) <= input(15);
output(0, 16) <= input(16);
output(0, 17) <= input(17);
output(0, 18) <= input(18);
output(0, 19) <= input(19);
output(0, 20) <= input(20);
output(0, 21) <= input(21);
output(0, 22) <= input(22);
output(0, 23) <= input(23);
output(0, 24) <= input(24);
output(0, 25) <= input(25);
output(0, 26) <= input(26);
output(0, 27) <= input(27);
output(0, 28) <= input(28);
output(0, 29) <= input(29);
output(0, 30) <= input(30);
output(0, 31) <= input(31);
output(0, 32) <= input(32);
output(0, 33) <= input(0);
output(0, 34) <= input(1);
output(0, 35) <= input(2);
output(0, 36) <= input(3);
output(0, 37) <= input(4);
output(0, 38) <= input(5);
output(0, 39) <= input(6);
output(0, 40) <= input(7);
output(0, 41) <= input(8);
output(0, 42) <= input(9);
output(0, 43) <= input(10);
output(0, 44) <= input(11);
output(0, 45) <= input(12);
output(0, 46) <= input(13);
output(0, 47) <= input(14);
output(0, 48) <= input(33);
output(0, 49) <= input(16);
output(0, 50) <= input(17);
output(0, 51) <= input(18);
output(0, 52) <= input(19);
output(0, 53) <= input(20);
output(0, 54) <= input(21);
output(0, 55) <= input(22);
output(0, 56) <= input(23);
output(0, 57) <= input(24);
output(0, 58) <= input(25);
output(0, 59) <= input(26);
output(0, 60) <= input(27);
output(0, 61) <= input(28);
output(0, 62) <= input(29);
output(0, 63) <= input(30);
output(0, 64) <= input(34);
output(0, 65) <= input(32);
output(0, 66) <= input(0);
output(0, 67) <= input(1);
output(0, 68) <= input(2);
output(0, 69) <= input(3);
output(0, 70) <= input(4);
output(0, 71) <= input(5);
output(0, 72) <= input(6);
output(0, 73) <= input(7);
output(0, 74) <= input(8);
output(0, 75) <= input(9);
output(0, 76) <= input(10);
output(0, 77) <= input(11);
output(0, 78) <= input(12);
output(0, 79) <= input(13);
output(0, 80) <= input(35);
output(0, 81) <= input(33);
output(0, 82) <= input(16);
output(0, 83) <= input(17);
output(0, 84) <= input(18);
output(0, 85) <= input(19);
output(0, 86) <= input(20);
output(0, 87) <= input(21);
output(0, 88) <= input(22);
output(0, 89) <= input(23);
output(0, 90) <= input(24);
output(0, 91) <= input(25);
output(0, 92) <= input(26);
output(0, 93) <= input(27);
output(0, 94) <= input(28);
output(0, 95) <= input(29);
output(0, 96) <= input(36);
output(0, 97) <= input(34);
output(0, 98) <= input(32);
output(0, 99) <= input(0);
output(0, 100) <= input(1);
output(0, 101) <= input(2);
output(0, 102) <= input(3);
output(0, 103) <= input(4);
output(0, 104) <= input(5);
output(0, 105) <= input(6);
output(0, 106) <= input(7);
output(0, 107) <= input(8);
output(0, 108) <= input(9);
output(0, 109) <= input(10);
output(0, 110) <= input(11);
output(0, 111) <= input(12);
output(0, 112) <= input(36);
output(0, 113) <= input(34);
output(0, 114) <= input(32);
output(0, 115) <= input(0);
output(0, 116) <= input(1);
output(0, 117) <= input(2);
output(0, 118) <= input(3);
output(0, 119) <= input(4);
output(0, 120) <= input(5);
output(0, 121) <= input(6);
output(0, 122) <= input(7);
output(0, 123) <= input(8);
output(0, 124) <= input(9);
output(0, 125) <= input(10);
output(0, 126) <= input(11);
output(0, 127) <= input(12);
output(0, 128) <= input(37);
output(0, 129) <= input(35);
output(0, 130) <= input(33);
output(0, 131) <= input(16);
output(0, 132) <= input(17);
output(0, 133) <= input(18);
output(0, 134) <= input(19);
output(0, 135) <= input(20);
output(0, 136) <= input(21);
output(0, 137) <= input(22);
output(0, 138) <= input(23);
output(0, 139) <= input(24);
output(0, 140) <= input(25);
output(0, 141) <= input(26);
output(0, 142) <= input(27);
output(0, 143) <= input(28);
output(0, 144) <= input(38);
output(0, 145) <= input(36);
output(0, 146) <= input(34);
output(0, 147) <= input(32);
output(0, 148) <= input(0);
output(0, 149) <= input(1);
output(0, 150) <= input(2);
output(0, 151) <= input(3);
output(0, 152) <= input(4);
output(0, 153) <= input(5);
output(0, 154) <= input(6);
output(0, 155) <= input(7);
output(0, 156) <= input(8);
output(0, 157) <= input(9);
output(0, 158) <= input(10);
output(0, 159) <= input(11);
output(0, 160) <= input(39);
output(0, 161) <= input(37);
output(0, 162) <= input(35);
output(0, 163) <= input(33);
output(0, 164) <= input(16);
output(0, 165) <= input(17);
output(0, 166) <= input(18);
output(0, 167) <= input(19);
output(0, 168) <= input(20);
output(0, 169) <= input(21);
output(0, 170) <= input(22);
output(0, 171) <= input(23);
output(0, 172) <= input(24);
output(0, 173) <= input(25);
output(0, 174) <= input(26);
output(0, 175) <= input(27);
output(0, 176) <= input(40);
output(0, 177) <= input(38);
output(0, 178) <= input(36);
output(0, 179) <= input(34);
output(0, 180) <= input(32);
output(0, 181) <= input(0);
output(0, 182) <= input(1);
output(0, 183) <= input(2);
output(0, 184) <= input(3);
output(0, 185) <= input(4);
output(0, 186) <= input(5);
output(0, 187) <= input(6);
output(0, 188) <= input(7);
output(0, 189) <= input(8);
output(0, 190) <= input(9);
output(0, 191) <= input(10);
output(0, 192) <= input(41);
output(0, 193) <= input(39);
output(0, 194) <= input(37);
output(0, 195) <= input(35);
output(0, 196) <= input(33);
output(0, 197) <= input(16);
output(0, 198) <= input(17);
output(0, 199) <= input(18);
output(0, 200) <= input(19);
output(0, 201) <= input(20);
output(0, 202) <= input(21);
output(0, 203) <= input(22);
output(0, 204) <= input(23);
output(0, 205) <= input(24);
output(0, 206) <= input(25);
output(0, 207) <= input(26);
output(0, 208) <= input(42);
output(0, 209) <= input(40);
output(0, 210) <= input(38);
output(0, 211) <= input(36);
output(0, 212) <= input(34);
output(0, 213) <= input(32);
output(0, 214) <= input(0);
output(0, 215) <= input(1);
output(0, 216) <= input(2);
output(0, 217) <= input(3);
output(0, 218) <= input(4);
output(0, 219) <= input(5);
output(0, 220) <= input(6);
output(0, 221) <= input(7);
output(0, 222) <= input(8);
output(0, 223) <= input(9);
output(0, 224) <= input(43);
output(0, 225) <= input(41);
output(0, 226) <= input(39);
output(0, 227) <= input(37);
output(0, 228) <= input(35);
output(0, 229) <= input(33);
output(0, 230) <= input(16);
output(0, 231) <= input(17);
output(0, 232) <= input(18);
output(0, 233) <= input(19);
output(0, 234) <= input(20);
output(0, 235) <= input(21);
output(0, 236) <= input(22);
output(0, 237) <= input(23);
output(0, 238) <= input(24);
output(0, 239) <= input(25);
output(0, 240) <= input(43);
output(0, 241) <= input(41);
output(0, 242) <= input(39);
output(0, 243) <= input(37);
output(0, 244) <= input(35);
output(0, 245) <= input(33);
output(0, 246) <= input(16);
output(0, 247) <= input(17);
output(0, 248) <= input(18);
output(0, 249) <= input(19);
output(0, 250) <= input(20);
output(0, 251) <= input(21);
output(0, 252) <= input(22);
output(0, 253) <= input(23);
output(0, 254) <= input(24);
output(0, 255) <= input(25);
output(1, 0) <= input(1);
output(1, 1) <= input(2);
output(1, 2) <= input(3);
output(1, 3) <= input(4);
output(1, 4) <= input(5);
output(1, 5) <= input(6);
output(1, 6) <= input(7);
output(1, 7) <= input(8);
output(1, 8) <= input(9);
output(1, 9) <= input(10);
output(1, 10) <= input(11);
output(1, 11) <= input(12);
output(1, 12) <= input(13);
output(1, 13) <= input(14);
output(1, 14) <= input(15);
output(1, 15) <= input(44);
output(1, 16) <= input(17);
output(1, 17) <= input(18);
output(1, 18) <= input(19);
output(1, 19) <= input(20);
output(1, 20) <= input(21);
output(1, 21) <= input(22);
output(1, 22) <= input(23);
output(1, 23) <= input(24);
output(1, 24) <= input(25);
output(1, 25) <= input(26);
output(1, 26) <= input(27);
output(1, 27) <= input(28);
output(1, 28) <= input(29);
output(1, 29) <= input(30);
output(1, 30) <= input(31);
output(1, 31) <= input(45);
output(1, 32) <= input(0);
output(1, 33) <= input(1);
output(1, 34) <= input(2);
output(1, 35) <= input(3);
output(1, 36) <= input(4);
output(1, 37) <= input(5);
output(1, 38) <= input(6);
output(1, 39) <= input(7);
output(1, 40) <= input(8);
output(1, 41) <= input(9);
output(1, 42) <= input(10);
output(1, 43) <= input(11);
output(1, 44) <= input(12);
output(1, 45) <= input(13);
output(1, 46) <= input(14);
output(1, 47) <= input(15);
output(1, 48) <= input(0);
output(1, 49) <= input(1);
output(1, 50) <= input(2);
output(1, 51) <= input(3);
output(1, 52) <= input(4);
output(1, 53) <= input(5);
output(1, 54) <= input(6);
output(1, 55) <= input(7);
output(1, 56) <= input(8);
output(1, 57) <= input(9);
output(1, 58) <= input(10);
output(1, 59) <= input(11);
output(1, 60) <= input(12);
output(1, 61) <= input(13);
output(1, 62) <= input(14);
output(1, 63) <= input(15);
output(1, 64) <= input(16);
output(1, 65) <= input(17);
output(1, 66) <= input(18);
output(1, 67) <= input(19);
output(1, 68) <= input(20);
output(1, 69) <= input(21);
output(1, 70) <= input(22);
output(1, 71) <= input(23);
output(1, 72) <= input(24);
output(1, 73) <= input(25);
output(1, 74) <= input(26);
output(1, 75) <= input(27);
output(1, 76) <= input(28);
output(1, 77) <= input(29);
output(1, 78) <= input(30);
output(1, 79) <= input(31);
output(1, 80) <= input(32);
output(1, 81) <= input(0);
output(1, 82) <= input(1);
output(1, 83) <= input(2);
output(1, 84) <= input(3);
output(1, 85) <= input(4);
output(1, 86) <= input(5);
output(1, 87) <= input(6);
output(1, 88) <= input(7);
output(1, 89) <= input(8);
output(1, 90) <= input(9);
output(1, 91) <= input(10);
output(1, 92) <= input(11);
output(1, 93) <= input(12);
output(1, 94) <= input(13);
output(1, 95) <= input(14);
output(1, 96) <= input(33);
output(1, 97) <= input(16);
output(1, 98) <= input(17);
output(1, 99) <= input(18);
output(1, 100) <= input(19);
output(1, 101) <= input(20);
output(1, 102) <= input(21);
output(1, 103) <= input(22);
output(1, 104) <= input(23);
output(1, 105) <= input(24);
output(1, 106) <= input(25);
output(1, 107) <= input(26);
output(1, 108) <= input(27);
output(1, 109) <= input(28);
output(1, 110) <= input(29);
output(1, 111) <= input(30);
output(1, 112) <= input(33);
output(1, 113) <= input(16);
output(1, 114) <= input(17);
output(1, 115) <= input(18);
output(1, 116) <= input(19);
output(1, 117) <= input(20);
output(1, 118) <= input(21);
output(1, 119) <= input(22);
output(1, 120) <= input(23);
output(1, 121) <= input(24);
output(1, 122) <= input(25);
output(1, 123) <= input(26);
output(1, 124) <= input(27);
output(1, 125) <= input(28);
output(1, 126) <= input(29);
output(1, 127) <= input(30);
output(1, 128) <= input(34);
output(1, 129) <= input(32);
output(1, 130) <= input(0);
output(1, 131) <= input(1);
output(1, 132) <= input(2);
output(1, 133) <= input(3);
output(1, 134) <= input(4);
output(1, 135) <= input(5);
output(1, 136) <= input(6);
output(1, 137) <= input(7);
output(1, 138) <= input(8);
output(1, 139) <= input(9);
output(1, 140) <= input(10);
output(1, 141) <= input(11);
output(1, 142) <= input(12);
output(1, 143) <= input(13);
output(1, 144) <= input(35);
output(1, 145) <= input(33);
output(1, 146) <= input(16);
output(1, 147) <= input(17);
output(1, 148) <= input(18);
output(1, 149) <= input(19);
output(1, 150) <= input(20);
output(1, 151) <= input(21);
output(1, 152) <= input(22);
output(1, 153) <= input(23);
output(1, 154) <= input(24);
output(1, 155) <= input(25);
output(1, 156) <= input(26);
output(1, 157) <= input(27);
output(1, 158) <= input(28);
output(1, 159) <= input(29);
output(1, 160) <= input(36);
output(1, 161) <= input(34);
output(1, 162) <= input(32);
output(1, 163) <= input(0);
output(1, 164) <= input(1);
output(1, 165) <= input(2);
output(1, 166) <= input(3);
output(1, 167) <= input(4);
output(1, 168) <= input(5);
output(1, 169) <= input(6);
output(1, 170) <= input(7);
output(1, 171) <= input(8);
output(1, 172) <= input(9);
output(1, 173) <= input(10);
output(1, 174) <= input(11);
output(1, 175) <= input(12);
output(1, 176) <= input(36);
output(1, 177) <= input(34);
output(1, 178) <= input(32);
output(1, 179) <= input(0);
output(1, 180) <= input(1);
output(1, 181) <= input(2);
output(1, 182) <= input(3);
output(1, 183) <= input(4);
output(1, 184) <= input(5);
output(1, 185) <= input(6);
output(1, 186) <= input(7);
output(1, 187) <= input(8);
output(1, 188) <= input(9);
output(1, 189) <= input(10);
output(1, 190) <= input(11);
output(1, 191) <= input(12);
output(1, 192) <= input(37);
output(1, 193) <= input(35);
output(1, 194) <= input(33);
output(1, 195) <= input(16);
output(1, 196) <= input(17);
output(1, 197) <= input(18);
output(1, 198) <= input(19);
output(1, 199) <= input(20);
output(1, 200) <= input(21);
output(1, 201) <= input(22);
output(1, 202) <= input(23);
output(1, 203) <= input(24);
output(1, 204) <= input(25);
output(1, 205) <= input(26);
output(1, 206) <= input(27);
output(1, 207) <= input(28);
output(1, 208) <= input(38);
output(1, 209) <= input(36);
output(1, 210) <= input(34);
output(1, 211) <= input(32);
output(1, 212) <= input(0);
output(1, 213) <= input(1);
output(1, 214) <= input(2);
output(1, 215) <= input(3);
output(1, 216) <= input(4);
output(1, 217) <= input(5);
output(1, 218) <= input(6);
output(1, 219) <= input(7);
output(1, 220) <= input(8);
output(1, 221) <= input(9);
output(1, 222) <= input(10);
output(1, 223) <= input(11);
output(1, 224) <= input(39);
output(1, 225) <= input(37);
output(1, 226) <= input(35);
output(1, 227) <= input(33);
output(1, 228) <= input(16);
output(1, 229) <= input(17);
output(1, 230) <= input(18);
output(1, 231) <= input(19);
output(1, 232) <= input(20);
output(1, 233) <= input(21);
output(1, 234) <= input(22);
output(1, 235) <= input(23);
output(1, 236) <= input(24);
output(1, 237) <= input(25);
output(1, 238) <= input(26);
output(1, 239) <= input(27);
output(1, 240) <= input(39);
output(1, 241) <= input(37);
output(1, 242) <= input(35);
output(1, 243) <= input(33);
output(1, 244) <= input(16);
output(1, 245) <= input(17);
output(1, 246) <= input(18);
output(1, 247) <= input(19);
output(1, 248) <= input(20);
output(1, 249) <= input(21);
output(1, 250) <= input(22);
output(1, 251) <= input(23);
output(1, 252) <= input(24);
output(1, 253) <= input(25);
output(1, 254) <= input(26);
output(1, 255) <= input(27);
output(2, 0) <= input(2);
output(2, 1) <= input(3);
output(2, 2) <= input(4);
output(2, 3) <= input(5);
output(2, 4) <= input(6);
output(2, 5) <= input(7);
output(2, 6) <= input(8);
output(2, 7) <= input(9);
output(2, 8) <= input(10);
output(2, 9) <= input(11);
output(2, 10) <= input(12);
output(2, 11) <= input(13);
output(2, 12) <= input(14);
output(2, 13) <= input(15);
output(2, 14) <= input(44);
output(2, 15) <= input(46);
output(2, 16) <= input(18);
output(2, 17) <= input(19);
output(2, 18) <= input(20);
output(2, 19) <= input(21);
output(2, 20) <= input(22);
output(2, 21) <= input(23);
output(2, 22) <= input(24);
output(2, 23) <= input(25);
output(2, 24) <= input(26);
output(2, 25) <= input(27);
output(2, 26) <= input(28);
output(2, 27) <= input(29);
output(2, 28) <= input(30);
output(2, 29) <= input(31);
output(2, 30) <= input(45);
output(2, 31) <= input(47);
output(2, 32) <= input(18);
output(2, 33) <= input(19);
output(2, 34) <= input(20);
output(2, 35) <= input(21);
output(2, 36) <= input(22);
output(2, 37) <= input(23);
output(2, 38) <= input(24);
output(2, 39) <= input(25);
output(2, 40) <= input(26);
output(2, 41) <= input(27);
output(2, 42) <= input(28);
output(2, 43) <= input(29);
output(2, 44) <= input(30);
output(2, 45) <= input(31);
output(2, 46) <= input(45);
output(2, 47) <= input(47);
output(2, 48) <= input(1);
output(2, 49) <= input(2);
output(2, 50) <= input(3);
output(2, 51) <= input(4);
output(2, 52) <= input(5);
output(2, 53) <= input(6);
output(2, 54) <= input(7);
output(2, 55) <= input(8);
output(2, 56) <= input(9);
output(2, 57) <= input(10);
output(2, 58) <= input(11);
output(2, 59) <= input(12);
output(2, 60) <= input(13);
output(2, 61) <= input(14);
output(2, 62) <= input(15);
output(2, 63) <= input(44);
output(2, 64) <= input(17);
output(2, 65) <= input(18);
output(2, 66) <= input(19);
output(2, 67) <= input(20);
output(2, 68) <= input(21);
output(2, 69) <= input(22);
output(2, 70) <= input(23);
output(2, 71) <= input(24);
output(2, 72) <= input(25);
output(2, 73) <= input(26);
output(2, 74) <= input(27);
output(2, 75) <= input(28);
output(2, 76) <= input(29);
output(2, 77) <= input(30);
output(2, 78) <= input(31);
output(2, 79) <= input(45);
output(2, 80) <= input(17);
output(2, 81) <= input(18);
output(2, 82) <= input(19);
output(2, 83) <= input(20);
output(2, 84) <= input(21);
output(2, 85) <= input(22);
output(2, 86) <= input(23);
output(2, 87) <= input(24);
output(2, 88) <= input(25);
output(2, 89) <= input(26);
output(2, 90) <= input(27);
output(2, 91) <= input(28);
output(2, 92) <= input(29);
output(2, 93) <= input(30);
output(2, 94) <= input(31);
output(2, 95) <= input(45);
output(2, 96) <= input(0);
output(2, 97) <= input(1);
output(2, 98) <= input(2);
output(2, 99) <= input(3);
output(2, 100) <= input(4);
output(2, 101) <= input(5);
output(2, 102) <= input(6);
output(2, 103) <= input(7);
output(2, 104) <= input(8);
output(2, 105) <= input(9);
output(2, 106) <= input(10);
output(2, 107) <= input(11);
output(2, 108) <= input(12);
output(2, 109) <= input(13);
output(2, 110) <= input(14);
output(2, 111) <= input(15);
output(2, 112) <= input(0);
output(2, 113) <= input(1);
output(2, 114) <= input(2);
output(2, 115) <= input(3);
output(2, 116) <= input(4);
output(2, 117) <= input(5);
output(2, 118) <= input(6);
output(2, 119) <= input(7);
output(2, 120) <= input(8);
output(2, 121) <= input(9);
output(2, 122) <= input(10);
output(2, 123) <= input(11);
output(2, 124) <= input(12);
output(2, 125) <= input(13);
output(2, 126) <= input(14);
output(2, 127) <= input(15);
output(2, 128) <= input(16);
output(2, 129) <= input(17);
output(2, 130) <= input(18);
output(2, 131) <= input(19);
output(2, 132) <= input(20);
output(2, 133) <= input(21);
output(2, 134) <= input(22);
output(2, 135) <= input(23);
output(2, 136) <= input(24);
output(2, 137) <= input(25);
output(2, 138) <= input(26);
output(2, 139) <= input(27);
output(2, 140) <= input(28);
output(2, 141) <= input(29);
output(2, 142) <= input(30);
output(2, 143) <= input(31);
output(2, 144) <= input(32);
output(2, 145) <= input(0);
output(2, 146) <= input(1);
output(2, 147) <= input(2);
output(2, 148) <= input(3);
output(2, 149) <= input(4);
output(2, 150) <= input(5);
output(2, 151) <= input(6);
output(2, 152) <= input(7);
output(2, 153) <= input(8);
output(2, 154) <= input(9);
output(2, 155) <= input(10);
output(2, 156) <= input(11);
output(2, 157) <= input(12);
output(2, 158) <= input(13);
output(2, 159) <= input(14);
output(2, 160) <= input(32);
output(2, 161) <= input(0);
output(2, 162) <= input(1);
output(2, 163) <= input(2);
output(2, 164) <= input(3);
output(2, 165) <= input(4);
output(2, 166) <= input(5);
output(2, 167) <= input(6);
output(2, 168) <= input(7);
output(2, 169) <= input(8);
output(2, 170) <= input(9);
output(2, 171) <= input(10);
output(2, 172) <= input(11);
output(2, 173) <= input(12);
output(2, 174) <= input(13);
output(2, 175) <= input(14);
output(2, 176) <= input(33);
output(2, 177) <= input(16);
output(2, 178) <= input(17);
output(2, 179) <= input(18);
output(2, 180) <= input(19);
output(2, 181) <= input(20);
output(2, 182) <= input(21);
output(2, 183) <= input(22);
output(2, 184) <= input(23);
output(2, 185) <= input(24);
output(2, 186) <= input(25);
output(2, 187) <= input(26);
output(2, 188) <= input(27);
output(2, 189) <= input(28);
output(2, 190) <= input(29);
output(2, 191) <= input(30);
output(2, 192) <= input(34);
output(2, 193) <= input(32);
output(2, 194) <= input(0);
output(2, 195) <= input(1);
output(2, 196) <= input(2);
output(2, 197) <= input(3);
output(2, 198) <= input(4);
output(2, 199) <= input(5);
output(2, 200) <= input(6);
output(2, 201) <= input(7);
output(2, 202) <= input(8);
output(2, 203) <= input(9);
output(2, 204) <= input(10);
output(2, 205) <= input(11);
output(2, 206) <= input(12);
output(2, 207) <= input(13);
output(2, 208) <= input(34);
output(2, 209) <= input(32);
output(2, 210) <= input(0);
output(2, 211) <= input(1);
output(2, 212) <= input(2);
output(2, 213) <= input(3);
output(2, 214) <= input(4);
output(2, 215) <= input(5);
output(2, 216) <= input(6);
output(2, 217) <= input(7);
output(2, 218) <= input(8);
output(2, 219) <= input(9);
output(2, 220) <= input(10);
output(2, 221) <= input(11);
output(2, 222) <= input(12);
output(2, 223) <= input(13);
output(2, 224) <= input(35);
output(2, 225) <= input(33);
output(2, 226) <= input(16);
output(2, 227) <= input(17);
output(2, 228) <= input(18);
output(2, 229) <= input(19);
output(2, 230) <= input(20);
output(2, 231) <= input(21);
output(2, 232) <= input(22);
output(2, 233) <= input(23);
output(2, 234) <= input(24);
output(2, 235) <= input(25);
output(2, 236) <= input(26);
output(2, 237) <= input(27);
output(2, 238) <= input(28);
output(2, 239) <= input(29);
output(2, 240) <= input(35);
output(2, 241) <= input(33);
output(2, 242) <= input(16);
output(2, 243) <= input(17);
output(2, 244) <= input(18);
output(2, 245) <= input(19);
output(2, 246) <= input(20);
output(2, 247) <= input(21);
output(2, 248) <= input(22);
output(2, 249) <= input(23);
output(2, 250) <= input(24);
output(2, 251) <= input(25);
output(2, 252) <= input(26);
output(2, 253) <= input(27);
output(2, 254) <= input(28);
output(2, 255) <= input(29);
when "1100" =>
output(0, 0) <= input(0);
output(0, 1) <= input(1);
output(0, 2) <= input(2);
output(0, 3) <= input(3);
output(0, 4) <= input(4);
output(0, 5) <= input(5);
output(0, 6) <= input(6);
output(0, 7) <= input(7);
output(0, 8) <= input(8);
output(0, 9) <= input(9);
output(0, 10) <= input(10);
output(0, 11) <= input(11);
output(0, 12) <= input(12);
output(0, 13) <= input(13);
output(0, 14) <= input(14);
output(0, 15) <= input(15);
output(0, 16) <= input(0);
output(0, 17) <= input(1);
output(0, 18) <= input(2);
output(0, 19) <= input(3);
output(0, 20) <= input(4);
output(0, 21) <= input(5);
output(0, 22) <= input(6);
output(0, 23) <= input(7);
output(0, 24) <= input(8);
output(0, 25) <= input(9);
output(0, 26) <= input(10);
output(0, 27) <= input(11);
output(0, 28) <= input(12);
output(0, 29) <= input(13);
output(0, 30) <= input(14);
output(0, 31) <= input(15);
output(0, 32) <= input(16);
output(0, 33) <= input(17);
output(0, 34) <= input(18);
output(0, 35) <= input(19);
output(0, 36) <= input(20);
output(0, 37) <= input(21);
output(0, 38) <= input(22);
output(0, 39) <= input(23);
output(0, 40) <= input(24);
output(0, 41) <= input(25);
output(0, 42) <= input(26);
output(0, 43) <= input(27);
output(0, 44) <= input(28);
output(0, 45) <= input(29);
output(0, 46) <= input(30);
output(0, 47) <= input(31);
output(0, 48) <= input(16);
output(0, 49) <= input(17);
output(0, 50) <= input(18);
output(0, 51) <= input(19);
output(0, 52) <= input(20);
output(0, 53) <= input(21);
output(0, 54) <= input(22);
output(0, 55) <= input(23);
output(0, 56) <= input(24);
output(0, 57) <= input(25);
output(0, 58) <= input(26);
output(0, 59) <= input(27);
output(0, 60) <= input(28);
output(0, 61) <= input(29);
output(0, 62) <= input(30);
output(0, 63) <= input(31);
output(0, 64) <= input(32);
output(0, 65) <= input(0);
output(0, 66) <= input(1);
output(0, 67) <= input(2);
output(0, 68) <= input(3);
output(0, 69) <= input(4);
output(0, 70) <= input(5);
output(0, 71) <= input(6);
output(0, 72) <= input(7);
output(0, 73) <= input(8);
output(0, 74) <= input(9);
output(0, 75) <= input(10);
output(0, 76) <= input(11);
output(0, 77) <= input(12);
output(0, 78) <= input(13);
output(0, 79) <= input(14);
output(0, 80) <= input(32);
output(0, 81) <= input(0);
output(0, 82) <= input(1);
output(0, 83) <= input(2);
output(0, 84) <= input(3);
output(0, 85) <= input(4);
output(0, 86) <= input(5);
output(0, 87) <= input(6);
output(0, 88) <= input(7);
output(0, 89) <= input(8);
output(0, 90) <= input(9);
output(0, 91) <= input(10);
output(0, 92) <= input(11);
output(0, 93) <= input(12);
output(0, 94) <= input(13);
output(0, 95) <= input(14);
output(0, 96) <= input(33);
output(0, 97) <= input(16);
output(0, 98) <= input(17);
output(0, 99) <= input(18);
output(0, 100) <= input(19);
output(0, 101) <= input(20);
output(0, 102) <= input(21);
output(0, 103) <= input(22);
output(0, 104) <= input(23);
output(0, 105) <= input(24);
output(0, 106) <= input(25);
output(0, 107) <= input(26);
output(0, 108) <= input(27);
output(0, 109) <= input(28);
output(0, 110) <= input(29);
output(0, 111) <= input(30);
output(0, 112) <= input(33);
output(0, 113) <= input(16);
output(0, 114) <= input(17);
output(0, 115) <= input(18);
output(0, 116) <= input(19);
output(0, 117) <= input(20);
output(0, 118) <= input(21);
output(0, 119) <= input(22);
output(0, 120) <= input(23);
output(0, 121) <= input(24);
output(0, 122) <= input(25);
output(0, 123) <= input(26);
output(0, 124) <= input(27);
output(0, 125) <= input(28);
output(0, 126) <= input(29);
output(0, 127) <= input(30);
output(0, 128) <= input(34);
output(0, 129) <= input(32);
output(0, 130) <= input(0);
output(0, 131) <= input(1);
output(0, 132) <= input(2);
output(0, 133) <= input(3);
output(0, 134) <= input(4);
output(0, 135) <= input(5);
output(0, 136) <= input(6);
output(0, 137) <= input(7);
output(0, 138) <= input(8);
output(0, 139) <= input(9);
output(0, 140) <= input(10);
output(0, 141) <= input(11);
output(0, 142) <= input(12);
output(0, 143) <= input(13);
output(0, 144) <= input(34);
output(0, 145) <= input(32);
output(0, 146) <= input(0);
output(0, 147) <= input(1);
output(0, 148) <= input(2);
output(0, 149) <= input(3);
output(0, 150) <= input(4);
output(0, 151) <= input(5);
output(0, 152) <= input(6);
output(0, 153) <= input(7);
output(0, 154) <= input(8);
output(0, 155) <= input(9);
output(0, 156) <= input(10);
output(0, 157) <= input(11);
output(0, 158) <= input(12);
output(0, 159) <= input(13);
output(0, 160) <= input(35);
output(0, 161) <= input(33);
output(0, 162) <= input(16);
output(0, 163) <= input(17);
output(0, 164) <= input(18);
output(0, 165) <= input(19);
output(0, 166) <= input(20);
output(0, 167) <= input(21);
output(0, 168) <= input(22);
output(0, 169) <= input(23);
output(0, 170) <= input(24);
output(0, 171) <= input(25);
output(0, 172) <= input(26);
output(0, 173) <= input(27);
output(0, 174) <= input(28);
output(0, 175) <= input(29);
output(0, 176) <= input(35);
output(0, 177) <= input(33);
output(0, 178) <= input(16);
output(0, 179) <= input(17);
output(0, 180) <= input(18);
output(0, 181) <= input(19);
output(0, 182) <= input(20);
output(0, 183) <= input(21);
output(0, 184) <= input(22);
output(0, 185) <= input(23);
output(0, 186) <= input(24);
output(0, 187) <= input(25);
output(0, 188) <= input(26);
output(0, 189) <= input(27);
output(0, 190) <= input(28);
output(0, 191) <= input(29);
output(0, 192) <= input(36);
output(0, 193) <= input(34);
output(0, 194) <= input(32);
output(0, 195) <= input(0);
output(0, 196) <= input(1);
output(0, 197) <= input(2);
output(0, 198) <= input(3);
output(0, 199) <= input(4);
output(0, 200) <= input(5);
output(0, 201) <= input(6);
output(0, 202) <= input(7);
output(0, 203) <= input(8);
output(0, 204) <= input(9);
output(0, 205) <= input(10);
output(0, 206) <= input(11);
output(0, 207) <= input(12);
output(0, 208) <= input(36);
output(0, 209) <= input(34);
output(0, 210) <= input(32);
output(0, 211) <= input(0);
output(0, 212) <= input(1);
output(0, 213) <= input(2);
output(0, 214) <= input(3);
output(0, 215) <= input(4);
output(0, 216) <= input(5);
output(0, 217) <= input(6);
output(0, 218) <= input(7);
output(0, 219) <= input(8);
output(0, 220) <= input(9);
output(0, 221) <= input(10);
output(0, 222) <= input(11);
output(0, 223) <= input(12);
output(0, 224) <= input(37);
output(0, 225) <= input(35);
output(0, 226) <= input(33);
output(0, 227) <= input(16);
output(0, 228) <= input(17);
output(0, 229) <= input(18);
output(0, 230) <= input(19);
output(0, 231) <= input(20);
output(0, 232) <= input(21);
output(0, 233) <= input(22);
output(0, 234) <= input(23);
output(0, 235) <= input(24);
output(0, 236) <= input(25);
output(0, 237) <= input(26);
output(0, 238) <= input(27);
output(0, 239) <= input(28);
output(0, 240) <= input(37);
output(0, 241) <= input(35);
output(0, 242) <= input(33);
output(0, 243) <= input(16);
output(0, 244) <= input(17);
output(0, 245) <= input(18);
output(0, 246) <= input(19);
output(0, 247) <= input(20);
output(0, 248) <= input(21);
output(0, 249) <= input(22);
output(0, 250) <= input(23);
output(0, 251) <= input(24);
output(0, 252) <= input(25);
output(0, 253) <= input(26);
output(0, 254) <= input(27);
output(0, 255) <= input(28);
output(1, 0) <= input(1);
output(1, 1) <= input(2);
output(1, 2) <= input(3);
output(1, 3) <= input(4);
output(1, 4) <= input(5);
output(1, 5) <= input(6);
output(1, 6) <= input(7);
output(1, 7) <= input(8);
output(1, 8) <= input(9);
output(1, 9) <= input(10);
output(1, 10) <= input(11);
output(1, 11) <= input(12);
output(1, 12) <= input(13);
output(1, 13) <= input(14);
output(1, 14) <= input(15);
output(1, 15) <= input(38);
output(1, 16) <= input(1);
output(1, 17) <= input(2);
output(1, 18) <= input(3);
output(1, 19) <= input(4);
output(1, 20) <= input(5);
output(1, 21) <= input(6);
output(1, 22) <= input(7);
output(1, 23) <= input(8);
output(1, 24) <= input(9);
output(1, 25) <= input(10);
output(1, 26) <= input(11);
output(1, 27) <= input(12);
output(1, 28) <= input(13);
output(1, 29) <= input(14);
output(1, 30) <= input(15);
output(1, 31) <= input(38);
output(1, 32) <= input(17);
output(1, 33) <= input(18);
output(1, 34) <= input(19);
output(1, 35) <= input(20);
output(1, 36) <= input(21);
output(1, 37) <= input(22);
output(1, 38) <= input(23);
output(1, 39) <= input(24);
output(1, 40) <= input(25);
output(1, 41) <= input(26);
output(1, 42) <= input(27);
output(1, 43) <= input(28);
output(1, 44) <= input(29);
output(1, 45) <= input(30);
output(1, 46) <= input(31);
output(1, 47) <= input(39);
output(1, 48) <= input(17);
output(1, 49) <= input(18);
output(1, 50) <= input(19);
output(1, 51) <= input(20);
output(1, 52) <= input(21);
output(1, 53) <= input(22);
output(1, 54) <= input(23);
output(1, 55) <= input(24);
output(1, 56) <= input(25);
output(1, 57) <= input(26);
output(1, 58) <= input(27);
output(1, 59) <= input(28);
output(1, 60) <= input(29);
output(1, 61) <= input(30);
output(1, 62) <= input(31);
output(1, 63) <= input(39);
output(1, 64) <= input(17);
output(1, 65) <= input(18);
output(1, 66) <= input(19);
output(1, 67) <= input(20);
output(1, 68) <= input(21);
output(1, 69) <= input(22);
output(1, 70) <= input(23);
output(1, 71) <= input(24);
output(1, 72) <= input(25);
output(1, 73) <= input(26);
output(1, 74) <= input(27);
output(1, 75) <= input(28);
output(1, 76) <= input(29);
output(1, 77) <= input(30);
output(1, 78) <= input(31);
output(1, 79) <= input(39);
output(1, 80) <= input(0);
output(1, 81) <= input(1);
output(1, 82) <= input(2);
output(1, 83) <= input(3);
output(1, 84) <= input(4);
output(1, 85) <= input(5);
output(1, 86) <= input(6);
output(1, 87) <= input(7);
output(1, 88) <= input(8);
output(1, 89) <= input(9);
output(1, 90) <= input(10);
output(1, 91) <= input(11);
output(1, 92) <= input(12);
output(1, 93) <= input(13);
output(1, 94) <= input(14);
output(1, 95) <= input(15);
output(1, 96) <= input(0);
output(1, 97) <= input(1);
output(1, 98) <= input(2);
output(1, 99) <= input(3);
output(1, 100) <= input(4);
output(1, 101) <= input(5);
output(1, 102) <= input(6);
output(1, 103) <= input(7);
output(1, 104) <= input(8);
output(1, 105) <= input(9);
output(1, 106) <= input(10);
output(1, 107) <= input(11);
output(1, 108) <= input(12);
output(1, 109) <= input(13);
output(1, 110) <= input(14);
output(1, 111) <= input(15);
output(1, 112) <= input(0);
output(1, 113) <= input(1);
output(1, 114) <= input(2);
output(1, 115) <= input(3);
output(1, 116) <= input(4);
output(1, 117) <= input(5);
output(1, 118) <= input(6);
output(1, 119) <= input(7);
output(1, 120) <= input(8);
output(1, 121) <= input(9);
output(1, 122) <= input(10);
output(1, 123) <= input(11);
output(1, 124) <= input(12);
output(1, 125) <= input(13);
output(1, 126) <= input(14);
output(1, 127) <= input(15);
output(1, 128) <= input(16);
output(1, 129) <= input(17);
output(1, 130) <= input(18);
output(1, 131) <= input(19);
output(1, 132) <= input(20);
output(1, 133) <= input(21);
output(1, 134) <= input(22);
output(1, 135) <= input(23);
output(1, 136) <= input(24);
output(1, 137) <= input(25);
output(1, 138) <= input(26);
output(1, 139) <= input(27);
output(1, 140) <= input(28);
output(1, 141) <= input(29);
output(1, 142) <= input(30);
output(1, 143) <= input(31);
output(1, 144) <= input(16);
output(1, 145) <= input(17);
output(1, 146) <= input(18);
output(1, 147) <= input(19);
output(1, 148) <= input(20);
output(1, 149) <= input(21);
output(1, 150) <= input(22);
output(1, 151) <= input(23);
output(1, 152) <= input(24);
output(1, 153) <= input(25);
output(1, 154) <= input(26);
output(1, 155) <= input(27);
output(1, 156) <= input(28);
output(1, 157) <= input(29);
output(1, 158) <= input(30);
output(1, 159) <= input(31);
output(1, 160) <= input(32);
output(1, 161) <= input(0);
output(1, 162) <= input(1);
output(1, 163) <= input(2);
output(1, 164) <= input(3);
output(1, 165) <= input(4);
output(1, 166) <= input(5);
output(1, 167) <= input(6);
output(1, 168) <= input(7);
output(1, 169) <= input(8);
output(1, 170) <= input(9);
output(1, 171) <= input(10);
output(1, 172) <= input(11);
output(1, 173) <= input(12);
output(1, 174) <= input(13);
output(1, 175) <= input(14);
output(1, 176) <= input(32);
output(1, 177) <= input(0);
output(1, 178) <= input(1);
output(1, 179) <= input(2);
output(1, 180) <= input(3);
output(1, 181) <= input(4);
output(1, 182) <= input(5);
output(1, 183) <= input(6);
output(1, 184) <= input(7);
output(1, 185) <= input(8);
output(1, 186) <= input(9);
output(1, 187) <= input(10);
output(1, 188) <= input(11);
output(1, 189) <= input(12);
output(1, 190) <= input(13);
output(1, 191) <= input(14);
output(1, 192) <= input(32);
output(1, 193) <= input(0);
output(1, 194) <= input(1);
output(1, 195) <= input(2);
output(1, 196) <= input(3);
output(1, 197) <= input(4);
output(1, 198) <= input(5);
output(1, 199) <= input(6);
output(1, 200) <= input(7);
output(1, 201) <= input(8);
output(1, 202) <= input(9);
output(1, 203) <= input(10);
output(1, 204) <= input(11);
output(1, 205) <= input(12);
output(1, 206) <= input(13);
output(1, 207) <= input(14);
output(1, 208) <= input(33);
output(1, 209) <= input(16);
output(1, 210) <= input(17);
output(1, 211) <= input(18);
output(1, 212) <= input(19);
output(1, 213) <= input(20);
output(1, 214) <= input(21);
output(1, 215) <= input(22);
output(1, 216) <= input(23);
output(1, 217) <= input(24);
output(1, 218) <= input(25);
output(1, 219) <= input(26);
output(1, 220) <= input(27);
output(1, 221) <= input(28);
output(1, 222) <= input(29);
output(1, 223) <= input(30);
output(1, 224) <= input(33);
output(1, 225) <= input(16);
output(1, 226) <= input(17);
output(1, 227) <= input(18);
output(1, 228) <= input(19);
output(1, 229) <= input(20);
output(1, 230) <= input(21);
output(1, 231) <= input(22);
output(1, 232) <= input(23);
output(1, 233) <= input(24);
output(1, 234) <= input(25);
output(1, 235) <= input(26);
output(1, 236) <= input(27);
output(1, 237) <= input(28);
output(1, 238) <= input(29);
output(1, 239) <= input(30);
output(1, 240) <= input(33);
output(1, 241) <= input(16);
output(1, 242) <= input(17);
output(1, 243) <= input(18);
output(1, 244) <= input(19);
output(1, 245) <= input(20);
output(1, 246) <= input(21);
output(1, 247) <= input(22);
output(1, 248) <= input(23);
output(1, 249) <= input(24);
output(1, 250) <= input(25);
output(1, 251) <= input(26);
output(1, 252) <= input(27);
output(1, 253) <= input(28);
output(1, 254) <= input(29);
output(1, 255) <= input(30);
output(2, 0) <= input(2);
output(2, 1) <= input(3);
output(2, 2) <= input(4);
output(2, 3) <= input(5);
output(2, 4) <= input(6);
output(2, 5) <= input(7);
output(2, 6) <= input(8);
output(2, 7) <= input(9);
output(2, 8) <= input(10);
output(2, 9) <= input(11);
output(2, 10) <= input(12);
output(2, 11) <= input(13);
output(2, 12) <= input(14);
output(2, 13) <= input(15);
output(2, 14) <= input(38);
output(2, 15) <= input(40);
output(2, 16) <= input(2);
output(2, 17) <= input(3);
output(2, 18) <= input(4);
output(2, 19) <= input(5);
output(2, 20) <= input(6);
output(2, 21) <= input(7);
output(2, 22) <= input(8);
output(2, 23) <= input(9);
output(2, 24) <= input(10);
output(2, 25) <= input(11);
output(2, 26) <= input(12);
output(2, 27) <= input(13);
output(2, 28) <= input(14);
output(2, 29) <= input(15);
output(2, 30) <= input(38);
output(2, 31) <= input(40);
output(2, 32) <= input(2);
output(2, 33) <= input(3);
output(2, 34) <= input(4);
output(2, 35) <= input(5);
output(2, 36) <= input(6);
output(2, 37) <= input(7);
output(2, 38) <= input(8);
output(2, 39) <= input(9);
output(2, 40) <= input(10);
output(2, 41) <= input(11);
output(2, 42) <= input(12);
output(2, 43) <= input(13);
output(2, 44) <= input(14);
output(2, 45) <= input(15);
output(2, 46) <= input(38);
output(2, 47) <= input(40);
output(2, 48) <= input(2);
output(2, 49) <= input(3);
output(2, 50) <= input(4);
output(2, 51) <= input(5);
output(2, 52) <= input(6);
output(2, 53) <= input(7);
output(2, 54) <= input(8);
output(2, 55) <= input(9);
output(2, 56) <= input(10);
output(2, 57) <= input(11);
output(2, 58) <= input(12);
output(2, 59) <= input(13);
output(2, 60) <= input(14);
output(2, 61) <= input(15);
output(2, 62) <= input(38);
output(2, 63) <= input(40);
output(2, 64) <= input(18);
output(2, 65) <= input(19);
output(2, 66) <= input(20);
output(2, 67) <= input(21);
output(2, 68) <= input(22);
output(2, 69) <= input(23);
output(2, 70) <= input(24);
output(2, 71) <= input(25);
output(2, 72) <= input(26);
output(2, 73) <= input(27);
output(2, 74) <= input(28);
output(2, 75) <= input(29);
output(2, 76) <= input(30);
output(2, 77) <= input(31);
output(2, 78) <= input(39);
output(2, 79) <= input(41);
output(2, 80) <= input(18);
output(2, 81) <= input(19);
output(2, 82) <= input(20);
output(2, 83) <= input(21);
output(2, 84) <= input(22);
output(2, 85) <= input(23);
output(2, 86) <= input(24);
output(2, 87) <= input(25);
output(2, 88) <= input(26);
output(2, 89) <= input(27);
output(2, 90) <= input(28);
output(2, 91) <= input(29);
output(2, 92) <= input(30);
output(2, 93) <= input(31);
output(2, 94) <= input(39);
output(2, 95) <= input(41);
output(2, 96) <= input(18);
output(2, 97) <= input(19);
output(2, 98) <= input(20);
output(2, 99) <= input(21);
output(2, 100) <= input(22);
output(2, 101) <= input(23);
output(2, 102) <= input(24);
output(2, 103) <= input(25);
output(2, 104) <= input(26);
output(2, 105) <= input(27);
output(2, 106) <= input(28);
output(2, 107) <= input(29);
output(2, 108) <= input(30);
output(2, 109) <= input(31);
output(2, 110) <= input(39);
output(2, 111) <= input(41);
output(2, 112) <= input(18);
output(2, 113) <= input(19);
output(2, 114) <= input(20);
output(2, 115) <= input(21);
output(2, 116) <= input(22);
output(2, 117) <= input(23);
output(2, 118) <= input(24);
output(2, 119) <= input(25);
output(2, 120) <= input(26);
output(2, 121) <= input(27);
output(2, 122) <= input(28);
output(2, 123) <= input(29);
output(2, 124) <= input(30);
output(2, 125) <= input(31);
output(2, 126) <= input(39);
output(2, 127) <= input(41);
output(2, 128) <= input(1);
output(2, 129) <= input(2);
output(2, 130) <= input(3);
output(2, 131) <= input(4);
output(2, 132) <= input(5);
output(2, 133) <= input(6);
output(2, 134) <= input(7);
output(2, 135) <= input(8);
output(2, 136) <= input(9);
output(2, 137) <= input(10);
output(2, 138) <= input(11);
output(2, 139) <= input(12);
output(2, 140) <= input(13);
output(2, 141) <= input(14);
output(2, 142) <= input(15);
output(2, 143) <= input(38);
output(2, 144) <= input(1);
output(2, 145) <= input(2);
output(2, 146) <= input(3);
output(2, 147) <= input(4);
output(2, 148) <= input(5);
output(2, 149) <= input(6);
output(2, 150) <= input(7);
output(2, 151) <= input(8);
output(2, 152) <= input(9);
output(2, 153) <= input(10);
output(2, 154) <= input(11);
output(2, 155) <= input(12);
output(2, 156) <= input(13);
output(2, 157) <= input(14);
output(2, 158) <= input(15);
output(2, 159) <= input(38);
output(2, 160) <= input(1);
output(2, 161) <= input(2);
output(2, 162) <= input(3);
output(2, 163) <= input(4);
output(2, 164) <= input(5);
output(2, 165) <= input(6);
output(2, 166) <= input(7);
output(2, 167) <= input(8);
output(2, 168) <= input(9);
output(2, 169) <= input(10);
output(2, 170) <= input(11);
output(2, 171) <= input(12);
output(2, 172) <= input(13);
output(2, 173) <= input(14);
output(2, 174) <= input(15);
output(2, 175) <= input(38);
output(2, 176) <= input(1);
output(2, 177) <= input(2);
output(2, 178) <= input(3);
output(2, 179) <= input(4);
output(2, 180) <= input(5);
output(2, 181) <= input(6);
output(2, 182) <= input(7);
output(2, 183) <= input(8);
output(2, 184) <= input(9);
output(2, 185) <= input(10);
output(2, 186) <= input(11);
output(2, 187) <= input(12);
output(2, 188) <= input(13);
output(2, 189) <= input(14);
output(2, 190) <= input(15);
output(2, 191) <= input(38);
output(2, 192) <= input(17);
output(2, 193) <= input(18);
output(2, 194) <= input(19);
output(2, 195) <= input(20);
output(2, 196) <= input(21);
output(2, 197) <= input(22);
output(2, 198) <= input(23);
output(2, 199) <= input(24);
output(2, 200) <= input(25);
output(2, 201) <= input(26);
output(2, 202) <= input(27);
output(2, 203) <= input(28);
output(2, 204) <= input(29);
output(2, 205) <= input(30);
output(2, 206) <= input(31);
output(2, 207) <= input(39);
output(2, 208) <= input(17);
output(2, 209) <= input(18);
output(2, 210) <= input(19);
output(2, 211) <= input(20);
output(2, 212) <= input(21);
output(2, 213) <= input(22);
output(2, 214) <= input(23);
output(2, 215) <= input(24);
output(2, 216) <= input(25);
output(2, 217) <= input(26);
output(2, 218) <= input(27);
output(2, 219) <= input(28);
output(2, 220) <= input(29);
output(2, 221) <= input(30);
output(2, 222) <= input(31);
output(2, 223) <= input(39);
output(2, 224) <= input(17);
output(2, 225) <= input(18);
output(2, 226) <= input(19);
output(2, 227) <= input(20);
output(2, 228) <= input(21);
output(2, 229) <= input(22);
output(2, 230) <= input(23);
output(2, 231) <= input(24);
output(2, 232) <= input(25);
output(2, 233) <= input(26);
output(2, 234) <= input(27);
output(2, 235) <= input(28);
output(2, 236) <= input(29);
output(2, 237) <= input(30);
output(2, 238) <= input(31);
output(2, 239) <= input(39);
output(2, 240) <= input(17);
output(2, 241) <= input(18);
output(2, 242) <= input(19);
output(2, 243) <= input(20);
output(2, 244) <= input(21);
output(2, 245) <= input(22);
output(2, 246) <= input(23);
output(2, 247) <= input(24);
output(2, 248) <= input(25);
output(2, 249) <= input(26);
output(2, 250) <= input(27);
output(2, 251) <= input(28);
output(2, 252) <= input(29);
output(2, 253) <= input(30);
output(2, 254) <= input(31);
output(2, 255) <= input(39);
when "1101" =>
output(0, 0) <= input(0);
output(0, 1) <= input(1);
output(0, 2) <= input(2);
output(0, 3) <= input(3);
output(0, 4) <= input(4);
output(0, 5) <= input(5);
output(0, 6) <= input(6);
output(0, 7) <= input(7);
output(0, 8) <= input(8);
output(0, 9) <= input(9);
output(0, 10) <= input(10);
output(0, 11) <= input(11);
output(0, 12) <= input(12);
output(0, 13) <= input(13);
output(0, 14) <= input(14);
output(0, 15) <= input(15);
output(0, 16) <= input(0);
output(0, 17) <= input(1);
output(0, 18) <= input(2);
output(0, 19) <= input(3);
output(0, 20) <= input(4);
output(0, 21) <= input(5);
output(0, 22) <= input(6);
output(0, 23) <= input(7);
output(0, 24) <= input(8);
output(0, 25) <= input(9);
output(0, 26) <= input(10);
output(0, 27) <= input(11);
output(0, 28) <= input(12);
output(0, 29) <= input(13);
output(0, 30) <= input(14);
output(0, 31) <= input(15);
output(0, 32) <= input(0);
output(0, 33) <= input(1);
output(0, 34) <= input(2);
output(0, 35) <= input(3);
output(0, 36) <= input(4);
output(0, 37) <= input(5);
output(0, 38) <= input(6);
output(0, 39) <= input(7);
output(0, 40) <= input(8);
output(0, 41) <= input(9);
output(0, 42) <= input(10);
output(0, 43) <= input(11);
output(0, 44) <= input(12);
output(0, 45) <= input(13);
output(0, 46) <= input(14);
output(0, 47) <= input(15);
output(0, 48) <= input(0);
output(0, 49) <= input(1);
output(0, 50) <= input(2);
output(0, 51) <= input(3);
output(0, 52) <= input(4);
output(0, 53) <= input(5);
output(0, 54) <= input(6);
output(0, 55) <= input(7);
output(0, 56) <= input(8);
output(0, 57) <= input(9);
output(0, 58) <= input(10);
output(0, 59) <= input(11);
output(0, 60) <= input(12);
output(0, 61) <= input(13);
output(0, 62) <= input(14);
output(0, 63) <= input(15);
output(0, 64) <= input(0);
output(0, 65) <= input(1);
output(0, 66) <= input(2);
output(0, 67) <= input(3);
output(0, 68) <= input(4);
output(0, 69) <= input(5);
output(0, 70) <= input(6);
output(0, 71) <= input(7);
output(0, 72) <= input(8);
output(0, 73) <= input(9);
output(0, 74) <= input(10);
output(0, 75) <= input(11);
output(0, 76) <= input(12);
output(0, 77) <= input(13);
output(0, 78) <= input(14);
output(0, 79) <= input(15);
output(0, 80) <= input(16);
output(0, 81) <= input(17);
output(0, 82) <= input(18);
output(0, 83) <= input(19);
output(0, 84) <= input(20);
output(0, 85) <= input(21);
output(0, 86) <= input(22);
output(0, 87) <= input(23);
output(0, 88) <= input(24);
output(0, 89) <= input(25);
output(0, 90) <= input(26);
output(0, 91) <= input(27);
output(0, 92) <= input(28);
output(0, 93) <= input(29);
output(0, 94) <= input(30);
output(0, 95) <= input(31);
output(0, 96) <= input(16);
output(0, 97) <= input(17);
output(0, 98) <= input(18);
output(0, 99) <= input(19);
output(0, 100) <= input(20);
output(0, 101) <= input(21);
output(0, 102) <= input(22);
output(0, 103) <= input(23);
output(0, 104) <= input(24);
output(0, 105) <= input(25);
output(0, 106) <= input(26);
output(0, 107) <= input(27);
output(0, 108) <= input(28);
output(0, 109) <= input(29);
output(0, 110) <= input(30);
output(0, 111) <= input(31);
output(0, 112) <= input(16);
output(0, 113) <= input(17);
output(0, 114) <= input(18);
output(0, 115) <= input(19);
output(0, 116) <= input(20);
output(0, 117) <= input(21);
output(0, 118) <= input(22);
output(0, 119) <= input(23);
output(0, 120) <= input(24);
output(0, 121) <= input(25);
output(0, 122) <= input(26);
output(0, 123) <= input(27);
output(0, 124) <= input(28);
output(0, 125) <= input(29);
output(0, 126) <= input(30);
output(0, 127) <= input(31);
output(0, 128) <= input(16);
output(0, 129) <= input(17);
output(0, 130) <= input(18);
output(0, 131) <= input(19);
output(0, 132) <= input(20);
output(0, 133) <= input(21);
output(0, 134) <= input(22);
output(0, 135) <= input(23);
output(0, 136) <= input(24);
output(0, 137) <= input(25);
output(0, 138) <= input(26);
output(0, 139) <= input(27);
output(0, 140) <= input(28);
output(0, 141) <= input(29);
output(0, 142) <= input(30);
output(0, 143) <= input(31);
output(0, 144) <= input(16);
output(0, 145) <= input(17);
output(0, 146) <= input(18);
output(0, 147) <= input(19);
output(0, 148) <= input(20);
output(0, 149) <= input(21);
output(0, 150) <= input(22);
output(0, 151) <= input(23);
output(0, 152) <= input(24);
output(0, 153) <= input(25);
output(0, 154) <= input(26);
output(0, 155) <= input(27);
output(0, 156) <= input(28);
output(0, 157) <= input(29);
output(0, 158) <= input(30);
output(0, 159) <= input(31);
output(0, 160) <= input(32);
output(0, 161) <= input(0);
output(0, 162) <= input(1);
output(0, 163) <= input(2);
output(0, 164) <= input(3);
output(0, 165) <= input(4);
output(0, 166) <= input(5);
output(0, 167) <= input(6);
output(0, 168) <= input(7);
output(0, 169) <= input(8);
output(0, 170) <= input(9);
output(0, 171) <= input(10);
output(0, 172) <= input(11);
output(0, 173) <= input(12);
output(0, 174) <= input(13);
output(0, 175) <= input(14);
output(0, 176) <= input(32);
output(0, 177) <= input(0);
output(0, 178) <= input(1);
output(0, 179) <= input(2);
output(0, 180) <= input(3);
output(0, 181) <= input(4);
output(0, 182) <= input(5);
output(0, 183) <= input(6);
output(0, 184) <= input(7);
output(0, 185) <= input(8);
output(0, 186) <= input(9);
output(0, 187) <= input(10);
output(0, 188) <= input(11);
output(0, 189) <= input(12);
output(0, 190) <= input(13);
output(0, 191) <= input(14);
output(0, 192) <= input(32);
output(0, 193) <= input(0);
output(0, 194) <= input(1);
output(0, 195) <= input(2);
output(0, 196) <= input(3);
output(0, 197) <= input(4);
output(0, 198) <= input(5);
output(0, 199) <= input(6);
output(0, 200) <= input(7);
output(0, 201) <= input(8);
output(0, 202) <= input(9);
output(0, 203) <= input(10);
output(0, 204) <= input(11);
output(0, 205) <= input(12);
output(0, 206) <= input(13);
output(0, 207) <= input(14);
output(0, 208) <= input(32);
output(0, 209) <= input(0);
output(0, 210) <= input(1);
output(0, 211) <= input(2);
output(0, 212) <= input(3);
output(0, 213) <= input(4);
output(0, 214) <= input(5);
output(0, 215) <= input(6);
output(0, 216) <= input(7);
output(0, 217) <= input(8);
output(0, 218) <= input(9);
output(0, 219) <= input(10);
output(0, 220) <= input(11);
output(0, 221) <= input(12);
output(0, 222) <= input(13);
output(0, 223) <= input(14);
output(0, 224) <= input(32);
output(0, 225) <= input(0);
output(0, 226) <= input(1);
output(0, 227) <= input(2);
output(0, 228) <= input(3);
output(0, 229) <= input(4);
output(0, 230) <= input(5);
output(0, 231) <= input(6);
output(0, 232) <= input(7);
output(0, 233) <= input(8);
output(0, 234) <= input(9);
output(0, 235) <= input(10);
output(0, 236) <= input(11);
output(0, 237) <= input(12);
output(0, 238) <= input(13);
output(0, 239) <= input(14);
output(0, 240) <= input(32);
output(0, 241) <= input(0);
output(0, 242) <= input(1);
output(0, 243) <= input(2);
output(0, 244) <= input(3);
output(0, 245) <= input(4);
output(0, 246) <= input(5);
output(0, 247) <= input(6);
output(0, 248) <= input(7);
output(0, 249) <= input(8);
output(0, 250) <= input(9);
output(0, 251) <= input(10);
output(0, 252) <= input(11);
output(0, 253) <= input(12);
output(0, 254) <= input(13);
output(0, 255) <= input(14);
output(1, 0) <= input(17);
output(1, 1) <= input(18);
output(1, 2) <= input(19);
output(1, 3) <= input(20);
output(1, 4) <= input(21);
output(1, 5) <= input(22);
output(1, 6) <= input(23);
output(1, 7) <= input(24);
output(1, 8) <= input(25);
output(1, 9) <= input(26);
output(1, 10) <= input(27);
output(1, 11) <= input(28);
output(1, 12) <= input(29);
output(1, 13) <= input(30);
output(1, 14) <= input(31);
output(1, 15) <= input(33);
output(1, 16) <= input(17);
output(1, 17) <= input(18);
output(1, 18) <= input(19);
output(1, 19) <= input(20);
output(1, 20) <= input(21);
output(1, 21) <= input(22);
output(1, 22) <= input(23);
output(1, 23) <= input(24);
output(1, 24) <= input(25);
output(1, 25) <= input(26);
output(1, 26) <= input(27);
output(1, 27) <= input(28);
output(1, 28) <= input(29);
output(1, 29) <= input(30);
output(1, 30) <= input(31);
output(1, 31) <= input(33);
output(1, 32) <= input(17);
output(1, 33) <= input(18);
output(1, 34) <= input(19);
output(1, 35) <= input(20);
output(1, 36) <= input(21);
output(1, 37) <= input(22);
output(1, 38) <= input(23);
output(1, 39) <= input(24);
output(1, 40) <= input(25);
output(1, 41) <= input(26);
output(1, 42) <= input(27);
output(1, 43) <= input(28);
output(1, 44) <= input(29);
output(1, 45) <= input(30);
output(1, 46) <= input(31);
output(1, 47) <= input(33);
output(1, 48) <= input(17);
output(1, 49) <= input(18);
output(1, 50) <= input(19);
output(1, 51) <= input(20);
output(1, 52) <= input(21);
output(1, 53) <= input(22);
output(1, 54) <= input(23);
output(1, 55) <= input(24);
output(1, 56) <= input(25);
output(1, 57) <= input(26);
output(1, 58) <= input(27);
output(1, 59) <= input(28);
output(1, 60) <= input(29);
output(1, 61) <= input(30);
output(1, 62) <= input(31);
output(1, 63) <= input(33);
output(1, 64) <= input(17);
output(1, 65) <= input(18);
output(1, 66) <= input(19);
output(1, 67) <= input(20);
output(1, 68) <= input(21);
output(1, 69) <= input(22);
output(1, 70) <= input(23);
output(1, 71) <= input(24);
output(1, 72) <= input(25);
output(1, 73) <= input(26);
output(1, 74) <= input(27);
output(1, 75) <= input(28);
output(1, 76) <= input(29);
output(1, 77) <= input(30);
output(1, 78) <= input(31);
output(1, 79) <= input(33);
output(1, 80) <= input(17);
output(1, 81) <= input(18);
output(1, 82) <= input(19);
output(1, 83) <= input(20);
output(1, 84) <= input(21);
output(1, 85) <= input(22);
output(1, 86) <= input(23);
output(1, 87) <= input(24);
output(1, 88) <= input(25);
output(1, 89) <= input(26);
output(1, 90) <= input(27);
output(1, 91) <= input(28);
output(1, 92) <= input(29);
output(1, 93) <= input(30);
output(1, 94) <= input(31);
output(1, 95) <= input(33);
output(1, 96) <= input(17);
output(1, 97) <= input(18);
output(1, 98) <= input(19);
output(1, 99) <= input(20);
output(1, 100) <= input(21);
output(1, 101) <= input(22);
output(1, 102) <= input(23);
output(1, 103) <= input(24);
output(1, 104) <= input(25);
output(1, 105) <= input(26);
output(1, 106) <= input(27);
output(1, 107) <= input(28);
output(1, 108) <= input(29);
output(1, 109) <= input(30);
output(1, 110) <= input(31);
output(1, 111) <= input(33);
output(1, 112) <= input(17);
output(1, 113) <= input(18);
output(1, 114) <= input(19);
output(1, 115) <= input(20);
output(1, 116) <= input(21);
output(1, 117) <= input(22);
output(1, 118) <= input(23);
output(1, 119) <= input(24);
output(1, 120) <= input(25);
output(1, 121) <= input(26);
output(1, 122) <= input(27);
output(1, 123) <= input(28);
output(1, 124) <= input(29);
output(1, 125) <= input(30);
output(1, 126) <= input(31);
output(1, 127) <= input(33);
output(1, 128) <= input(0);
output(1, 129) <= input(1);
output(1, 130) <= input(2);
output(1, 131) <= input(3);
output(1, 132) <= input(4);
output(1, 133) <= input(5);
output(1, 134) <= input(6);
output(1, 135) <= input(7);
output(1, 136) <= input(8);
output(1, 137) <= input(9);
output(1, 138) <= input(10);
output(1, 139) <= input(11);
output(1, 140) <= input(12);
output(1, 141) <= input(13);
output(1, 142) <= input(14);
output(1, 143) <= input(15);
output(1, 144) <= input(0);
output(1, 145) <= input(1);
output(1, 146) <= input(2);
output(1, 147) <= input(3);
output(1, 148) <= input(4);
output(1, 149) <= input(5);
output(1, 150) <= input(6);
output(1, 151) <= input(7);
output(1, 152) <= input(8);
output(1, 153) <= input(9);
output(1, 154) <= input(10);
output(1, 155) <= input(11);
output(1, 156) <= input(12);
output(1, 157) <= input(13);
output(1, 158) <= input(14);
output(1, 159) <= input(15);
output(1, 160) <= input(0);
output(1, 161) <= input(1);
output(1, 162) <= input(2);
output(1, 163) <= input(3);
output(1, 164) <= input(4);
output(1, 165) <= input(5);
output(1, 166) <= input(6);
output(1, 167) <= input(7);
output(1, 168) <= input(8);
output(1, 169) <= input(9);
output(1, 170) <= input(10);
output(1, 171) <= input(11);
output(1, 172) <= input(12);
output(1, 173) <= input(13);
output(1, 174) <= input(14);
output(1, 175) <= input(15);
output(1, 176) <= input(0);
output(1, 177) <= input(1);
output(1, 178) <= input(2);
output(1, 179) <= input(3);
output(1, 180) <= input(4);
output(1, 181) <= input(5);
output(1, 182) <= input(6);
output(1, 183) <= input(7);
output(1, 184) <= input(8);
output(1, 185) <= input(9);
output(1, 186) <= input(10);
output(1, 187) <= input(11);
output(1, 188) <= input(12);
output(1, 189) <= input(13);
output(1, 190) <= input(14);
output(1, 191) <= input(15);
output(1, 192) <= input(0);
output(1, 193) <= input(1);
output(1, 194) <= input(2);
output(1, 195) <= input(3);
output(1, 196) <= input(4);
output(1, 197) <= input(5);
output(1, 198) <= input(6);
output(1, 199) <= input(7);
output(1, 200) <= input(8);
output(1, 201) <= input(9);
output(1, 202) <= input(10);
output(1, 203) <= input(11);
output(1, 204) <= input(12);
output(1, 205) <= input(13);
output(1, 206) <= input(14);
output(1, 207) <= input(15);
output(1, 208) <= input(0);
output(1, 209) <= input(1);
output(1, 210) <= input(2);
output(1, 211) <= input(3);
output(1, 212) <= input(4);
output(1, 213) <= input(5);
output(1, 214) <= input(6);
output(1, 215) <= input(7);
output(1, 216) <= input(8);
output(1, 217) <= input(9);
output(1, 218) <= input(10);
output(1, 219) <= input(11);
output(1, 220) <= input(12);
output(1, 221) <= input(13);
output(1, 222) <= input(14);
output(1, 223) <= input(15);
output(1, 224) <= input(0);
output(1, 225) <= input(1);
output(1, 226) <= input(2);
output(1, 227) <= input(3);
output(1, 228) <= input(4);
output(1, 229) <= input(5);
output(1, 230) <= input(6);
output(1, 231) <= input(7);
output(1, 232) <= input(8);
output(1, 233) <= input(9);
output(1, 234) <= input(10);
output(1, 235) <= input(11);
output(1, 236) <= input(12);
output(1, 237) <= input(13);
output(1, 238) <= input(14);
output(1, 239) <= input(15);
output(1, 240) <= input(0);
output(1, 241) <= input(1);
output(1, 242) <= input(2);
output(1, 243) <= input(3);
output(1, 244) <= input(4);
output(1, 245) <= input(5);
output(1, 246) <= input(6);
output(1, 247) <= input(7);
output(1, 248) <= input(8);
output(1, 249) <= input(9);
output(1, 250) <= input(10);
output(1, 251) <= input(11);
output(1, 252) <= input(12);
output(1, 253) <= input(13);
output(1, 254) <= input(14);
output(1, 255) <= input(15);
output(2, 0) <= input(1);
output(2, 1) <= input(2);
output(2, 2) <= input(3);
output(2, 3) <= input(4);
output(2, 4) <= input(5);
output(2, 5) <= input(6);
output(2, 6) <= input(7);
output(2, 7) <= input(8);
output(2, 8) <= input(9);
output(2, 9) <= input(10);
output(2, 10) <= input(11);
output(2, 11) <= input(12);
output(2, 12) <= input(13);
output(2, 13) <= input(14);
output(2, 14) <= input(15);
output(2, 15) <= input(34);
output(2, 16) <= input(1);
output(2, 17) <= input(2);
output(2, 18) <= input(3);
output(2, 19) <= input(4);
output(2, 20) <= input(5);
output(2, 21) <= input(6);
output(2, 22) <= input(7);
output(2, 23) <= input(8);
output(2, 24) <= input(9);
output(2, 25) <= input(10);
output(2, 26) <= input(11);
output(2, 27) <= input(12);
output(2, 28) <= input(13);
output(2, 29) <= input(14);
output(2, 30) <= input(15);
output(2, 31) <= input(34);
output(2, 32) <= input(1);
output(2, 33) <= input(2);
output(2, 34) <= input(3);
output(2, 35) <= input(4);
output(2, 36) <= input(5);
output(2, 37) <= input(6);
output(2, 38) <= input(7);
output(2, 39) <= input(8);
output(2, 40) <= input(9);
output(2, 41) <= input(10);
output(2, 42) <= input(11);
output(2, 43) <= input(12);
output(2, 44) <= input(13);
output(2, 45) <= input(14);
output(2, 46) <= input(15);
output(2, 47) <= input(34);
output(2, 48) <= input(1);
output(2, 49) <= input(2);
output(2, 50) <= input(3);
output(2, 51) <= input(4);
output(2, 52) <= input(5);
output(2, 53) <= input(6);
output(2, 54) <= input(7);
output(2, 55) <= input(8);
output(2, 56) <= input(9);
output(2, 57) <= input(10);
output(2, 58) <= input(11);
output(2, 59) <= input(12);
output(2, 60) <= input(13);
output(2, 61) <= input(14);
output(2, 62) <= input(15);
output(2, 63) <= input(34);
output(2, 64) <= input(1);
output(2, 65) <= input(2);
output(2, 66) <= input(3);
output(2, 67) <= input(4);
output(2, 68) <= input(5);
output(2, 69) <= input(6);
output(2, 70) <= input(7);
output(2, 71) <= input(8);
output(2, 72) <= input(9);
output(2, 73) <= input(10);
output(2, 74) <= input(11);
output(2, 75) <= input(12);
output(2, 76) <= input(13);
output(2, 77) <= input(14);
output(2, 78) <= input(15);
output(2, 79) <= input(34);
output(2, 80) <= input(1);
output(2, 81) <= input(2);
output(2, 82) <= input(3);
output(2, 83) <= input(4);
output(2, 84) <= input(5);
output(2, 85) <= input(6);
output(2, 86) <= input(7);
output(2, 87) <= input(8);
output(2, 88) <= input(9);
output(2, 89) <= input(10);
output(2, 90) <= input(11);
output(2, 91) <= input(12);
output(2, 92) <= input(13);
output(2, 93) <= input(14);
output(2, 94) <= input(15);
output(2, 95) <= input(34);
output(2, 96) <= input(1);
output(2, 97) <= input(2);
output(2, 98) <= input(3);
output(2, 99) <= input(4);
output(2, 100) <= input(5);
output(2, 101) <= input(6);
output(2, 102) <= input(7);
output(2, 103) <= input(8);
output(2, 104) <= input(9);
output(2, 105) <= input(10);
output(2, 106) <= input(11);
output(2, 107) <= input(12);
output(2, 108) <= input(13);
output(2, 109) <= input(14);
output(2, 110) <= input(15);
output(2, 111) <= input(34);
output(2, 112) <= input(1);
output(2, 113) <= input(2);
output(2, 114) <= input(3);
output(2, 115) <= input(4);
output(2, 116) <= input(5);
output(2, 117) <= input(6);
output(2, 118) <= input(7);
output(2, 119) <= input(8);
output(2, 120) <= input(9);
output(2, 121) <= input(10);
output(2, 122) <= input(11);
output(2, 123) <= input(12);
output(2, 124) <= input(13);
output(2, 125) <= input(14);
output(2, 126) <= input(15);
output(2, 127) <= input(34);
output(2, 128) <= input(1);
output(2, 129) <= input(2);
output(2, 130) <= input(3);
output(2, 131) <= input(4);
output(2, 132) <= input(5);
output(2, 133) <= input(6);
output(2, 134) <= input(7);
output(2, 135) <= input(8);
output(2, 136) <= input(9);
output(2, 137) <= input(10);
output(2, 138) <= input(11);
output(2, 139) <= input(12);
output(2, 140) <= input(13);
output(2, 141) <= input(14);
output(2, 142) <= input(15);
output(2, 143) <= input(34);
output(2, 144) <= input(1);
output(2, 145) <= input(2);
output(2, 146) <= input(3);
output(2, 147) <= input(4);
output(2, 148) <= input(5);
output(2, 149) <= input(6);
output(2, 150) <= input(7);
output(2, 151) <= input(8);
output(2, 152) <= input(9);
output(2, 153) <= input(10);
output(2, 154) <= input(11);
output(2, 155) <= input(12);
output(2, 156) <= input(13);
output(2, 157) <= input(14);
output(2, 158) <= input(15);
output(2, 159) <= input(34);
output(2, 160) <= input(1);
output(2, 161) <= input(2);
output(2, 162) <= input(3);
output(2, 163) <= input(4);
output(2, 164) <= input(5);
output(2, 165) <= input(6);
output(2, 166) <= input(7);
output(2, 167) <= input(8);
output(2, 168) <= input(9);
output(2, 169) <= input(10);
output(2, 170) <= input(11);
output(2, 171) <= input(12);
output(2, 172) <= input(13);
output(2, 173) <= input(14);
output(2, 174) <= input(15);
output(2, 175) <= input(34);
output(2, 176) <= input(1);
output(2, 177) <= input(2);
output(2, 178) <= input(3);
output(2, 179) <= input(4);
output(2, 180) <= input(5);
output(2, 181) <= input(6);
output(2, 182) <= input(7);
output(2, 183) <= input(8);
output(2, 184) <= input(9);
output(2, 185) <= input(10);
output(2, 186) <= input(11);
output(2, 187) <= input(12);
output(2, 188) <= input(13);
output(2, 189) <= input(14);
output(2, 190) <= input(15);
output(2, 191) <= input(34);
output(2, 192) <= input(1);
output(2, 193) <= input(2);
output(2, 194) <= input(3);
output(2, 195) <= input(4);
output(2, 196) <= input(5);
output(2, 197) <= input(6);
output(2, 198) <= input(7);
output(2, 199) <= input(8);
output(2, 200) <= input(9);
output(2, 201) <= input(10);
output(2, 202) <= input(11);
output(2, 203) <= input(12);
output(2, 204) <= input(13);
output(2, 205) <= input(14);
output(2, 206) <= input(15);
output(2, 207) <= input(34);
output(2, 208) <= input(1);
output(2, 209) <= input(2);
output(2, 210) <= input(3);
output(2, 211) <= input(4);
output(2, 212) <= input(5);
output(2, 213) <= input(6);
output(2, 214) <= input(7);
output(2, 215) <= input(8);
output(2, 216) <= input(9);
output(2, 217) <= input(10);
output(2, 218) <= input(11);
output(2, 219) <= input(12);
output(2, 220) <= input(13);
output(2, 221) <= input(14);
output(2, 222) <= input(15);
output(2, 223) <= input(34);
output(2, 224) <= input(1);
output(2, 225) <= input(2);
output(2, 226) <= input(3);
output(2, 227) <= input(4);
output(2, 228) <= input(5);
output(2, 229) <= input(6);
output(2, 230) <= input(7);
output(2, 231) <= input(8);
output(2, 232) <= input(9);
output(2, 233) <= input(10);
output(2, 234) <= input(11);
output(2, 235) <= input(12);
output(2, 236) <= input(13);
output(2, 237) <= input(14);
output(2, 238) <= input(15);
output(2, 239) <= input(34);
output(2, 240) <= input(1);
output(2, 241) <= input(2);
output(2, 242) <= input(3);
output(2, 243) <= input(4);
output(2, 244) <= input(5);
output(2, 245) <= input(6);
output(2, 246) <= input(7);
output(2, 247) <= input(8);
output(2, 248) <= input(9);
output(2, 249) <= input(10);
output(2, 250) <= input(11);
output(2, 251) <= input(12);
output(2, 252) <= input(13);
output(2, 253) <= input(14);
output(2, 254) <= input(15);
output(2, 255) <= input(34);
output(3, 0) <= input(2);
output(3, 1) <= input(3);
output(3, 2) <= input(4);
output(3, 3) <= input(5);
output(3, 4) <= input(6);
output(3, 5) <= input(7);
output(3, 6) <= input(8);
output(3, 7) <= input(9);
output(3, 8) <= input(10);
output(3, 9) <= input(11);
output(3, 10) <= input(12);
output(3, 11) <= input(13);
output(3, 12) <= input(14);
output(3, 13) <= input(15);
output(3, 14) <= input(34);
output(3, 15) <= input(35);
output(3, 16) <= input(2);
output(3, 17) <= input(3);
output(3, 18) <= input(4);
output(3, 19) <= input(5);
output(3, 20) <= input(6);
output(3, 21) <= input(7);
output(3, 22) <= input(8);
output(3, 23) <= input(9);
output(3, 24) <= input(10);
output(3, 25) <= input(11);
output(3, 26) <= input(12);
output(3, 27) <= input(13);
output(3, 28) <= input(14);
output(3, 29) <= input(15);
output(3, 30) <= input(34);
output(3, 31) <= input(35);
output(3, 32) <= input(2);
output(3, 33) <= input(3);
output(3, 34) <= input(4);
output(3, 35) <= input(5);
output(3, 36) <= input(6);
output(3, 37) <= input(7);
output(3, 38) <= input(8);
output(3, 39) <= input(9);
output(3, 40) <= input(10);
output(3, 41) <= input(11);
output(3, 42) <= input(12);
output(3, 43) <= input(13);
output(3, 44) <= input(14);
output(3, 45) <= input(15);
output(3, 46) <= input(34);
output(3, 47) <= input(35);
output(3, 48) <= input(2);
output(3, 49) <= input(3);
output(3, 50) <= input(4);
output(3, 51) <= input(5);
output(3, 52) <= input(6);
output(3, 53) <= input(7);
output(3, 54) <= input(8);
output(3, 55) <= input(9);
output(3, 56) <= input(10);
output(3, 57) <= input(11);
output(3, 58) <= input(12);
output(3, 59) <= input(13);
output(3, 60) <= input(14);
output(3, 61) <= input(15);
output(3, 62) <= input(34);
output(3, 63) <= input(35);
output(3, 64) <= input(2);
output(3, 65) <= input(3);
output(3, 66) <= input(4);
output(3, 67) <= input(5);
output(3, 68) <= input(6);
output(3, 69) <= input(7);
output(3, 70) <= input(8);
output(3, 71) <= input(9);
output(3, 72) <= input(10);
output(3, 73) <= input(11);
output(3, 74) <= input(12);
output(3, 75) <= input(13);
output(3, 76) <= input(14);
output(3, 77) <= input(15);
output(3, 78) <= input(34);
output(3, 79) <= input(35);
output(3, 80) <= input(2);
output(3, 81) <= input(3);
output(3, 82) <= input(4);
output(3, 83) <= input(5);
output(3, 84) <= input(6);
output(3, 85) <= input(7);
output(3, 86) <= input(8);
output(3, 87) <= input(9);
output(3, 88) <= input(10);
output(3, 89) <= input(11);
output(3, 90) <= input(12);
output(3, 91) <= input(13);
output(3, 92) <= input(14);
output(3, 93) <= input(15);
output(3, 94) <= input(34);
output(3, 95) <= input(35);
output(3, 96) <= input(2);
output(3, 97) <= input(3);
output(3, 98) <= input(4);
output(3, 99) <= input(5);
output(3, 100) <= input(6);
output(3, 101) <= input(7);
output(3, 102) <= input(8);
output(3, 103) <= input(9);
output(3, 104) <= input(10);
output(3, 105) <= input(11);
output(3, 106) <= input(12);
output(3, 107) <= input(13);
output(3, 108) <= input(14);
output(3, 109) <= input(15);
output(3, 110) <= input(34);
output(3, 111) <= input(35);
output(3, 112) <= input(2);
output(3, 113) <= input(3);
output(3, 114) <= input(4);
output(3, 115) <= input(5);
output(3, 116) <= input(6);
output(3, 117) <= input(7);
output(3, 118) <= input(8);
output(3, 119) <= input(9);
output(3, 120) <= input(10);
output(3, 121) <= input(11);
output(3, 122) <= input(12);
output(3, 123) <= input(13);
output(3, 124) <= input(14);
output(3, 125) <= input(15);
output(3, 126) <= input(34);
output(3, 127) <= input(35);
output(3, 128) <= input(2);
output(3, 129) <= input(3);
output(3, 130) <= input(4);
output(3, 131) <= input(5);
output(3, 132) <= input(6);
output(3, 133) <= input(7);
output(3, 134) <= input(8);
output(3, 135) <= input(9);
output(3, 136) <= input(10);
output(3, 137) <= input(11);
output(3, 138) <= input(12);
output(3, 139) <= input(13);
output(3, 140) <= input(14);
output(3, 141) <= input(15);
output(3, 142) <= input(34);
output(3, 143) <= input(35);
output(3, 144) <= input(2);
output(3, 145) <= input(3);
output(3, 146) <= input(4);
output(3, 147) <= input(5);
output(3, 148) <= input(6);
output(3, 149) <= input(7);
output(3, 150) <= input(8);
output(3, 151) <= input(9);
output(3, 152) <= input(10);
output(3, 153) <= input(11);
output(3, 154) <= input(12);
output(3, 155) <= input(13);
output(3, 156) <= input(14);
output(3, 157) <= input(15);
output(3, 158) <= input(34);
output(3, 159) <= input(35);
output(3, 160) <= input(2);
output(3, 161) <= input(3);
output(3, 162) <= input(4);
output(3, 163) <= input(5);
output(3, 164) <= input(6);
output(3, 165) <= input(7);
output(3, 166) <= input(8);
output(3, 167) <= input(9);
output(3, 168) <= input(10);
output(3, 169) <= input(11);
output(3, 170) <= input(12);
output(3, 171) <= input(13);
output(3, 172) <= input(14);
output(3, 173) <= input(15);
output(3, 174) <= input(34);
output(3, 175) <= input(35);
output(3, 176) <= input(2);
output(3, 177) <= input(3);
output(3, 178) <= input(4);
output(3, 179) <= input(5);
output(3, 180) <= input(6);
output(3, 181) <= input(7);
output(3, 182) <= input(8);
output(3, 183) <= input(9);
output(3, 184) <= input(10);
output(3, 185) <= input(11);
output(3, 186) <= input(12);
output(3, 187) <= input(13);
output(3, 188) <= input(14);
output(3, 189) <= input(15);
output(3, 190) <= input(34);
output(3, 191) <= input(35);
output(3, 192) <= input(2);
output(3, 193) <= input(3);
output(3, 194) <= input(4);
output(3, 195) <= input(5);
output(3, 196) <= input(6);
output(3, 197) <= input(7);
output(3, 198) <= input(8);
output(3, 199) <= input(9);
output(3, 200) <= input(10);
output(3, 201) <= input(11);
output(3, 202) <= input(12);
output(3, 203) <= input(13);
output(3, 204) <= input(14);
output(3, 205) <= input(15);
output(3, 206) <= input(34);
output(3, 207) <= input(35);
output(3, 208) <= input(2);
output(3, 209) <= input(3);
output(3, 210) <= input(4);
output(3, 211) <= input(5);
output(3, 212) <= input(6);
output(3, 213) <= input(7);
output(3, 214) <= input(8);
output(3, 215) <= input(9);
output(3, 216) <= input(10);
output(3, 217) <= input(11);
output(3, 218) <= input(12);
output(3, 219) <= input(13);
output(3, 220) <= input(14);
output(3, 221) <= input(15);
output(3, 222) <= input(34);
output(3, 223) <= input(35);
output(3, 224) <= input(2);
output(3, 225) <= input(3);
output(3, 226) <= input(4);
output(3, 227) <= input(5);
output(3, 228) <= input(6);
output(3, 229) <= input(7);
output(3, 230) <= input(8);
output(3, 231) <= input(9);
output(3, 232) <= input(10);
output(3, 233) <= input(11);
output(3, 234) <= input(12);
output(3, 235) <= input(13);
output(3, 236) <= input(14);
output(3, 237) <= input(15);
output(3, 238) <= input(34);
output(3, 239) <= input(35);
output(3, 240) <= input(2);
output(3, 241) <= input(3);
output(3, 242) <= input(4);
output(3, 243) <= input(5);
output(3, 244) <= input(6);
output(3, 245) <= input(7);
output(3, 246) <= input(8);
output(3, 247) <= input(9);
output(3, 248) <= input(10);
output(3, 249) <= input(11);
output(3, 250) <= input(12);
output(3, 251) <= input(13);
output(3, 252) <= input(14);
output(3, 253) <= input(15);
output(3, 254) <= input(34);
output(3, 255) <= input(35);
output(4, 0) <= input(19);
output(4, 1) <= input(20);
output(4, 2) <= input(21);
output(4, 3) <= input(22);
output(4, 4) <= input(23);
output(4, 5) <= input(24);
output(4, 6) <= input(25);
output(4, 7) <= input(26);
output(4, 8) <= input(27);
output(4, 9) <= input(28);
output(4, 10) <= input(29);
output(4, 11) <= input(30);
output(4, 12) <= input(31);
output(4, 13) <= input(33);
output(4, 14) <= input(36);
output(4, 15) <= input(37);
output(4, 16) <= input(19);
output(4, 17) <= input(20);
output(4, 18) <= input(21);
output(4, 19) <= input(22);
output(4, 20) <= input(23);
output(4, 21) <= input(24);
output(4, 22) <= input(25);
output(4, 23) <= input(26);
output(4, 24) <= input(27);
output(4, 25) <= input(28);
output(4, 26) <= input(29);
output(4, 27) <= input(30);
output(4, 28) <= input(31);
output(4, 29) <= input(33);
output(4, 30) <= input(36);
output(4, 31) <= input(37);
output(4, 32) <= input(19);
output(4, 33) <= input(20);
output(4, 34) <= input(21);
output(4, 35) <= input(22);
output(4, 36) <= input(23);
output(4, 37) <= input(24);
output(4, 38) <= input(25);
output(4, 39) <= input(26);
output(4, 40) <= input(27);
output(4, 41) <= input(28);
output(4, 42) <= input(29);
output(4, 43) <= input(30);
output(4, 44) <= input(31);
output(4, 45) <= input(33);
output(4, 46) <= input(36);
output(4, 47) <= input(37);
output(4, 48) <= input(19);
output(4, 49) <= input(20);
output(4, 50) <= input(21);
output(4, 51) <= input(22);
output(4, 52) <= input(23);
output(4, 53) <= input(24);
output(4, 54) <= input(25);
output(4, 55) <= input(26);
output(4, 56) <= input(27);
output(4, 57) <= input(28);
output(4, 58) <= input(29);
output(4, 59) <= input(30);
output(4, 60) <= input(31);
output(4, 61) <= input(33);
output(4, 62) <= input(36);
output(4, 63) <= input(37);
output(4, 64) <= input(19);
output(4, 65) <= input(20);
output(4, 66) <= input(21);
output(4, 67) <= input(22);
output(4, 68) <= input(23);
output(4, 69) <= input(24);
output(4, 70) <= input(25);
output(4, 71) <= input(26);
output(4, 72) <= input(27);
output(4, 73) <= input(28);
output(4, 74) <= input(29);
output(4, 75) <= input(30);
output(4, 76) <= input(31);
output(4, 77) <= input(33);
output(4, 78) <= input(36);
output(4, 79) <= input(37);
output(4, 80) <= input(19);
output(4, 81) <= input(20);
output(4, 82) <= input(21);
output(4, 83) <= input(22);
output(4, 84) <= input(23);
output(4, 85) <= input(24);
output(4, 86) <= input(25);
output(4, 87) <= input(26);
output(4, 88) <= input(27);
output(4, 89) <= input(28);
output(4, 90) <= input(29);
output(4, 91) <= input(30);
output(4, 92) <= input(31);
output(4, 93) <= input(33);
output(4, 94) <= input(36);
output(4, 95) <= input(37);
output(4, 96) <= input(19);
output(4, 97) <= input(20);
output(4, 98) <= input(21);
output(4, 99) <= input(22);
output(4, 100) <= input(23);
output(4, 101) <= input(24);
output(4, 102) <= input(25);
output(4, 103) <= input(26);
output(4, 104) <= input(27);
output(4, 105) <= input(28);
output(4, 106) <= input(29);
output(4, 107) <= input(30);
output(4, 108) <= input(31);
output(4, 109) <= input(33);
output(4, 110) <= input(36);
output(4, 111) <= input(37);
output(4, 112) <= input(19);
output(4, 113) <= input(20);
output(4, 114) <= input(21);
output(4, 115) <= input(22);
output(4, 116) <= input(23);
output(4, 117) <= input(24);
output(4, 118) <= input(25);
output(4, 119) <= input(26);
output(4, 120) <= input(27);
output(4, 121) <= input(28);
output(4, 122) <= input(29);
output(4, 123) <= input(30);
output(4, 124) <= input(31);
output(4, 125) <= input(33);
output(4, 126) <= input(36);
output(4, 127) <= input(37);
output(4, 128) <= input(19);
output(4, 129) <= input(20);
output(4, 130) <= input(21);
output(4, 131) <= input(22);
output(4, 132) <= input(23);
output(4, 133) <= input(24);
output(4, 134) <= input(25);
output(4, 135) <= input(26);
output(4, 136) <= input(27);
output(4, 137) <= input(28);
output(4, 138) <= input(29);
output(4, 139) <= input(30);
output(4, 140) <= input(31);
output(4, 141) <= input(33);
output(4, 142) <= input(36);
output(4, 143) <= input(37);
output(4, 144) <= input(19);
output(4, 145) <= input(20);
output(4, 146) <= input(21);
output(4, 147) <= input(22);
output(4, 148) <= input(23);
output(4, 149) <= input(24);
output(4, 150) <= input(25);
output(4, 151) <= input(26);
output(4, 152) <= input(27);
output(4, 153) <= input(28);
output(4, 154) <= input(29);
output(4, 155) <= input(30);
output(4, 156) <= input(31);
output(4, 157) <= input(33);
output(4, 158) <= input(36);
output(4, 159) <= input(37);
output(4, 160) <= input(19);
output(4, 161) <= input(20);
output(4, 162) <= input(21);
output(4, 163) <= input(22);
output(4, 164) <= input(23);
output(4, 165) <= input(24);
output(4, 166) <= input(25);
output(4, 167) <= input(26);
output(4, 168) <= input(27);
output(4, 169) <= input(28);
output(4, 170) <= input(29);
output(4, 171) <= input(30);
output(4, 172) <= input(31);
output(4, 173) <= input(33);
output(4, 174) <= input(36);
output(4, 175) <= input(37);
output(4, 176) <= input(19);
output(4, 177) <= input(20);
output(4, 178) <= input(21);
output(4, 179) <= input(22);
output(4, 180) <= input(23);
output(4, 181) <= input(24);
output(4, 182) <= input(25);
output(4, 183) <= input(26);
output(4, 184) <= input(27);
output(4, 185) <= input(28);
output(4, 186) <= input(29);
output(4, 187) <= input(30);
output(4, 188) <= input(31);
output(4, 189) <= input(33);
output(4, 190) <= input(36);
output(4, 191) <= input(37);
output(4, 192) <= input(19);
output(4, 193) <= input(20);
output(4, 194) <= input(21);
output(4, 195) <= input(22);
output(4, 196) <= input(23);
output(4, 197) <= input(24);
output(4, 198) <= input(25);
output(4, 199) <= input(26);
output(4, 200) <= input(27);
output(4, 201) <= input(28);
output(4, 202) <= input(29);
output(4, 203) <= input(30);
output(4, 204) <= input(31);
output(4, 205) <= input(33);
output(4, 206) <= input(36);
output(4, 207) <= input(37);
output(4, 208) <= input(19);
output(4, 209) <= input(20);
output(4, 210) <= input(21);
output(4, 211) <= input(22);
output(4, 212) <= input(23);
output(4, 213) <= input(24);
output(4, 214) <= input(25);
output(4, 215) <= input(26);
output(4, 216) <= input(27);
output(4, 217) <= input(28);
output(4, 218) <= input(29);
output(4, 219) <= input(30);
output(4, 220) <= input(31);
output(4, 221) <= input(33);
output(4, 222) <= input(36);
output(4, 223) <= input(37);
output(4, 224) <= input(19);
output(4, 225) <= input(20);
output(4, 226) <= input(21);
output(4, 227) <= input(22);
output(4, 228) <= input(23);
output(4, 229) <= input(24);
output(4, 230) <= input(25);
output(4, 231) <= input(26);
output(4, 232) <= input(27);
output(4, 233) <= input(28);
output(4, 234) <= input(29);
output(4, 235) <= input(30);
output(4, 236) <= input(31);
output(4, 237) <= input(33);
output(4, 238) <= input(36);
output(4, 239) <= input(37);
output(4, 240) <= input(3);
output(4, 241) <= input(4);
output(4, 242) <= input(5);
output(4, 243) <= input(6);
output(4, 244) <= input(7);
output(4, 245) <= input(8);
output(4, 246) <= input(9);
output(4, 247) <= input(10);
output(4, 248) <= input(11);
output(4, 249) <= input(12);
output(4, 250) <= input(13);
output(4, 251) <= input(14);
output(4, 252) <= input(15);
output(4, 253) <= input(34);
output(4, 254) <= input(35);
output(4, 255) <= input(38);
output(5, 0) <= input(3);
output(5, 1) <= input(4);
output(5, 2) <= input(5);
output(5, 3) <= input(6);
output(5, 4) <= input(7);
output(5, 5) <= input(8);
output(5, 6) <= input(9);
output(5, 7) <= input(10);
output(5, 8) <= input(11);
output(5, 9) <= input(12);
output(5, 10) <= input(13);
output(5, 11) <= input(14);
output(5, 12) <= input(15);
output(5, 13) <= input(34);
output(5, 14) <= input(35);
output(5, 15) <= input(38);
output(5, 16) <= input(3);
output(5, 17) <= input(4);
output(5, 18) <= input(5);
output(5, 19) <= input(6);
output(5, 20) <= input(7);
output(5, 21) <= input(8);
output(5, 22) <= input(9);
output(5, 23) <= input(10);
output(5, 24) <= input(11);
output(5, 25) <= input(12);
output(5, 26) <= input(13);
output(5, 27) <= input(14);
output(5, 28) <= input(15);
output(5, 29) <= input(34);
output(5, 30) <= input(35);
output(5, 31) <= input(38);
output(5, 32) <= input(3);
output(5, 33) <= input(4);
output(5, 34) <= input(5);
output(5, 35) <= input(6);
output(5, 36) <= input(7);
output(5, 37) <= input(8);
output(5, 38) <= input(9);
output(5, 39) <= input(10);
output(5, 40) <= input(11);
output(5, 41) <= input(12);
output(5, 42) <= input(13);
output(5, 43) <= input(14);
output(5, 44) <= input(15);
output(5, 45) <= input(34);
output(5, 46) <= input(35);
output(5, 47) <= input(38);
output(5, 48) <= input(3);
output(5, 49) <= input(4);
output(5, 50) <= input(5);
output(5, 51) <= input(6);
output(5, 52) <= input(7);
output(5, 53) <= input(8);
output(5, 54) <= input(9);
output(5, 55) <= input(10);
output(5, 56) <= input(11);
output(5, 57) <= input(12);
output(5, 58) <= input(13);
output(5, 59) <= input(14);
output(5, 60) <= input(15);
output(5, 61) <= input(34);
output(5, 62) <= input(35);
output(5, 63) <= input(38);
output(5, 64) <= input(3);
output(5, 65) <= input(4);
output(5, 66) <= input(5);
output(5, 67) <= input(6);
output(5, 68) <= input(7);
output(5, 69) <= input(8);
output(5, 70) <= input(9);
output(5, 71) <= input(10);
output(5, 72) <= input(11);
output(5, 73) <= input(12);
output(5, 74) <= input(13);
output(5, 75) <= input(14);
output(5, 76) <= input(15);
output(5, 77) <= input(34);
output(5, 78) <= input(35);
output(5, 79) <= input(38);
output(5, 80) <= input(3);
output(5, 81) <= input(4);
output(5, 82) <= input(5);
output(5, 83) <= input(6);
output(5, 84) <= input(7);
output(5, 85) <= input(8);
output(5, 86) <= input(9);
output(5, 87) <= input(10);
output(5, 88) <= input(11);
output(5, 89) <= input(12);
output(5, 90) <= input(13);
output(5, 91) <= input(14);
output(5, 92) <= input(15);
output(5, 93) <= input(34);
output(5, 94) <= input(35);
output(5, 95) <= input(38);
output(5, 96) <= input(3);
output(5, 97) <= input(4);
output(5, 98) <= input(5);
output(5, 99) <= input(6);
output(5, 100) <= input(7);
output(5, 101) <= input(8);
output(5, 102) <= input(9);
output(5, 103) <= input(10);
output(5, 104) <= input(11);
output(5, 105) <= input(12);
output(5, 106) <= input(13);
output(5, 107) <= input(14);
output(5, 108) <= input(15);
output(5, 109) <= input(34);
output(5, 110) <= input(35);
output(5, 111) <= input(38);
output(5, 112) <= input(20);
output(5, 113) <= input(21);
output(5, 114) <= input(22);
output(5, 115) <= input(23);
output(5, 116) <= input(24);
output(5, 117) <= input(25);
output(5, 118) <= input(26);
output(5, 119) <= input(27);
output(5, 120) <= input(28);
output(5, 121) <= input(29);
output(5, 122) <= input(30);
output(5, 123) <= input(31);
output(5, 124) <= input(33);
output(5, 125) <= input(36);
output(5, 126) <= input(37);
output(5, 127) <= input(39);
output(5, 128) <= input(20);
output(5, 129) <= input(21);
output(5, 130) <= input(22);
output(5, 131) <= input(23);
output(5, 132) <= input(24);
output(5, 133) <= input(25);
output(5, 134) <= input(26);
output(5, 135) <= input(27);
output(5, 136) <= input(28);
output(5, 137) <= input(29);
output(5, 138) <= input(30);
output(5, 139) <= input(31);
output(5, 140) <= input(33);
output(5, 141) <= input(36);
output(5, 142) <= input(37);
output(5, 143) <= input(39);
output(5, 144) <= input(20);
output(5, 145) <= input(21);
output(5, 146) <= input(22);
output(5, 147) <= input(23);
output(5, 148) <= input(24);
output(5, 149) <= input(25);
output(5, 150) <= input(26);
output(5, 151) <= input(27);
output(5, 152) <= input(28);
output(5, 153) <= input(29);
output(5, 154) <= input(30);
output(5, 155) <= input(31);
output(5, 156) <= input(33);
output(5, 157) <= input(36);
output(5, 158) <= input(37);
output(5, 159) <= input(39);
output(5, 160) <= input(20);
output(5, 161) <= input(21);
output(5, 162) <= input(22);
output(5, 163) <= input(23);
output(5, 164) <= input(24);
output(5, 165) <= input(25);
output(5, 166) <= input(26);
output(5, 167) <= input(27);
output(5, 168) <= input(28);
output(5, 169) <= input(29);
output(5, 170) <= input(30);
output(5, 171) <= input(31);
output(5, 172) <= input(33);
output(5, 173) <= input(36);
output(5, 174) <= input(37);
output(5, 175) <= input(39);
output(5, 176) <= input(20);
output(5, 177) <= input(21);
output(5, 178) <= input(22);
output(5, 179) <= input(23);
output(5, 180) <= input(24);
output(5, 181) <= input(25);
output(5, 182) <= input(26);
output(5, 183) <= input(27);
output(5, 184) <= input(28);
output(5, 185) <= input(29);
output(5, 186) <= input(30);
output(5, 187) <= input(31);
output(5, 188) <= input(33);
output(5, 189) <= input(36);
output(5, 190) <= input(37);
output(5, 191) <= input(39);
output(5, 192) <= input(20);
output(5, 193) <= input(21);
output(5, 194) <= input(22);
output(5, 195) <= input(23);
output(5, 196) <= input(24);
output(5, 197) <= input(25);
output(5, 198) <= input(26);
output(5, 199) <= input(27);
output(5, 200) <= input(28);
output(5, 201) <= input(29);
output(5, 202) <= input(30);
output(5, 203) <= input(31);
output(5, 204) <= input(33);
output(5, 205) <= input(36);
output(5, 206) <= input(37);
output(5, 207) <= input(39);
output(5, 208) <= input(20);
output(5, 209) <= input(21);
output(5, 210) <= input(22);
output(5, 211) <= input(23);
output(5, 212) <= input(24);
output(5, 213) <= input(25);
output(5, 214) <= input(26);
output(5, 215) <= input(27);
output(5, 216) <= input(28);
output(5, 217) <= input(29);
output(5, 218) <= input(30);
output(5, 219) <= input(31);
output(5, 220) <= input(33);
output(5, 221) <= input(36);
output(5, 222) <= input(37);
output(5, 223) <= input(39);
output(5, 224) <= input(20);
output(5, 225) <= input(21);
output(5, 226) <= input(22);
output(5, 227) <= input(23);
output(5, 228) <= input(24);
output(5, 229) <= input(25);
output(5, 230) <= input(26);
output(5, 231) <= input(27);
output(5, 232) <= input(28);
output(5, 233) <= input(29);
output(5, 234) <= input(30);
output(5, 235) <= input(31);
output(5, 236) <= input(33);
output(5, 237) <= input(36);
output(5, 238) <= input(37);
output(5, 239) <= input(39);
output(5, 240) <= input(4);
output(5, 241) <= input(5);
output(5, 242) <= input(6);
output(5, 243) <= input(7);
output(5, 244) <= input(8);
output(5, 245) <= input(9);
output(5, 246) <= input(10);
output(5, 247) <= input(11);
output(5, 248) <= input(12);
output(5, 249) <= input(13);
output(5, 250) <= input(14);
output(5, 251) <= input(15);
output(5, 252) <= input(34);
output(5, 253) <= input(35);
output(5, 254) <= input(38);
output(5, 255) <= input(40);
output(6, 0) <= input(20);
output(6, 1) <= input(21);
output(6, 2) <= input(22);
output(6, 3) <= input(23);
output(6, 4) <= input(24);
output(6, 5) <= input(25);
output(6, 6) <= input(26);
output(6, 7) <= input(27);
output(6, 8) <= input(28);
output(6, 9) <= input(29);
output(6, 10) <= input(30);
output(6, 11) <= input(31);
output(6, 12) <= input(33);
output(6, 13) <= input(36);
output(6, 14) <= input(37);
output(6, 15) <= input(39);
output(6, 16) <= input(20);
output(6, 17) <= input(21);
output(6, 18) <= input(22);
output(6, 19) <= input(23);
output(6, 20) <= input(24);
output(6, 21) <= input(25);
output(6, 22) <= input(26);
output(6, 23) <= input(27);
output(6, 24) <= input(28);
output(6, 25) <= input(29);
output(6, 26) <= input(30);
output(6, 27) <= input(31);
output(6, 28) <= input(33);
output(6, 29) <= input(36);
output(6, 30) <= input(37);
output(6, 31) <= input(39);
output(6, 32) <= input(20);
output(6, 33) <= input(21);
output(6, 34) <= input(22);
output(6, 35) <= input(23);
output(6, 36) <= input(24);
output(6, 37) <= input(25);
output(6, 38) <= input(26);
output(6, 39) <= input(27);
output(6, 40) <= input(28);
output(6, 41) <= input(29);
output(6, 42) <= input(30);
output(6, 43) <= input(31);
output(6, 44) <= input(33);
output(6, 45) <= input(36);
output(6, 46) <= input(37);
output(6, 47) <= input(39);
output(6, 48) <= input(20);
output(6, 49) <= input(21);
output(6, 50) <= input(22);
output(6, 51) <= input(23);
output(6, 52) <= input(24);
output(6, 53) <= input(25);
output(6, 54) <= input(26);
output(6, 55) <= input(27);
output(6, 56) <= input(28);
output(6, 57) <= input(29);
output(6, 58) <= input(30);
output(6, 59) <= input(31);
output(6, 60) <= input(33);
output(6, 61) <= input(36);
output(6, 62) <= input(37);
output(6, 63) <= input(39);
output(6, 64) <= input(20);
output(6, 65) <= input(21);
output(6, 66) <= input(22);
output(6, 67) <= input(23);
output(6, 68) <= input(24);
output(6, 69) <= input(25);
output(6, 70) <= input(26);
output(6, 71) <= input(27);
output(6, 72) <= input(28);
output(6, 73) <= input(29);
output(6, 74) <= input(30);
output(6, 75) <= input(31);
output(6, 76) <= input(33);
output(6, 77) <= input(36);
output(6, 78) <= input(37);
output(6, 79) <= input(39);
output(6, 80) <= input(4);
output(6, 81) <= input(5);
output(6, 82) <= input(6);
output(6, 83) <= input(7);
output(6, 84) <= input(8);
output(6, 85) <= input(9);
output(6, 86) <= input(10);
output(6, 87) <= input(11);
output(6, 88) <= input(12);
output(6, 89) <= input(13);
output(6, 90) <= input(14);
output(6, 91) <= input(15);
output(6, 92) <= input(34);
output(6, 93) <= input(35);
output(6, 94) <= input(38);
output(6, 95) <= input(40);
output(6, 96) <= input(4);
output(6, 97) <= input(5);
output(6, 98) <= input(6);
output(6, 99) <= input(7);
output(6, 100) <= input(8);
output(6, 101) <= input(9);
output(6, 102) <= input(10);
output(6, 103) <= input(11);
output(6, 104) <= input(12);
output(6, 105) <= input(13);
output(6, 106) <= input(14);
output(6, 107) <= input(15);
output(6, 108) <= input(34);
output(6, 109) <= input(35);
output(6, 110) <= input(38);
output(6, 111) <= input(40);
output(6, 112) <= input(4);
output(6, 113) <= input(5);
output(6, 114) <= input(6);
output(6, 115) <= input(7);
output(6, 116) <= input(8);
output(6, 117) <= input(9);
output(6, 118) <= input(10);
output(6, 119) <= input(11);
output(6, 120) <= input(12);
output(6, 121) <= input(13);
output(6, 122) <= input(14);
output(6, 123) <= input(15);
output(6, 124) <= input(34);
output(6, 125) <= input(35);
output(6, 126) <= input(38);
output(6, 127) <= input(40);
output(6, 128) <= input(4);
output(6, 129) <= input(5);
output(6, 130) <= input(6);
output(6, 131) <= input(7);
output(6, 132) <= input(8);
output(6, 133) <= input(9);
output(6, 134) <= input(10);
output(6, 135) <= input(11);
output(6, 136) <= input(12);
output(6, 137) <= input(13);
output(6, 138) <= input(14);
output(6, 139) <= input(15);
output(6, 140) <= input(34);
output(6, 141) <= input(35);
output(6, 142) <= input(38);
output(6, 143) <= input(40);
output(6, 144) <= input(4);
output(6, 145) <= input(5);
output(6, 146) <= input(6);
output(6, 147) <= input(7);
output(6, 148) <= input(8);
output(6, 149) <= input(9);
output(6, 150) <= input(10);
output(6, 151) <= input(11);
output(6, 152) <= input(12);
output(6, 153) <= input(13);
output(6, 154) <= input(14);
output(6, 155) <= input(15);
output(6, 156) <= input(34);
output(6, 157) <= input(35);
output(6, 158) <= input(38);
output(6, 159) <= input(40);
output(6, 160) <= input(21);
output(6, 161) <= input(22);
output(6, 162) <= input(23);
output(6, 163) <= input(24);
output(6, 164) <= input(25);
output(6, 165) <= input(26);
output(6, 166) <= input(27);
output(6, 167) <= input(28);
output(6, 168) <= input(29);
output(6, 169) <= input(30);
output(6, 170) <= input(31);
output(6, 171) <= input(33);
output(6, 172) <= input(36);
output(6, 173) <= input(37);
output(6, 174) <= input(39);
output(6, 175) <= input(41);
output(6, 176) <= input(21);
output(6, 177) <= input(22);
output(6, 178) <= input(23);
output(6, 179) <= input(24);
output(6, 180) <= input(25);
output(6, 181) <= input(26);
output(6, 182) <= input(27);
output(6, 183) <= input(28);
output(6, 184) <= input(29);
output(6, 185) <= input(30);
output(6, 186) <= input(31);
output(6, 187) <= input(33);
output(6, 188) <= input(36);
output(6, 189) <= input(37);
output(6, 190) <= input(39);
output(6, 191) <= input(41);
output(6, 192) <= input(21);
output(6, 193) <= input(22);
output(6, 194) <= input(23);
output(6, 195) <= input(24);
output(6, 196) <= input(25);
output(6, 197) <= input(26);
output(6, 198) <= input(27);
output(6, 199) <= input(28);
output(6, 200) <= input(29);
output(6, 201) <= input(30);
output(6, 202) <= input(31);
output(6, 203) <= input(33);
output(6, 204) <= input(36);
output(6, 205) <= input(37);
output(6, 206) <= input(39);
output(6, 207) <= input(41);
output(6, 208) <= input(21);
output(6, 209) <= input(22);
output(6, 210) <= input(23);
output(6, 211) <= input(24);
output(6, 212) <= input(25);
output(6, 213) <= input(26);
output(6, 214) <= input(27);
output(6, 215) <= input(28);
output(6, 216) <= input(29);
output(6, 217) <= input(30);
output(6, 218) <= input(31);
output(6, 219) <= input(33);
output(6, 220) <= input(36);
output(6, 221) <= input(37);
output(6, 222) <= input(39);
output(6, 223) <= input(41);
output(6, 224) <= input(21);
output(6, 225) <= input(22);
output(6, 226) <= input(23);
output(6, 227) <= input(24);
output(6, 228) <= input(25);
output(6, 229) <= input(26);
output(6, 230) <= input(27);
output(6, 231) <= input(28);
output(6, 232) <= input(29);
output(6, 233) <= input(30);
output(6, 234) <= input(31);
output(6, 235) <= input(33);
output(6, 236) <= input(36);
output(6, 237) <= input(37);
output(6, 238) <= input(39);
output(6, 239) <= input(41);
output(6, 240) <= input(5);
output(6, 241) <= input(6);
output(6, 242) <= input(7);
output(6, 243) <= input(8);
output(6, 244) <= input(9);
output(6, 245) <= input(10);
output(6, 246) <= input(11);
output(6, 247) <= input(12);
output(6, 248) <= input(13);
output(6, 249) <= input(14);
output(6, 250) <= input(15);
output(6, 251) <= input(34);
output(6, 252) <= input(35);
output(6, 253) <= input(38);
output(6, 254) <= input(40);
output(6, 255) <= input(42);
output(7, 0) <= input(4);
output(7, 1) <= input(5);
output(7, 2) <= input(6);
output(7, 3) <= input(7);
output(7, 4) <= input(8);
output(7, 5) <= input(9);
output(7, 6) <= input(10);
output(7, 7) <= input(11);
output(7, 8) <= input(12);
output(7, 9) <= input(13);
output(7, 10) <= input(14);
output(7, 11) <= input(15);
output(7, 12) <= input(34);
output(7, 13) <= input(35);
output(7, 14) <= input(38);
output(7, 15) <= input(40);
output(7, 16) <= input(4);
output(7, 17) <= input(5);
output(7, 18) <= input(6);
output(7, 19) <= input(7);
output(7, 20) <= input(8);
output(7, 21) <= input(9);
output(7, 22) <= input(10);
output(7, 23) <= input(11);
output(7, 24) <= input(12);
output(7, 25) <= input(13);
output(7, 26) <= input(14);
output(7, 27) <= input(15);
output(7, 28) <= input(34);
output(7, 29) <= input(35);
output(7, 30) <= input(38);
output(7, 31) <= input(40);
output(7, 32) <= input(4);
output(7, 33) <= input(5);
output(7, 34) <= input(6);
output(7, 35) <= input(7);
output(7, 36) <= input(8);
output(7, 37) <= input(9);
output(7, 38) <= input(10);
output(7, 39) <= input(11);
output(7, 40) <= input(12);
output(7, 41) <= input(13);
output(7, 42) <= input(14);
output(7, 43) <= input(15);
output(7, 44) <= input(34);
output(7, 45) <= input(35);
output(7, 46) <= input(38);
output(7, 47) <= input(40);
output(7, 48) <= input(21);
output(7, 49) <= input(22);
output(7, 50) <= input(23);
output(7, 51) <= input(24);
output(7, 52) <= input(25);
output(7, 53) <= input(26);
output(7, 54) <= input(27);
output(7, 55) <= input(28);
output(7, 56) <= input(29);
output(7, 57) <= input(30);
output(7, 58) <= input(31);
output(7, 59) <= input(33);
output(7, 60) <= input(36);
output(7, 61) <= input(37);
output(7, 62) <= input(39);
output(7, 63) <= input(41);
output(7, 64) <= input(21);
output(7, 65) <= input(22);
output(7, 66) <= input(23);
output(7, 67) <= input(24);
output(7, 68) <= input(25);
output(7, 69) <= input(26);
output(7, 70) <= input(27);
output(7, 71) <= input(28);
output(7, 72) <= input(29);
output(7, 73) <= input(30);
output(7, 74) <= input(31);
output(7, 75) <= input(33);
output(7, 76) <= input(36);
output(7, 77) <= input(37);
output(7, 78) <= input(39);
output(7, 79) <= input(41);
output(7, 80) <= input(21);
output(7, 81) <= input(22);
output(7, 82) <= input(23);
output(7, 83) <= input(24);
output(7, 84) <= input(25);
output(7, 85) <= input(26);
output(7, 86) <= input(27);
output(7, 87) <= input(28);
output(7, 88) <= input(29);
output(7, 89) <= input(30);
output(7, 90) <= input(31);
output(7, 91) <= input(33);
output(7, 92) <= input(36);
output(7, 93) <= input(37);
output(7, 94) <= input(39);
output(7, 95) <= input(41);
output(7, 96) <= input(21);
output(7, 97) <= input(22);
output(7, 98) <= input(23);
output(7, 99) <= input(24);
output(7, 100) <= input(25);
output(7, 101) <= input(26);
output(7, 102) <= input(27);
output(7, 103) <= input(28);
output(7, 104) <= input(29);
output(7, 105) <= input(30);
output(7, 106) <= input(31);
output(7, 107) <= input(33);
output(7, 108) <= input(36);
output(7, 109) <= input(37);
output(7, 110) <= input(39);
output(7, 111) <= input(41);
output(7, 112) <= input(5);
output(7, 113) <= input(6);
output(7, 114) <= input(7);
output(7, 115) <= input(8);
output(7, 116) <= input(9);
output(7, 117) <= input(10);
output(7, 118) <= input(11);
output(7, 119) <= input(12);
output(7, 120) <= input(13);
output(7, 121) <= input(14);
output(7, 122) <= input(15);
output(7, 123) <= input(34);
output(7, 124) <= input(35);
output(7, 125) <= input(38);
output(7, 126) <= input(40);
output(7, 127) <= input(42);
output(7, 128) <= input(5);
output(7, 129) <= input(6);
output(7, 130) <= input(7);
output(7, 131) <= input(8);
output(7, 132) <= input(9);
output(7, 133) <= input(10);
output(7, 134) <= input(11);
output(7, 135) <= input(12);
output(7, 136) <= input(13);
output(7, 137) <= input(14);
output(7, 138) <= input(15);
output(7, 139) <= input(34);
output(7, 140) <= input(35);
output(7, 141) <= input(38);
output(7, 142) <= input(40);
output(7, 143) <= input(42);
output(7, 144) <= input(5);
output(7, 145) <= input(6);
output(7, 146) <= input(7);
output(7, 147) <= input(8);
output(7, 148) <= input(9);
output(7, 149) <= input(10);
output(7, 150) <= input(11);
output(7, 151) <= input(12);
output(7, 152) <= input(13);
output(7, 153) <= input(14);
output(7, 154) <= input(15);
output(7, 155) <= input(34);
output(7, 156) <= input(35);
output(7, 157) <= input(38);
output(7, 158) <= input(40);
output(7, 159) <= input(42);
output(7, 160) <= input(5);
output(7, 161) <= input(6);
output(7, 162) <= input(7);
output(7, 163) <= input(8);
output(7, 164) <= input(9);
output(7, 165) <= input(10);
output(7, 166) <= input(11);
output(7, 167) <= input(12);
output(7, 168) <= input(13);
output(7, 169) <= input(14);
output(7, 170) <= input(15);
output(7, 171) <= input(34);
output(7, 172) <= input(35);
output(7, 173) <= input(38);
output(7, 174) <= input(40);
output(7, 175) <= input(42);
output(7, 176) <= input(22);
output(7, 177) <= input(23);
output(7, 178) <= input(24);
output(7, 179) <= input(25);
output(7, 180) <= input(26);
output(7, 181) <= input(27);
output(7, 182) <= input(28);
output(7, 183) <= input(29);
output(7, 184) <= input(30);
output(7, 185) <= input(31);
output(7, 186) <= input(33);
output(7, 187) <= input(36);
output(7, 188) <= input(37);
output(7, 189) <= input(39);
output(7, 190) <= input(41);
output(7, 191) <= input(43);
output(7, 192) <= input(22);
output(7, 193) <= input(23);
output(7, 194) <= input(24);
output(7, 195) <= input(25);
output(7, 196) <= input(26);
output(7, 197) <= input(27);
output(7, 198) <= input(28);
output(7, 199) <= input(29);
output(7, 200) <= input(30);
output(7, 201) <= input(31);
output(7, 202) <= input(33);
output(7, 203) <= input(36);
output(7, 204) <= input(37);
output(7, 205) <= input(39);
output(7, 206) <= input(41);
output(7, 207) <= input(43);
output(7, 208) <= input(22);
output(7, 209) <= input(23);
output(7, 210) <= input(24);
output(7, 211) <= input(25);
output(7, 212) <= input(26);
output(7, 213) <= input(27);
output(7, 214) <= input(28);
output(7, 215) <= input(29);
output(7, 216) <= input(30);
output(7, 217) <= input(31);
output(7, 218) <= input(33);
output(7, 219) <= input(36);
output(7, 220) <= input(37);
output(7, 221) <= input(39);
output(7, 222) <= input(41);
output(7, 223) <= input(43);
output(7, 224) <= input(22);
output(7, 225) <= input(23);
output(7, 226) <= input(24);
output(7, 227) <= input(25);
output(7, 228) <= input(26);
output(7, 229) <= input(27);
output(7, 230) <= input(28);
output(7, 231) <= input(29);
output(7, 232) <= input(30);
output(7, 233) <= input(31);
output(7, 234) <= input(33);
output(7, 235) <= input(36);
output(7, 236) <= input(37);
output(7, 237) <= input(39);
output(7, 238) <= input(41);
output(7, 239) <= input(43);
output(7, 240) <= input(6);
output(7, 241) <= input(7);
output(7, 242) <= input(8);
output(7, 243) <= input(9);
output(7, 244) <= input(10);
output(7, 245) <= input(11);
output(7, 246) <= input(12);
output(7, 247) <= input(13);
output(7, 248) <= input(14);
output(7, 249) <= input(15);
output(7, 250) <= input(34);
output(7, 251) <= input(35);
output(7, 252) <= input(38);
output(7, 253) <= input(40);
output(7, 254) <= input(42);
output(7, 255) <= input(44);
when "1110" =>
output(0, 0) <= input(0);
output(0, 1) <= input(1);
output(0, 2) <= input(2);
output(0, 3) <= input(3);
output(0, 4) <= input(4);
output(0, 5) <= input(5);
output(0, 6) <= input(6);
output(0, 7) <= input(7);
output(0, 8) <= input(8);
output(0, 9) <= input(9);
output(0, 10) <= input(10);
output(0, 11) <= input(11);
output(0, 12) <= input(12);
output(0, 13) <= input(13);
output(0, 14) <= input(14);
output(0, 15) <= input(15);
output(0, 16) <= input(0);
output(0, 17) <= input(1);
output(0, 18) <= input(2);
output(0, 19) <= input(3);
output(0, 20) <= input(4);
output(0, 21) <= input(5);
output(0, 22) <= input(6);
output(0, 23) <= input(7);
output(0, 24) <= input(8);
output(0, 25) <= input(9);
output(0, 26) <= input(10);
output(0, 27) <= input(11);
output(0, 28) <= input(12);
output(0, 29) <= input(13);
output(0, 30) <= input(14);
output(0, 31) <= input(15);
output(0, 32) <= input(16);
output(0, 33) <= input(17);
output(0, 34) <= input(18);
output(0, 35) <= input(19);
output(0, 36) <= input(20);
output(0, 37) <= input(21);
output(0, 38) <= input(22);
output(0, 39) <= input(23);
output(0, 40) <= input(24);
output(0, 41) <= input(25);
output(0, 42) <= input(26);
output(0, 43) <= input(27);
output(0, 44) <= input(28);
output(0, 45) <= input(29);
output(0, 46) <= input(30);
output(0, 47) <= input(31);
output(0, 48) <= input(16);
output(0, 49) <= input(17);
output(0, 50) <= input(18);
output(0, 51) <= input(19);
output(0, 52) <= input(20);
output(0, 53) <= input(21);
output(0, 54) <= input(22);
output(0, 55) <= input(23);
output(0, 56) <= input(24);
output(0, 57) <= input(25);
output(0, 58) <= input(26);
output(0, 59) <= input(27);
output(0, 60) <= input(28);
output(0, 61) <= input(29);
output(0, 62) <= input(30);
output(0, 63) <= input(31);
output(0, 64) <= input(16);
output(0, 65) <= input(17);
output(0, 66) <= input(18);
output(0, 67) <= input(19);
output(0, 68) <= input(20);
output(0, 69) <= input(21);
output(0, 70) <= input(22);
output(0, 71) <= input(23);
output(0, 72) <= input(24);
output(0, 73) <= input(25);
output(0, 74) <= input(26);
output(0, 75) <= input(27);
output(0, 76) <= input(28);
output(0, 77) <= input(29);
output(0, 78) <= input(30);
output(0, 79) <= input(31);
output(0, 80) <= input(1);
output(0, 81) <= input(2);
output(0, 82) <= input(3);
output(0, 83) <= input(4);
output(0, 84) <= input(5);
output(0, 85) <= input(6);
output(0, 86) <= input(7);
output(0, 87) <= input(8);
output(0, 88) <= input(9);
output(0, 89) <= input(10);
output(0, 90) <= input(11);
output(0, 91) <= input(12);
output(0, 92) <= input(13);
output(0, 93) <= input(14);
output(0, 94) <= input(15);
output(0, 95) <= input(32);
output(0, 96) <= input(1);
output(0, 97) <= input(2);
output(0, 98) <= input(3);
output(0, 99) <= input(4);
output(0, 100) <= input(5);
output(0, 101) <= input(6);
output(0, 102) <= input(7);
output(0, 103) <= input(8);
output(0, 104) <= input(9);
output(0, 105) <= input(10);
output(0, 106) <= input(11);
output(0, 107) <= input(12);
output(0, 108) <= input(13);
output(0, 109) <= input(14);
output(0, 110) <= input(15);
output(0, 111) <= input(32);
output(0, 112) <= input(17);
output(0, 113) <= input(18);
output(0, 114) <= input(19);
output(0, 115) <= input(20);
output(0, 116) <= input(21);
output(0, 117) <= input(22);
output(0, 118) <= input(23);
output(0, 119) <= input(24);
output(0, 120) <= input(25);
output(0, 121) <= input(26);
output(0, 122) <= input(27);
output(0, 123) <= input(28);
output(0, 124) <= input(29);
output(0, 125) <= input(30);
output(0, 126) <= input(31);
output(0, 127) <= input(33);
output(0, 128) <= input(17);
output(0, 129) <= input(18);
output(0, 130) <= input(19);
output(0, 131) <= input(20);
output(0, 132) <= input(21);
output(0, 133) <= input(22);
output(0, 134) <= input(23);
output(0, 135) <= input(24);
output(0, 136) <= input(25);
output(0, 137) <= input(26);
output(0, 138) <= input(27);
output(0, 139) <= input(28);
output(0, 140) <= input(29);
output(0, 141) <= input(30);
output(0, 142) <= input(31);
output(0, 143) <= input(33);
output(0, 144) <= input(17);
output(0, 145) <= input(18);
output(0, 146) <= input(19);
output(0, 147) <= input(20);
output(0, 148) <= input(21);
output(0, 149) <= input(22);
output(0, 150) <= input(23);
output(0, 151) <= input(24);
output(0, 152) <= input(25);
output(0, 153) <= input(26);
output(0, 154) <= input(27);
output(0, 155) <= input(28);
output(0, 156) <= input(29);
output(0, 157) <= input(30);
output(0, 158) <= input(31);
output(0, 159) <= input(33);
output(0, 160) <= input(2);
output(0, 161) <= input(3);
output(0, 162) <= input(4);
output(0, 163) <= input(5);
output(0, 164) <= input(6);
output(0, 165) <= input(7);
output(0, 166) <= input(8);
output(0, 167) <= input(9);
output(0, 168) <= input(10);
output(0, 169) <= input(11);
output(0, 170) <= input(12);
output(0, 171) <= input(13);
output(0, 172) <= input(14);
output(0, 173) <= input(15);
output(0, 174) <= input(32);
output(0, 175) <= input(34);
output(0, 176) <= input(2);
output(0, 177) <= input(3);
output(0, 178) <= input(4);
output(0, 179) <= input(5);
output(0, 180) <= input(6);
output(0, 181) <= input(7);
output(0, 182) <= input(8);
output(0, 183) <= input(9);
output(0, 184) <= input(10);
output(0, 185) <= input(11);
output(0, 186) <= input(12);
output(0, 187) <= input(13);
output(0, 188) <= input(14);
output(0, 189) <= input(15);
output(0, 190) <= input(32);
output(0, 191) <= input(34);
output(0, 192) <= input(2);
output(0, 193) <= input(3);
output(0, 194) <= input(4);
output(0, 195) <= input(5);
output(0, 196) <= input(6);
output(0, 197) <= input(7);
output(0, 198) <= input(8);
output(0, 199) <= input(9);
output(0, 200) <= input(10);
output(0, 201) <= input(11);
output(0, 202) <= input(12);
output(0, 203) <= input(13);
output(0, 204) <= input(14);
output(0, 205) <= input(15);
output(0, 206) <= input(32);
output(0, 207) <= input(34);
output(0, 208) <= input(18);
output(0, 209) <= input(19);
output(0, 210) <= input(20);
output(0, 211) <= input(21);
output(0, 212) <= input(22);
output(0, 213) <= input(23);
output(0, 214) <= input(24);
output(0, 215) <= input(25);
output(0, 216) <= input(26);
output(0, 217) <= input(27);
output(0, 218) <= input(28);
output(0, 219) <= input(29);
output(0, 220) <= input(30);
output(0, 221) <= input(31);
output(0, 222) <= input(33);
output(0, 223) <= input(35);
output(0, 224) <= input(18);
output(0, 225) <= input(19);
output(0, 226) <= input(20);
output(0, 227) <= input(21);
output(0, 228) <= input(22);
output(0, 229) <= input(23);
output(0, 230) <= input(24);
output(0, 231) <= input(25);
output(0, 232) <= input(26);
output(0, 233) <= input(27);
output(0, 234) <= input(28);
output(0, 235) <= input(29);
output(0, 236) <= input(30);
output(0, 237) <= input(31);
output(0, 238) <= input(33);
output(0, 239) <= input(35);
output(0, 240) <= input(3);
output(0, 241) <= input(4);
output(0, 242) <= input(5);
output(0, 243) <= input(6);
output(0, 244) <= input(7);
output(0, 245) <= input(8);
output(0, 246) <= input(9);
output(0, 247) <= input(10);
output(0, 248) <= input(11);
output(0, 249) <= input(12);
output(0, 250) <= input(13);
output(0, 251) <= input(14);
output(0, 252) <= input(15);
output(0, 253) <= input(32);
output(0, 254) <= input(34);
output(0, 255) <= input(36);
output(1, 0) <= input(1);
output(1, 1) <= input(2);
output(1, 2) <= input(3);
output(1, 3) <= input(4);
output(1, 4) <= input(5);
output(1, 5) <= input(6);
output(1, 6) <= input(7);
output(1, 7) <= input(8);
output(1, 8) <= input(9);
output(1, 9) <= input(10);
output(1, 10) <= input(11);
output(1, 11) <= input(12);
output(1, 12) <= input(13);
output(1, 13) <= input(14);
output(1, 14) <= input(15);
output(1, 15) <= input(32);
output(1, 16) <= input(17);
output(1, 17) <= input(18);
output(1, 18) <= input(19);
output(1, 19) <= input(20);
output(1, 20) <= input(21);
output(1, 21) <= input(22);
output(1, 22) <= input(23);
output(1, 23) <= input(24);
output(1, 24) <= input(25);
output(1, 25) <= input(26);
output(1, 26) <= input(27);
output(1, 27) <= input(28);
output(1, 28) <= input(29);
output(1, 29) <= input(30);
output(1, 30) <= input(31);
output(1, 31) <= input(33);
output(1, 32) <= input(17);
output(1, 33) <= input(18);
output(1, 34) <= input(19);
output(1, 35) <= input(20);
output(1, 36) <= input(21);
output(1, 37) <= input(22);
output(1, 38) <= input(23);
output(1, 39) <= input(24);
output(1, 40) <= input(25);
output(1, 41) <= input(26);
output(1, 42) <= input(27);
output(1, 43) <= input(28);
output(1, 44) <= input(29);
output(1, 45) <= input(30);
output(1, 46) <= input(31);
output(1, 47) <= input(33);
output(1, 48) <= input(2);
output(1, 49) <= input(3);
output(1, 50) <= input(4);
output(1, 51) <= input(5);
output(1, 52) <= input(6);
output(1, 53) <= input(7);
output(1, 54) <= input(8);
output(1, 55) <= input(9);
output(1, 56) <= input(10);
output(1, 57) <= input(11);
output(1, 58) <= input(12);
output(1, 59) <= input(13);
output(1, 60) <= input(14);
output(1, 61) <= input(15);
output(1, 62) <= input(32);
output(1, 63) <= input(34);
output(1, 64) <= input(2);
output(1, 65) <= input(3);
output(1, 66) <= input(4);
output(1, 67) <= input(5);
output(1, 68) <= input(6);
output(1, 69) <= input(7);
output(1, 70) <= input(8);
output(1, 71) <= input(9);
output(1, 72) <= input(10);
output(1, 73) <= input(11);
output(1, 74) <= input(12);
output(1, 75) <= input(13);
output(1, 76) <= input(14);
output(1, 77) <= input(15);
output(1, 78) <= input(32);
output(1, 79) <= input(34);
output(1, 80) <= input(18);
output(1, 81) <= input(19);
output(1, 82) <= input(20);
output(1, 83) <= input(21);
output(1, 84) <= input(22);
output(1, 85) <= input(23);
output(1, 86) <= input(24);
output(1, 87) <= input(25);
output(1, 88) <= input(26);
output(1, 89) <= input(27);
output(1, 90) <= input(28);
output(1, 91) <= input(29);
output(1, 92) <= input(30);
output(1, 93) <= input(31);
output(1, 94) <= input(33);
output(1, 95) <= input(35);
output(1, 96) <= input(18);
output(1, 97) <= input(19);
output(1, 98) <= input(20);
output(1, 99) <= input(21);
output(1, 100) <= input(22);
output(1, 101) <= input(23);
output(1, 102) <= input(24);
output(1, 103) <= input(25);
output(1, 104) <= input(26);
output(1, 105) <= input(27);
output(1, 106) <= input(28);
output(1, 107) <= input(29);
output(1, 108) <= input(30);
output(1, 109) <= input(31);
output(1, 110) <= input(33);
output(1, 111) <= input(35);
output(1, 112) <= input(3);
output(1, 113) <= input(4);
output(1, 114) <= input(5);
output(1, 115) <= input(6);
output(1, 116) <= input(7);
output(1, 117) <= input(8);
output(1, 118) <= input(9);
output(1, 119) <= input(10);
output(1, 120) <= input(11);
output(1, 121) <= input(12);
output(1, 122) <= input(13);
output(1, 123) <= input(14);
output(1, 124) <= input(15);
output(1, 125) <= input(32);
output(1, 126) <= input(34);
output(1, 127) <= input(36);
output(1, 128) <= input(3);
output(1, 129) <= input(4);
output(1, 130) <= input(5);
output(1, 131) <= input(6);
output(1, 132) <= input(7);
output(1, 133) <= input(8);
output(1, 134) <= input(9);
output(1, 135) <= input(10);
output(1, 136) <= input(11);
output(1, 137) <= input(12);
output(1, 138) <= input(13);
output(1, 139) <= input(14);
output(1, 140) <= input(15);
output(1, 141) <= input(32);
output(1, 142) <= input(34);
output(1, 143) <= input(36);
output(1, 144) <= input(19);
output(1, 145) <= input(20);
output(1, 146) <= input(21);
output(1, 147) <= input(22);
output(1, 148) <= input(23);
output(1, 149) <= input(24);
output(1, 150) <= input(25);
output(1, 151) <= input(26);
output(1, 152) <= input(27);
output(1, 153) <= input(28);
output(1, 154) <= input(29);
output(1, 155) <= input(30);
output(1, 156) <= input(31);
output(1, 157) <= input(33);
output(1, 158) <= input(35);
output(1, 159) <= input(37);
output(1, 160) <= input(19);
output(1, 161) <= input(20);
output(1, 162) <= input(21);
output(1, 163) <= input(22);
output(1, 164) <= input(23);
output(1, 165) <= input(24);
output(1, 166) <= input(25);
output(1, 167) <= input(26);
output(1, 168) <= input(27);
output(1, 169) <= input(28);
output(1, 170) <= input(29);
output(1, 171) <= input(30);
output(1, 172) <= input(31);
output(1, 173) <= input(33);
output(1, 174) <= input(35);
output(1, 175) <= input(37);
output(1, 176) <= input(4);
output(1, 177) <= input(5);
output(1, 178) <= input(6);
output(1, 179) <= input(7);
output(1, 180) <= input(8);
output(1, 181) <= input(9);
output(1, 182) <= input(10);
output(1, 183) <= input(11);
output(1, 184) <= input(12);
output(1, 185) <= input(13);
output(1, 186) <= input(14);
output(1, 187) <= input(15);
output(1, 188) <= input(32);
output(1, 189) <= input(34);
output(1, 190) <= input(36);
output(1, 191) <= input(38);
output(1, 192) <= input(4);
output(1, 193) <= input(5);
output(1, 194) <= input(6);
output(1, 195) <= input(7);
output(1, 196) <= input(8);
output(1, 197) <= input(9);
output(1, 198) <= input(10);
output(1, 199) <= input(11);
output(1, 200) <= input(12);
output(1, 201) <= input(13);
output(1, 202) <= input(14);
output(1, 203) <= input(15);
output(1, 204) <= input(32);
output(1, 205) <= input(34);
output(1, 206) <= input(36);
output(1, 207) <= input(38);
output(1, 208) <= input(20);
output(1, 209) <= input(21);
output(1, 210) <= input(22);
output(1, 211) <= input(23);
output(1, 212) <= input(24);
output(1, 213) <= input(25);
output(1, 214) <= input(26);
output(1, 215) <= input(27);
output(1, 216) <= input(28);
output(1, 217) <= input(29);
output(1, 218) <= input(30);
output(1, 219) <= input(31);
output(1, 220) <= input(33);
output(1, 221) <= input(35);
output(1, 222) <= input(37);
output(1, 223) <= input(39);
output(1, 224) <= input(20);
output(1, 225) <= input(21);
output(1, 226) <= input(22);
output(1, 227) <= input(23);
output(1, 228) <= input(24);
output(1, 229) <= input(25);
output(1, 230) <= input(26);
output(1, 231) <= input(27);
output(1, 232) <= input(28);
output(1, 233) <= input(29);
output(1, 234) <= input(30);
output(1, 235) <= input(31);
output(1, 236) <= input(33);
output(1, 237) <= input(35);
output(1, 238) <= input(37);
output(1, 239) <= input(39);
output(1, 240) <= input(5);
output(1, 241) <= input(6);
output(1, 242) <= input(7);
output(1, 243) <= input(8);
output(1, 244) <= input(9);
output(1, 245) <= input(10);
output(1, 246) <= input(11);
output(1, 247) <= input(12);
output(1, 248) <= input(13);
output(1, 249) <= input(14);
output(1, 250) <= input(15);
output(1, 251) <= input(32);
output(1, 252) <= input(34);
output(1, 253) <= input(36);
output(1, 254) <= input(38);
output(1, 255) <= input(40);
output(2, 0) <= input(2);
output(2, 1) <= input(3);
output(2, 2) <= input(4);
output(2, 3) <= input(5);
output(2, 4) <= input(6);
output(2, 5) <= input(7);
output(2, 6) <= input(8);
output(2, 7) <= input(9);
output(2, 8) <= input(10);
output(2, 9) <= input(11);
output(2, 10) <= input(12);
output(2, 11) <= input(13);
output(2, 12) <= input(14);
output(2, 13) <= input(15);
output(2, 14) <= input(32);
output(2, 15) <= input(34);
output(2, 16) <= input(18);
output(2, 17) <= input(19);
output(2, 18) <= input(20);
output(2, 19) <= input(21);
output(2, 20) <= input(22);
output(2, 21) <= input(23);
output(2, 22) <= input(24);
output(2, 23) <= input(25);
output(2, 24) <= input(26);
output(2, 25) <= input(27);
output(2, 26) <= input(28);
output(2, 27) <= input(29);
output(2, 28) <= input(30);
output(2, 29) <= input(31);
output(2, 30) <= input(33);
output(2, 31) <= input(35);
output(2, 32) <= input(18);
output(2, 33) <= input(19);
output(2, 34) <= input(20);
output(2, 35) <= input(21);
output(2, 36) <= input(22);
output(2, 37) <= input(23);
output(2, 38) <= input(24);
output(2, 39) <= input(25);
output(2, 40) <= input(26);
output(2, 41) <= input(27);
output(2, 42) <= input(28);
output(2, 43) <= input(29);
output(2, 44) <= input(30);
output(2, 45) <= input(31);
output(2, 46) <= input(33);
output(2, 47) <= input(35);
output(2, 48) <= input(3);
output(2, 49) <= input(4);
output(2, 50) <= input(5);
output(2, 51) <= input(6);
output(2, 52) <= input(7);
output(2, 53) <= input(8);
output(2, 54) <= input(9);
output(2, 55) <= input(10);
output(2, 56) <= input(11);
output(2, 57) <= input(12);
output(2, 58) <= input(13);
output(2, 59) <= input(14);
output(2, 60) <= input(15);
output(2, 61) <= input(32);
output(2, 62) <= input(34);
output(2, 63) <= input(36);
output(2, 64) <= input(19);
output(2, 65) <= input(20);
output(2, 66) <= input(21);
output(2, 67) <= input(22);
output(2, 68) <= input(23);
output(2, 69) <= input(24);
output(2, 70) <= input(25);
output(2, 71) <= input(26);
output(2, 72) <= input(27);
output(2, 73) <= input(28);
output(2, 74) <= input(29);
output(2, 75) <= input(30);
output(2, 76) <= input(31);
output(2, 77) <= input(33);
output(2, 78) <= input(35);
output(2, 79) <= input(37);
output(2, 80) <= input(19);
output(2, 81) <= input(20);
output(2, 82) <= input(21);
output(2, 83) <= input(22);
output(2, 84) <= input(23);
output(2, 85) <= input(24);
output(2, 86) <= input(25);
output(2, 87) <= input(26);
output(2, 88) <= input(27);
output(2, 89) <= input(28);
output(2, 90) <= input(29);
output(2, 91) <= input(30);
output(2, 92) <= input(31);
output(2, 93) <= input(33);
output(2, 94) <= input(35);
output(2, 95) <= input(37);
output(2, 96) <= input(4);
output(2, 97) <= input(5);
output(2, 98) <= input(6);
output(2, 99) <= input(7);
output(2, 100) <= input(8);
output(2, 101) <= input(9);
output(2, 102) <= input(10);
output(2, 103) <= input(11);
output(2, 104) <= input(12);
output(2, 105) <= input(13);
output(2, 106) <= input(14);
output(2, 107) <= input(15);
output(2, 108) <= input(32);
output(2, 109) <= input(34);
output(2, 110) <= input(36);
output(2, 111) <= input(38);
output(2, 112) <= input(20);
output(2, 113) <= input(21);
output(2, 114) <= input(22);
output(2, 115) <= input(23);
output(2, 116) <= input(24);
output(2, 117) <= input(25);
output(2, 118) <= input(26);
output(2, 119) <= input(27);
output(2, 120) <= input(28);
output(2, 121) <= input(29);
output(2, 122) <= input(30);
output(2, 123) <= input(31);
output(2, 124) <= input(33);
output(2, 125) <= input(35);
output(2, 126) <= input(37);
output(2, 127) <= input(39);
output(2, 128) <= input(20);
output(2, 129) <= input(21);
output(2, 130) <= input(22);
output(2, 131) <= input(23);
output(2, 132) <= input(24);
output(2, 133) <= input(25);
output(2, 134) <= input(26);
output(2, 135) <= input(27);
output(2, 136) <= input(28);
output(2, 137) <= input(29);
output(2, 138) <= input(30);
output(2, 139) <= input(31);
output(2, 140) <= input(33);
output(2, 141) <= input(35);
output(2, 142) <= input(37);
output(2, 143) <= input(39);
output(2, 144) <= input(5);
output(2, 145) <= input(6);
output(2, 146) <= input(7);
output(2, 147) <= input(8);
output(2, 148) <= input(9);
output(2, 149) <= input(10);
output(2, 150) <= input(11);
output(2, 151) <= input(12);
output(2, 152) <= input(13);
output(2, 153) <= input(14);
output(2, 154) <= input(15);
output(2, 155) <= input(32);
output(2, 156) <= input(34);
output(2, 157) <= input(36);
output(2, 158) <= input(38);
output(2, 159) <= input(40);
output(2, 160) <= input(5);
output(2, 161) <= input(6);
output(2, 162) <= input(7);
output(2, 163) <= input(8);
output(2, 164) <= input(9);
output(2, 165) <= input(10);
output(2, 166) <= input(11);
output(2, 167) <= input(12);
output(2, 168) <= input(13);
output(2, 169) <= input(14);
output(2, 170) <= input(15);
output(2, 171) <= input(32);
output(2, 172) <= input(34);
output(2, 173) <= input(36);
output(2, 174) <= input(38);
output(2, 175) <= input(40);
output(2, 176) <= input(21);
output(2, 177) <= input(22);
output(2, 178) <= input(23);
output(2, 179) <= input(24);
output(2, 180) <= input(25);
output(2, 181) <= input(26);
output(2, 182) <= input(27);
output(2, 183) <= input(28);
output(2, 184) <= input(29);
output(2, 185) <= input(30);
output(2, 186) <= input(31);
output(2, 187) <= input(33);
output(2, 188) <= input(35);
output(2, 189) <= input(37);
output(2, 190) <= input(39);
output(2, 191) <= input(41);
output(2, 192) <= input(6);
output(2, 193) <= input(7);
output(2, 194) <= input(8);
output(2, 195) <= input(9);
output(2, 196) <= input(10);
output(2, 197) <= input(11);
output(2, 198) <= input(12);
output(2, 199) <= input(13);
output(2, 200) <= input(14);
output(2, 201) <= input(15);
output(2, 202) <= input(32);
output(2, 203) <= input(34);
output(2, 204) <= input(36);
output(2, 205) <= input(38);
output(2, 206) <= input(40);
output(2, 207) <= input(42);
output(2, 208) <= input(6);
output(2, 209) <= input(7);
output(2, 210) <= input(8);
output(2, 211) <= input(9);
output(2, 212) <= input(10);
output(2, 213) <= input(11);
output(2, 214) <= input(12);
output(2, 215) <= input(13);
output(2, 216) <= input(14);
output(2, 217) <= input(15);
output(2, 218) <= input(32);
output(2, 219) <= input(34);
output(2, 220) <= input(36);
output(2, 221) <= input(38);
output(2, 222) <= input(40);
output(2, 223) <= input(42);
output(2, 224) <= input(22);
output(2, 225) <= input(23);
output(2, 226) <= input(24);
output(2, 227) <= input(25);
output(2, 228) <= input(26);
output(2, 229) <= input(27);
output(2, 230) <= input(28);
output(2, 231) <= input(29);
output(2, 232) <= input(30);
output(2, 233) <= input(31);
output(2, 234) <= input(33);
output(2, 235) <= input(35);
output(2, 236) <= input(37);
output(2, 237) <= input(39);
output(2, 238) <= input(41);
output(2, 239) <= input(43);
output(2, 240) <= input(7);
output(2, 241) <= input(8);
output(2, 242) <= input(9);
output(2, 243) <= input(10);
output(2, 244) <= input(11);
output(2, 245) <= input(12);
output(2, 246) <= input(13);
output(2, 247) <= input(14);
output(2, 248) <= input(15);
output(2, 249) <= input(32);
output(2, 250) <= input(34);
output(2, 251) <= input(36);
output(2, 252) <= input(38);
output(2, 253) <= input(40);
output(2, 254) <= input(42);
output(2, 255) <= input(44);
output(3, 0) <= input(3);
output(3, 1) <= input(4);
output(3, 2) <= input(5);
output(3, 3) <= input(6);
output(3, 4) <= input(7);
output(3, 5) <= input(8);
output(3, 6) <= input(9);
output(3, 7) <= input(10);
output(3, 8) <= input(11);
output(3, 9) <= input(12);
output(3, 10) <= input(13);
output(3, 11) <= input(14);
output(3, 12) <= input(15);
output(3, 13) <= input(32);
output(3, 14) <= input(34);
output(3, 15) <= input(36);
output(3, 16) <= input(19);
output(3, 17) <= input(20);
output(3, 18) <= input(21);
output(3, 19) <= input(22);
output(3, 20) <= input(23);
output(3, 21) <= input(24);
output(3, 22) <= input(25);
output(3, 23) <= input(26);
output(3, 24) <= input(27);
output(3, 25) <= input(28);
output(3, 26) <= input(29);
output(3, 27) <= input(30);
output(3, 28) <= input(31);
output(3, 29) <= input(33);
output(3, 30) <= input(35);
output(3, 31) <= input(37);
output(3, 32) <= input(4);
output(3, 33) <= input(5);
output(3, 34) <= input(6);
output(3, 35) <= input(7);
output(3, 36) <= input(8);
output(3, 37) <= input(9);
output(3, 38) <= input(10);
output(3, 39) <= input(11);
output(3, 40) <= input(12);
output(3, 41) <= input(13);
output(3, 42) <= input(14);
output(3, 43) <= input(15);
output(3, 44) <= input(32);
output(3, 45) <= input(34);
output(3, 46) <= input(36);
output(3, 47) <= input(38);
output(3, 48) <= input(20);
output(3, 49) <= input(21);
output(3, 50) <= input(22);
output(3, 51) <= input(23);
output(3, 52) <= input(24);
output(3, 53) <= input(25);
output(3, 54) <= input(26);
output(3, 55) <= input(27);
output(3, 56) <= input(28);
output(3, 57) <= input(29);
output(3, 58) <= input(30);
output(3, 59) <= input(31);
output(3, 60) <= input(33);
output(3, 61) <= input(35);
output(3, 62) <= input(37);
output(3, 63) <= input(39);
output(3, 64) <= input(20);
output(3, 65) <= input(21);
output(3, 66) <= input(22);
output(3, 67) <= input(23);
output(3, 68) <= input(24);
output(3, 69) <= input(25);
output(3, 70) <= input(26);
output(3, 71) <= input(27);
output(3, 72) <= input(28);
output(3, 73) <= input(29);
output(3, 74) <= input(30);
output(3, 75) <= input(31);
output(3, 76) <= input(33);
output(3, 77) <= input(35);
output(3, 78) <= input(37);
output(3, 79) <= input(39);
output(3, 80) <= input(5);
output(3, 81) <= input(6);
output(3, 82) <= input(7);
output(3, 83) <= input(8);
output(3, 84) <= input(9);
output(3, 85) <= input(10);
output(3, 86) <= input(11);
output(3, 87) <= input(12);
output(3, 88) <= input(13);
output(3, 89) <= input(14);
output(3, 90) <= input(15);
output(3, 91) <= input(32);
output(3, 92) <= input(34);
output(3, 93) <= input(36);
output(3, 94) <= input(38);
output(3, 95) <= input(40);
output(3, 96) <= input(21);
output(3, 97) <= input(22);
output(3, 98) <= input(23);
output(3, 99) <= input(24);
output(3, 100) <= input(25);
output(3, 101) <= input(26);
output(3, 102) <= input(27);
output(3, 103) <= input(28);
output(3, 104) <= input(29);
output(3, 105) <= input(30);
output(3, 106) <= input(31);
output(3, 107) <= input(33);
output(3, 108) <= input(35);
output(3, 109) <= input(37);
output(3, 110) <= input(39);
output(3, 111) <= input(41);
output(3, 112) <= input(6);
output(3, 113) <= input(7);
output(3, 114) <= input(8);
output(3, 115) <= input(9);
output(3, 116) <= input(10);
output(3, 117) <= input(11);
output(3, 118) <= input(12);
output(3, 119) <= input(13);
output(3, 120) <= input(14);
output(3, 121) <= input(15);
output(3, 122) <= input(32);
output(3, 123) <= input(34);
output(3, 124) <= input(36);
output(3, 125) <= input(38);
output(3, 126) <= input(40);
output(3, 127) <= input(42);
output(3, 128) <= input(6);
output(3, 129) <= input(7);
output(3, 130) <= input(8);
output(3, 131) <= input(9);
output(3, 132) <= input(10);
output(3, 133) <= input(11);
output(3, 134) <= input(12);
output(3, 135) <= input(13);
output(3, 136) <= input(14);
output(3, 137) <= input(15);
output(3, 138) <= input(32);
output(3, 139) <= input(34);
output(3, 140) <= input(36);
output(3, 141) <= input(38);
output(3, 142) <= input(40);
output(3, 143) <= input(42);
output(3, 144) <= input(22);
output(3, 145) <= input(23);
output(3, 146) <= input(24);
output(3, 147) <= input(25);
output(3, 148) <= input(26);
output(3, 149) <= input(27);
output(3, 150) <= input(28);
output(3, 151) <= input(29);
output(3, 152) <= input(30);
output(3, 153) <= input(31);
output(3, 154) <= input(33);
output(3, 155) <= input(35);
output(3, 156) <= input(37);
output(3, 157) <= input(39);
output(3, 158) <= input(41);
output(3, 159) <= input(43);
output(3, 160) <= input(7);
output(3, 161) <= input(8);
output(3, 162) <= input(9);
output(3, 163) <= input(10);
output(3, 164) <= input(11);
output(3, 165) <= input(12);
output(3, 166) <= input(13);
output(3, 167) <= input(14);
output(3, 168) <= input(15);
output(3, 169) <= input(32);
output(3, 170) <= input(34);
output(3, 171) <= input(36);
output(3, 172) <= input(38);
output(3, 173) <= input(40);
output(3, 174) <= input(42);
output(3, 175) <= input(44);
output(3, 176) <= input(23);
output(3, 177) <= input(24);
output(3, 178) <= input(25);
output(3, 179) <= input(26);
output(3, 180) <= input(27);
output(3, 181) <= input(28);
output(3, 182) <= input(29);
output(3, 183) <= input(30);
output(3, 184) <= input(31);
output(3, 185) <= input(33);
output(3, 186) <= input(35);
output(3, 187) <= input(37);
output(3, 188) <= input(39);
output(3, 189) <= input(41);
output(3, 190) <= input(43);
output(3, 191) <= input(45);
output(3, 192) <= input(23);
output(3, 193) <= input(24);
output(3, 194) <= input(25);
output(3, 195) <= input(26);
output(3, 196) <= input(27);
output(3, 197) <= input(28);
output(3, 198) <= input(29);
output(3, 199) <= input(30);
output(3, 200) <= input(31);
output(3, 201) <= input(33);
output(3, 202) <= input(35);
output(3, 203) <= input(37);
output(3, 204) <= input(39);
output(3, 205) <= input(41);
output(3, 206) <= input(43);
output(3, 207) <= input(45);
output(3, 208) <= input(8);
output(3, 209) <= input(9);
output(3, 210) <= input(10);
output(3, 211) <= input(11);
output(3, 212) <= input(12);
output(3, 213) <= input(13);
output(3, 214) <= input(14);
output(3, 215) <= input(15);
output(3, 216) <= input(32);
output(3, 217) <= input(34);
output(3, 218) <= input(36);
output(3, 219) <= input(38);
output(3, 220) <= input(40);
output(3, 221) <= input(42);
output(3, 222) <= input(44);
output(3, 223) <= input(46);
output(3, 224) <= input(24);
output(3, 225) <= input(25);
output(3, 226) <= input(26);
output(3, 227) <= input(27);
output(3, 228) <= input(28);
output(3, 229) <= input(29);
output(3, 230) <= input(30);
output(3, 231) <= input(31);
output(3, 232) <= input(33);
output(3, 233) <= input(35);
output(3, 234) <= input(37);
output(3, 235) <= input(39);
output(3, 236) <= input(41);
output(3, 237) <= input(43);
output(3, 238) <= input(45);
output(3, 239) <= input(47);
output(3, 240) <= input(9);
output(3, 241) <= input(10);
output(3, 242) <= input(11);
output(3, 243) <= input(12);
output(3, 244) <= input(13);
output(3, 245) <= input(14);
output(3, 246) <= input(15);
output(3, 247) <= input(32);
output(3, 248) <= input(34);
output(3, 249) <= input(36);
output(3, 250) <= input(38);
output(3, 251) <= input(40);
output(3, 252) <= input(42);
output(3, 253) <= input(44);
output(3, 254) <= input(46);
output(3, 255) <= input(48);
output(4, 0) <= input(4);
output(4, 1) <= input(5);
output(4, 2) <= input(6);
output(4, 3) <= input(7);
output(4, 4) <= input(8);
output(4, 5) <= input(9);
output(4, 6) <= input(10);
output(4, 7) <= input(11);
output(4, 8) <= input(12);
output(4, 9) <= input(13);
output(4, 10) <= input(14);
output(4, 11) <= input(15);
output(4, 12) <= input(32);
output(4, 13) <= input(34);
output(4, 14) <= input(36);
output(4, 15) <= input(38);
output(4, 16) <= input(20);
output(4, 17) <= input(21);
output(4, 18) <= input(22);
output(4, 19) <= input(23);
output(4, 20) <= input(24);
output(4, 21) <= input(25);
output(4, 22) <= input(26);
output(4, 23) <= input(27);
output(4, 24) <= input(28);
output(4, 25) <= input(29);
output(4, 26) <= input(30);
output(4, 27) <= input(31);
output(4, 28) <= input(33);
output(4, 29) <= input(35);
output(4, 30) <= input(37);
output(4, 31) <= input(39);
output(4, 32) <= input(5);
output(4, 33) <= input(6);
output(4, 34) <= input(7);
output(4, 35) <= input(8);
output(4, 36) <= input(9);
output(4, 37) <= input(10);
output(4, 38) <= input(11);
output(4, 39) <= input(12);
output(4, 40) <= input(13);
output(4, 41) <= input(14);
output(4, 42) <= input(15);
output(4, 43) <= input(32);
output(4, 44) <= input(34);
output(4, 45) <= input(36);
output(4, 46) <= input(38);
output(4, 47) <= input(40);
output(4, 48) <= input(21);
output(4, 49) <= input(22);
output(4, 50) <= input(23);
output(4, 51) <= input(24);
output(4, 52) <= input(25);
output(4, 53) <= input(26);
output(4, 54) <= input(27);
output(4, 55) <= input(28);
output(4, 56) <= input(29);
output(4, 57) <= input(30);
output(4, 58) <= input(31);
output(4, 59) <= input(33);
output(4, 60) <= input(35);
output(4, 61) <= input(37);
output(4, 62) <= input(39);
output(4, 63) <= input(41);
output(4, 64) <= input(6);
output(4, 65) <= input(7);
output(4, 66) <= input(8);
output(4, 67) <= input(9);
output(4, 68) <= input(10);
output(4, 69) <= input(11);
output(4, 70) <= input(12);
output(4, 71) <= input(13);
output(4, 72) <= input(14);
output(4, 73) <= input(15);
output(4, 74) <= input(32);
output(4, 75) <= input(34);
output(4, 76) <= input(36);
output(4, 77) <= input(38);
output(4, 78) <= input(40);
output(4, 79) <= input(42);
output(4, 80) <= input(22);
output(4, 81) <= input(23);
output(4, 82) <= input(24);
output(4, 83) <= input(25);
output(4, 84) <= input(26);
output(4, 85) <= input(27);
output(4, 86) <= input(28);
output(4, 87) <= input(29);
output(4, 88) <= input(30);
output(4, 89) <= input(31);
output(4, 90) <= input(33);
output(4, 91) <= input(35);
output(4, 92) <= input(37);
output(4, 93) <= input(39);
output(4, 94) <= input(41);
output(4, 95) <= input(43);
output(4, 96) <= input(7);
output(4, 97) <= input(8);
output(4, 98) <= input(9);
output(4, 99) <= input(10);
output(4, 100) <= input(11);
output(4, 101) <= input(12);
output(4, 102) <= input(13);
output(4, 103) <= input(14);
output(4, 104) <= input(15);
output(4, 105) <= input(32);
output(4, 106) <= input(34);
output(4, 107) <= input(36);
output(4, 108) <= input(38);
output(4, 109) <= input(40);
output(4, 110) <= input(42);
output(4, 111) <= input(44);
output(4, 112) <= input(23);
output(4, 113) <= input(24);
output(4, 114) <= input(25);
output(4, 115) <= input(26);
output(4, 116) <= input(27);
output(4, 117) <= input(28);
output(4, 118) <= input(29);
output(4, 119) <= input(30);
output(4, 120) <= input(31);
output(4, 121) <= input(33);
output(4, 122) <= input(35);
output(4, 123) <= input(37);
output(4, 124) <= input(39);
output(4, 125) <= input(41);
output(4, 126) <= input(43);
output(4, 127) <= input(45);
output(4, 128) <= input(23);
output(4, 129) <= input(24);
output(4, 130) <= input(25);
output(4, 131) <= input(26);
output(4, 132) <= input(27);
output(4, 133) <= input(28);
output(4, 134) <= input(29);
output(4, 135) <= input(30);
output(4, 136) <= input(31);
output(4, 137) <= input(33);
output(4, 138) <= input(35);
output(4, 139) <= input(37);
output(4, 140) <= input(39);
output(4, 141) <= input(41);
output(4, 142) <= input(43);
output(4, 143) <= input(45);
output(4, 144) <= input(8);
output(4, 145) <= input(9);
output(4, 146) <= input(10);
output(4, 147) <= input(11);
output(4, 148) <= input(12);
output(4, 149) <= input(13);
output(4, 150) <= input(14);
output(4, 151) <= input(15);
output(4, 152) <= input(32);
output(4, 153) <= input(34);
output(4, 154) <= input(36);
output(4, 155) <= input(38);
output(4, 156) <= input(40);
output(4, 157) <= input(42);
output(4, 158) <= input(44);
output(4, 159) <= input(46);
output(4, 160) <= input(24);
output(4, 161) <= input(25);
output(4, 162) <= input(26);
output(4, 163) <= input(27);
output(4, 164) <= input(28);
output(4, 165) <= input(29);
output(4, 166) <= input(30);
output(4, 167) <= input(31);
output(4, 168) <= input(33);
output(4, 169) <= input(35);
output(4, 170) <= input(37);
output(4, 171) <= input(39);
output(4, 172) <= input(41);
output(4, 173) <= input(43);
output(4, 174) <= input(45);
output(4, 175) <= input(47);
output(4, 176) <= input(9);
output(4, 177) <= input(10);
output(4, 178) <= input(11);
output(4, 179) <= input(12);
output(4, 180) <= input(13);
output(4, 181) <= input(14);
output(4, 182) <= input(15);
output(4, 183) <= input(32);
output(4, 184) <= input(34);
output(4, 185) <= input(36);
output(4, 186) <= input(38);
output(4, 187) <= input(40);
output(4, 188) <= input(42);
output(4, 189) <= input(44);
output(4, 190) <= input(46);
output(4, 191) <= input(48);
output(4, 192) <= input(25);
output(4, 193) <= input(26);
output(4, 194) <= input(27);
output(4, 195) <= input(28);
output(4, 196) <= input(29);
output(4, 197) <= input(30);
output(4, 198) <= input(31);
output(4, 199) <= input(33);
output(4, 200) <= input(35);
output(4, 201) <= input(37);
output(4, 202) <= input(39);
output(4, 203) <= input(41);
output(4, 204) <= input(43);
output(4, 205) <= input(45);
output(4, 206) <= input(47);
output(4, 207) <= input(49);
output(4, 208) <= input(10);
output(4, 209) <= input(11);
output(4, 210) <= input(12);
output(4, 211) <= input(13);
output(4, 212) <= input(14);
output(4, 213) <= input(15);
output(4, 214) <= input(32);
output(4, 215) <= input(34);
output(4, 216) <= input(36);
output(4, 217) <= input(38);
output(4, 218) <= input(40);
output(4, 219) <= input(42);
output(4, 220) <= input(44);
output(4, 221) <= input(46);
output(4, 222) <= input(48);
output(4, 223) <= input(50);
output(4, 224) <= input(26);
output(4, 225) <= input(27);
output(4, 226) <= input(28);
output(4, 227) <= input(29);
output(4, 228) <= input(30);
output(4, 229) <= input(31);
output(4, 230) <= input(33);
output(4, 231) <= input(35);
output(4, 232) <= input(37);
output(4, 233) <= input(39);
output(4, 234) <= input(41);
output(4, 235) <= input(43);
output(4, 236) <= input(45);
output(4, 237) <= input(47);
output(4, 238) <= input(49);
output(4, 239) <= input(51);
output(4, 240) <= input(11);
output(4, 241) <= input(12);
output(4, 242) <= input(13);
output(4, 243) <= input(14);
output(4, 244) <= input(15);
output(4, 245) <= input(32);
output(4, 246) <= input(34);
output(4, 247) <= input(36);
output(4, 248) <= input(38);
output(4, 249) <= input(40);
output(4, 250) <= input(42);
output(4, 251) <= input(44);
output(4, 252) <= input(46);
output(4, 253) <= input(48);
output(4, 254) <= input(50);
output(4, 255) <= input(52);
output(5, 0) <= input(21);
output(5, 1) <= input(22);
output(5, 2) <= input(23);
output(5, 3) <= input(24);
output(5, 4) <= input(25);
output(5, 5) <= input(26);
output(5, 6) <= input(27);
output(5, 7) <= input(28);
output(5, 8) <= input(29);
output(5, 9) <= input(30);
output(5, 10) <= input(31);
output(5, 11) <= input(33);
output(5, 12) <= input(35);
output(5, 13) <= input(37);
output(5, 14) <= input(39);
output(5, 15) <= input(41);
output(5, 16) <= input(6);
output(5, 17) <= input(7);
output(5, 18) <= input(8);
output(5, 19) <= input(9);
output(5, 20) <= input(10);
output(5, 21) <= input(11);
output(5, 22) <= input(12);
output(5, 23) <= input(13);
output(5, 24) <= input(14);
output(5, 25) <= input(15);
output(5, 26) <= input(32);
output(5, 27) <= input(34);
output(5, 28) <= input(36);
output(5, 29) <= input(38);
output(5, 30) <= input(40);
output(5, 31) <= input(42);
output(5, 32) <= input(22);
output(5, 33) <= input(23);
output(5, 34) <= input(24);
output(5, 35) <= input(25);
output(5, 36) <= input(26);
output(5, 37) <= input(27);
output(5, 38) <= input(28);
output(5, 39) <= input(29);
output(5, 40) <= input(30);
output(5, 41) <= input(31);
output(5, 42) <= input(33);
output(5, 43) <= input(35);
output(5, 44) <= input(37);
output(5, 45) <= input(39);
output(5, 46) <= input(41);
output(5, 47) <= input(43);
output(5, 48) <= input(7);
output(5, 49) <= input(8);
output(5, 50) <= input(9);
output(5, 51) <= input(10);
output(5, 52) <= input(11);
output(5, 53) <= input(12);
output(5, 54) <= input(13);
output(5, 55) <= input(14);
output(5, 56) <= input(15);
output(5, 57) <= input(32);
output(5, 58) <= input(34);
output(5, 59) <= input(36);
output(5, 60) <= input(38);
output(5, 61) <= input(40);
output(5, 62) <= input(42);
output(5, 63) <= input(44);
output(5, 64) <= input(23);
output(5, 65) <= input(24);
output(5, 66) <= input(25);
output(5, 67) <= input(26);
output(5, 68) <= input(27);
output(5, 69) <= input(28);
output(5, 70) <= input(29);
output(5, 71) <= input(30);
output(5, 72) <= input(31);
output(5, 73) <= input(33);
output(5, 74) <= input(35);
output(5, 75) <= input(37);
output(5, 76) <= input(39);
output(5, 77) <= input(41);
output(5, 78) <= input(43);
output(5, 79) <= input(45);
output(5, 80) <= input(8);
output(5, 81) <= input(9);
output(5, 82) <= input(10);
output(5, 83) <= input(11);
output(5, 84) <= input(12);
output(5, 85) <= input(13);
output(5, 86) <= input(14);
output(5, 87) <= input(15);
output(5, 88) <= input(32);
output(5, 89) <= input(34);
output(5, 90) <= input(36);
output(5, 91) <= input(38);
output(5, 92) <= input(40);
output(5, 93) <= input(42);
output(5, 94) <= input(44);
output(5, 95) <= input(46);
output(5, 96) <= input(24);
output(5, 97) <= input(25);
output(5, 98) <= input(26);
output(5, 99) <= input(27);
output(5, 100) <= input(28);
output(5, 101) <= input(29);
output(5, 102) <= input(30);
output(5, 103) <= input(31);
output(5, 104) <= input(33);
output(5, 105) <= input(35);
output(5, 106) <= input(37);
output(5, 107) <= input(39);
output(5, 108) <= input(41);
output(5, 109) <= input(43);
output(5, 110) <= input(45);
output(5, 111) <= input(47);
output(5, 112) <= input(9);
output(5, 113) <= input(10);
output(5, 114) <= input(11);
output(5, 115) <= input(12);
output(5, 116) <= input(13);
output(5, 117) <= input(14);
output(5, 118) <= input(15);
output(5, 119) <= input(32);
output(5, 120) <= input(34);
output(5, 121) <= input(36);
output(5, 122) <= input(38);
output(5, 123) <= input(40);
output(5, 124) <= input(42);
output(5, 125) <= input(44);
output(5, 126) <= input(46);
output(5, 127) <= input(48);
output(5, 128) <= input(25);
output(5, 129) <= input(26);
output(5, 130) <= input(27);
output(5, 131) <= input(28);
output(5, 132) <= input(29);
output(5, 133) <= input(30);
output(5, 134) <= input(31);
output(5, 135) <= input(33);
output(5, 136) <= input(35);
output(5, 137) <= input(37);
output(5, 138) <= input(39);
output(5, 139) <= input(41);
output(5, 140) <= input(43);
output(5, 141) <= input(45);
output(5, 142) <= input(47);
output(5, 143) <= input(49);
output(5, 144) <= input(10);
output(5, 145) <= input(11);
output(5, 146) <= input(12);
output(5, 147) <= input(13);
output(5, 148) <= input(14);
output(5, 149) <= input(15);
output(5, 150) <= input(32);
output(5, 151) <= input(34);
output(5, 152) <= input(36);
output(5, 153) <= input(38);
output(5, 154) <= input(40);
output(5, 155) <= input(42);
output(5, 156) <= input(44);
output(5, 157) <= input(46);
output(5, 158) <= input(48);
output(5, 159) <= input(50);
output(5, 160) <= input(26);
output(5, 161) <= input(27);
output(5, 162) <= input(28);
output(5, 163) <= input(29);
output(5, 164) <= input(30);
output(5, 165) <= input(31);
output(5, 166) <= input(33);
output(5, 167) <= input(35);
output(5, 168) <= input(37);
output(5, 169) <= input(39);
output(5, 170) <= input(41);
output(5, 171) <= input(43);
output(5, 172) <= input(45);
output(5, 173) <= input(47);
output(5, 174) <= input(49);
output(5, 175) <= input(51);
output(5, 176) <= input(11);
output(5, 177) <= input(12);
output(5, 178) <= input(13);
output(5, 179) <= input(14);
output(5, 180) <= input(15);
output(5, 181) <= input(32);
output(5, 182) <= input(34);
output(5, 183) <= input(36);
output(5, 184) <= input(38);
output(5, 185) <= input(40);
output(5, 186) <= input(42);
output(5, 187) <= input(44);
output(5, 188) <= input(46);
output(5, 189) <= input(48);
output(5, 190) <= input(50);
output(5, 191) <= input(52);
output(5, 192) <= input(27);
output(5, 193) <= input(28);
output(5, 194) <= input(29);
output(5, 195) <= input(30);
output(5, 196) <= input(31);
output(5, 197) <= input(33);
output(5, 198) <= input(35);
output(5, 199) <= input(37);
output(5, 200) <= input(39);
output(5, 201) <= input(41);
output(5, 202) <= input(43);
output(5, 203) <= input(45);
output(5, 204) <= input(47);
output(5, 205) <= input(49);
output(5, 206) <= input(51);
output(5, 207) <= input(53);
output(5, 208) <= input(12);
output(5, 209) <= input(13);
output(5, 210) <= input(14);
output(5, 211) <= input(15);
output(5, 212) <= input(32);
output(5, 213) <= input(34);
output(5, 214) <= input(36);
output(5, 215) <= input(38);
output(5, 216) <= input(40);
output(5, 217) <= input(42);
output(5, 218) <= input(44);
output(5, 219) <= input(46);
output(5, 220) <= input(48);
output(5, 221) <= input(50);
output(5, 222) <= input(52);
output(5, 223) <= input(54);
output(5, 224) <= input(28);
output(5, 225) <= input(29);
output(5, 226) <= input(30);
output(5, 227) <= input(31);
output(5, 228) <= input(33);
output(5, 229) <= input(35);
output(5, 230) <= input(37);
output(5, 231) <= input(39);
output(5, 232) <= input(41);
output(5, 233) <= input(43);
output(5, 234) <= input(45);
output(5, 235) <= input(47);
output(5, 236) <= input(49);
output(5, 237) <= input(51);
output(5, 238) <= input(53);
output(5, 239) <= input(55);
output(5, 240) <= input(13);
output(5, 241) <= input(14);
output(5, 242) <= input(15);
output(5, 243) <= input(32);
output(5, 244) <= input(34);
output(5, 245) <= input(36);
output(5, 246) <= input(38);
output(5, 247) <= input(40);
output(5, 248) <= input(42);
output(5, 249) <= input(44);
output(5, 250) <= input(46);
output(5, 251) <= input(48);
output(5, 252) <= input(50);
output(5, 253) <= input(52);
output(5, 254) <= input(54);
output(5, 255) <= input(56);
when "1111" =>
output(0, 0) <= input(0);
output(0, 1) <= input(1);
output(0, 2) <= input(2);
output(0, 3) <= input(3);
output(0, 4) <= input(4);
output(0, 5) <= input(5);
output(0, 6) <= input(6);
output(0, 7) <= input(7);
output(0, 8) <= input(8);
output(0, 9) <= input(9);
output(0, 10) <= input(10);
output(0, 11) <= input(11);
output(0, 12) <= input(12);
output(0, 13) <= input(13);
output(0, 14) <= input(14);
output(0, 15) <= input(15);
output(0, 16) <= input(16);
output(0, 17) <= input(17);
output(0, 18) <= input(18);
output(0, 19) <= input(19);
output(0, 20) <= input(20);
output(0, 21) <= input(21);
output(0, 22) <= input(22);
output(0, 23) <= input(23);
output(0, 24) <= input(24);
output(0, 25) <= input(25);
output(0, 26) <= input(26);
output(0, 27) <= input(27);
output(0, 28) <= input(28);
output(0, 29) <= input(29);
output(0, 30) <= input(30);
output(0, 31) <= input(31);
output(0, 32) <= input(1);
output(0, 33) <= input(2);
output(0, 34) <= input(3);
output(0, 35) <= input(4);
output(0, 36) <= input(5);
output(0, 37) <= input(6);
output(0, 38) <= input(7);
output(0, 39) <= input(8);
output(0, 40) <= input(9);
output(0, 41) <= input(10);
output(0, 42) <= input(11);
output(0, 43) <= input(12);
output(0, 44) <= input(13);
output(0, 45) <= input(14);
output(0, 46) <= input(15);
output(0, 47) <= input(32);
output(0, 48) <= input(17);
output(0, 49) <= input(18);
output(0, 50) <= input(19);
output(0, 51) <= input(20);
output(0, 52) <= input(21);
output(0, 53) <= input(22);
output(0, 54) <= input(23);
output(0, 55) <= input(24);
output(0, 56) <= input(25);
output(0, 57) <= input(26);
output(0, 58) <= input(27);
output(0, 59) <= input(28);
output(0, 60) <= input(29);
output(0, 61) <= input(30);
output(0, 62) <= input(31);
output(0, 63) <= input(33);
output(0, 64) <= input(2);
output(0, 65) <= input(3);
output(0, 66) <= input(4);
output(0, 67) <= input(5);
output(0, 68) <= input(6);
output(0, 69) <= input(7);
output(0, 70) <= input(8);
output(0, 71) <= input(9);
output(0, 72) <= input(10);
output(0, 73) <= input(11);
output(0, 74) <= input(12);
output(0, 75) <= input(13);
output(0, 76) <= input(14);
output(0, 77) <= input(15);
output(0, 78) <= input(32);
output(0, 79) <= input(34);
output(0, 80) <= input(18);
output(0, 81) <= input(19);
output(0, 82) <= input(20);
output(0, 83) <= input(21);
output(0, 84) <= input(22);
output(0, 85) <= input(23);
output(0, 86) <= input(24);
output(0, 87) <= input(25);
output(0, 88) <= input(26);
output(0, 89) <= input(27);
output(0, 90) <= input(28);
output(0, 91) <= input(29);
output(0, 92) <= input(30);
output(0, 93) <= input(31);
output(0, 94) <= input(33);
output(0, 95) <= input(35);
output(0, 96) <= input(3);
output(0, 97) <= input(4);
output(0, 98) <= input(5);
output(0, 99) <= input(6);
output(0, 100) <= input(7);
output(0, 101) <= input(8);
output(0, 102) <= input(9);
output(0, 103) <= input(10);
output(0, 104) <= input(11);
output(0, 105) <= input(12);
output(0, 106) <= input(13);
output(0, 107) <= input(14);
output(0, 108) <= input(15);
output(0, 109) <= input(32);
output(0, 110) <= input(34);
output(0, 111) <= input(36);
output(0, 112) <= input(4);
output(0, 113) <= input(5);
output(0, 114) <= input(6);
output(0, 115) <= input(7);
output(0, 116) <= input(8);
output(0, 117) <= input(9);
output(0, 118) <= input(10);
output(0, 119) <= input(11);
output(0, 120) <= input(12);
output(0, 121) <= input(13);
output(0, 122) <= input(14);
output(0, 123) <= input(15);
output(0, 124) <= input(32);
output(0, 125) <= input(34);
output(0, 126) <= input(36);
output(0, 127) <= input(37);
output(0, 128) <= input(20);
output(0, 129) <= input(21);
output(0, 130) <= input(22);
output(0, 131) <= input(23);
output(0, 132) <= input(24);
output(0, 133) <= input(25);
output(0, 134) <= input(26);
output(0, 135) <= input(27);
output(0, 136) <= input(28);
output(0, 137) <= input(29);
output(0, 138) <= input(30);
output(0, 139) <= input(31);
output(0, 140) <= input(33);
output(0, 141) <= input(35);
output(0, 142) <= input(38);
output(0, 143) <= input(39);
output(0, 144) <= input(5);
output(0, 145) <= input(6);
output(0, 146) <= input(7);
output(0, 147) <= input(8);
output(0, 148) <= input(9);
output(0, 149) <= input(10);
output(0, 150) <= input(11);
output(0, 151) <= input(12);
output(0, 152) <= input(13);
output(0, 153) <= input(14);
output(0, 154) <= input(15);
output(0, 155) <= input(32);
output(0, 156) <= input(34);
output(0, 157) <= input(36);
output(0, 158) <= input(37);
output(0, 159) <= input(40);
output(0, 160) <= input(21);
output(0, 161) <= input(22);
output(0, 162) <= input(23);
output(0, 163) <= input(24);
output(0, 164) <= input(25);
output(0, 165) <= input(26);
output(0, 166) <= input(27);
output(0, 167) <= input(28);
output(0, 168) <= input(29);
output(0, 169) <= input(30);
output(0, 170) <= input(31);
output(0, 171) <= input(33);
output(0, 172) <= input(35);
output(0, 173) <= input(38);
output(0, 174) <= input(39);
output(0, 175) <= input(41);
output(0, 176) <= input(6);
output(0, 177) <= input(7);
output(0, 178) <= input(8);
output(0, 179) <= input(9);
output(0, 180) <= input(10);
output(0, 181) <= input(11);
output(0, 182) <= input(12);
output(0, 183) <= input(13);
output(0, 184) <= input(14);
output(0, 185) <= input(15);
output(0, 186) <= input(32);
output(0, 187) <= input(34);
output(0, 188) <= input(36);
output(0, 189) <= input(37);
output(0, 190) <= input(40);
output(0, 191) <= input(42);
output(0, 192) <= input(22);
output(0, 193) <= input(23);
output(0, 194) <= input(24);
output(0, 195) <= input(25);
output(0, 196) <= input(26);
output(0, 197) <= input(27);
output(0, 198) <= input(28);
output(0, 199) <= input(29);
output(0, 200) <= input(30);
output(0, 201) <= input(31);
output(0, 202) <= input(33);
output(0, 203) <= input(35);
output(0, 204) <= input(38);
output(0, 205) <= input(39);
output(0, 206) <= input(41);
output(0, 207) <= input(43);
output(0, 208) <= input(7);
output(0, 209) <= input(8);
output(0, 210) <= input(9);
output(0, 211) <= input(10);
output(0, 212) <= input(11);
output(0, 213) <= input(12);
output(0, 214) <= input(13);
output(0, 215) <= input(14);
output(0, 216) <= input(15);
output(0, 217) <= input(32);
output(0, 218) <= input(34);
output(0, 219) <= input(36);
output(0, 220) <= input(37);
output(0, 221) <= input(40);
output(0, 222) <= input(42);
output(0, 223) <= input(44);
output(0, 224) <= input(23);
output(0, 225) <= input(24);
output(0, 226) <= input(25);
output(0, 227) <= input(26);
output(0, 228) <= input(27);
output(0, 229) <= input(28);
output(0, 230) <= input(29);
output(0, 231) <= input(30);
output(0, 232) <= input(31);
output(0, 233) <= input(33);
output(0, 234) <= input(35);
output(0, 235) <= input(38);
output(0, 236) <= input(39);
output(0, 237) <= input(41);
output(0, 238) <= input(43);
output(0, 239) <= input(45);
output(0, 240) <= input(24);
output(0, 241) <= input(25);
output(0, 242) <= input(26);
output(0, 243) <= input(27);
output(0, 244) <= input(28);
output(0, 245) <= input(29);
output(0, 246) <= input(30);
output(0, 247) <= input(31);
output(0, 248) <= input(33);
output(0, 249) <= input(35);
output(0, 250) <= input(38);
output(0, 251) <= input(39);
output(0, 252) <= input(41);
output(0, 253) <= input(43);
output(0, 254) <= input(45);
output(0, 255) <= input(46);
output(1, 0) <= input(1);
output(1, 1) <= input(2);
output(1, 2) <= input(3);
output(1, 3) <= input(4);
output(1, 4) <= input(5);
output(1, 5) <= input(6);
output(1, 6) <= input(7);
output(1, 7) <= input(8);
output(1, 8) <= input(9);
output(1, 9) <= input(10);
output(1, 10) <= input(11);
output(1, 11) <= input(12);
output(1, 12) <= input(13);
output(1, 13) <= input(14);
output(1, 14) <= input(15);
output(1, 15) <= input(32);
output(1, 16) <= input(17);
output(1, 17) <= input(18);
output(1, 18) <= input(19);
output(1, 19) <= input(20);
output(1, 20) <= input(21);
output(1, 21) <= input(22);
output(1, 22) <= input(23);
output(1, 23) <= input(24);
output(1, 24) <= input(25);
output(1, 25) <= input(26);
output(1, 26) <= input(27);
output(1, 27) <= input(28);
output(1, 28) <= input(29);
output(1, 29) <= input(30);
output(1, 30) <= input(31);
output(1, 31) <= input(33);
output(1, 32) <= input(2);
output(1, 33) <= input(3);
output(1, 34) <= input(4);
output(1, 35) <= input(5);
output(1, 36) <= input(6);
output(1, 37) <= input(7);
output(1, 38) <= input(8);
output(1, 39) <= input(9);
output(1, 40) <= input(10);
output(1, 41) <= input(11);
output(1, 42) <= input(12);
output(1, 43) <= input(13);
output(1, 44) <= input(14);
output(1, 45) <= input(15);
output(1, 46) <= input(32);
output(1, 47) <= input(34);
output(1, 48) <= input(3);
output(1, 49) <= input(4);
output(1, 50) <= input(5);
output(1, 51) <= input(6);
output(1, 52) <= input(7);
output(1, 53) <= input(8);
output(1, 54) <= input(9);
output(1, 55) <= input(10);
output(1, 56) <= input(11);
output(1, 57) <= input(12);
output(1, 58) <= input(13);
output(1, 59) <= input(14);
output(1, 60) <= input(15);
output(1, 61) <= input(32);
output(1, 62) <= input(34);
output(1, 63) <= input(36);
output(1, 64) <= input(19);
output(1, 65) <= input(20);
output(1, 66) <= input(21);
output(1, 67) <= input(22);
output(1, 68) <= input(23);
output(1, 69) <= input(24);
output(1, 70) <= input(25);
output(1, 71) <= input(26);
output(1, 72) <= input(27);
output(1, 73) <= input(28);
output(1, 74) <= input(29);
output(1, 75) <= input(30);
output(1, 76) <= input(31);
output(1, 77) <= input(33);
output(1, 78) <= input(35);
output(1, 79) <= input(38);
output(1, 80) <= input(4);
output(1, 81) <= input(5);
output(1, 82) <= input(6);
output(1, 83) <= input(7);
output(1, 84) <= input(8);
output(1, 85) <= input(9);
output(1, 86) <= input(10);
output(1, 87) <= input(11);
output(1, 88) <= input(12);
output(1, 89) <= input(13);
output(1, 90) <= input(14);
output(1, 91) <= input(15);
output(1, 92) <= input(32);
output(1, 93) <= input(34);
output(1, 94) <= input(36);
output(1, 95) <= input(37);
output(1, 96) <= input(20);
output(1, 97) <= input(21);
output(1, 98) <= input(22);
output(1, 99) <= input(23);
output(1, 100) <= input(24);
output(1, 101) <= input(25);
output(1, 102) <= input(26);
output(1, 103) <= input(27);
output(1, 104) <= input(28);
output(1, 105) <= input(29);
output(1, 106) <= input(30);
output(1, 107) <= input(31);
output(1, 108) <= input(33);
output(1, 109) <= input(35);
output(1, 110) <= input(38);
output(1, 111) <= input(39);
output(1, 112) <= input(21);
output(1, 113) <= input(22);
output(1, 114) <= input(23);
output(1, 115) <= input(24);
output(1, 116) <= input(25);
output(1, 117) <= input(26);
output(1, 118) <= input(27);
output(1, 119) <= input(28);
output(1, 120) <= input(29);
output(1, 121) <= input(30);
output(1, 122) <= input(31);
output(1, 123) <= input(33);
output(1, 124) <= input(35);
output(1, 125) <= input(38);
output(1, 126) <= input(39);
output(1, 127) <= input(41);
output(1, 128) <= input(6);
output(1, 129) <= input(7);
output(1, 130) <= input(8);
output(1, 131) <= input(9);
output(1, 132) <= input(10);
output(1, 133) <= input(11);
output(1, 134) <= input(12);
output(1, 135) <= input(13);
output(1, 136) <= input(14);
output(1, 137) <= input(15);
output(1, 138) <= input(32);
output(1, 139) <= input(34);
output(1, 140) <= input(36);
output(1, 141) <= input(37);
output(1, 142) <= input(40);
output(1, 143) <= input(42);
output(1, 144) <= input(22);
output(1, 145) <= input(23);
output(1, 146) <= input(24);
output(1, 147) <= input(25);
output(1, 148) <= input(26);
output(1, 149) <= input(27);
output(1, 150) <= input(28);
output(1, 151) <= input(29);
output(1, 152) <= input(30);
output(1, 153) <= input(31);
output(1, 154) <= input(33);
output(1, 155) <= input(35);
output(1, 156) <= input(38);
output(1, 157) <= input(39);
output(1, 158) <= input(41);
output(1, 159) <= input(43);
output(1, 160) <= input(7);
output(1, 161) <= input(8);
output(1, 162) <= input(9);
output(1, 163) <= input(10);
output(1, 164) <= input(11);
output(1, 165) <= input(12);
output(1, 166) <= input(13);
output(1, 167) <= input(14);
output(1, 168) <= input(15);
output(1, 169) <= input(32);
output(1, 170) <= input(34);
output(1, 171) <= input(36);
output(1, 172) <= input(37);
output(1, 173) <= input(40);
output(1, 174) <= input(42);
output(1, 175) <= input(44);
output(1, 176) <= input(8);
output(1, 177) <= input(9);
output(1, 178) <= input(10);
output(1, 179) <= input(11);
output(1, 180) <= input(12);
output(1, 181) <= input(13);
output(1, 182) <= input(14);
output(1, 183) <= input(15);
output(1, 184) <= input(32);
output(1, 185) <= input(34);
output(1, 186) <= input(36);
output(1, 187) <= input(37);
output(1, 188) <= input(40);
output(1, 189) <= input(42);
output(1, 190) <= input(44);
output(1, 191) <= input(47);
output(1, 192) <= input(24);
output(1, 193) <= input(25);
output(1, 194) <= input(26);
output(1, 195) <= input(27);
output(1, 196) <= input(28);
output(1, 197) <= input(29);
output(1, 198) <= input(30);
output(1, 199) <= input(31);
output(1, 200) <= input(33);
output(1, 201) <= input(35);
output(1, 202) <= input(38);
output(1, 203) <= input(39);
output(1, 204) <= input(41);
output(1, 205) <= input(43);
output(1, 206) <= input(45);
output(1, 207) <= input(46);
output(1, 208) <= input(9);
output(1, 209) <= input(10);
output(1, 210) <= input(11);
output(1, 211) <= input(12);
output(1, 212) <= input(13);
output(1, 213) <= input(14);
output(1, 214) <= input(15);
output(1, 215) <= input(32);
output(1, 216) <= input(34);
output(1, 217) <= input(36);
output(1, 218) <= input(37);
output(1, 219) <= input(40);
output(1, 220) <= input(42);
output(1, 221) <= input(44);
output(1, 222) <= input(47);
output(1, 223) <= input(48);
output(1, 224) <= input(25);
output(1, 225) <= input(26);
output(1, 226) <= input(27);
output(1, 227) <= input(28);
output(1, 228) <= input(29);
output(1, 229) <= input(30);
output(1, 230) <= input(31);
output(1, 231) <= input(33);
output(1, 232) <= input(35);
output(1, 233) <= input(38);
output(1, 234) <= input(39);
output(1, 235) <= input(41);
output(1, 236) <= input(43);
output(1, 237) <= input(45);
output(1, 238) <= input(46);
output(1, 239) <= input(49);
output(1, 240) <= input(26);
output(1, 241) <= input(27);
output(1, 242) <= input(28);
output(1, 243) <= input(29);
output(1, 244) <= input(30);
output(1, 245) <= input(31);
output(1, 246) <= input(33);
output(1, 247) <= input(35);
output(1, 248) <= input(38);
output(1, 249) <= input(39);
output(1, 250) <= input(41);
output(1, 251) <= input(43);
output(1, 252) <= input(45);
output(1, 253) <= input(46);
output(1, 254) <= input(49);
output(1, 255) <= input(50);
output(2, 0) <= input(18);
output(2, 1) <= input(19);
output(2, 2) <= input(20);
output(2, 3) <= input(21);
output(2, 4) <= input(22);
output(2, 5) <= input(23);
output(2, 6) <= input(24);
output(2, 7) <= input(25);
output(2, 8) <= input(26);
output(2, 9) <= input(27);
output(2, 10) <= input(28);
output(2, 11) <= input(29);
output(2, 12) <= input(30);
output(2, 13) <= input(31);
output(2, 14) <= input(33);
output(2, 15) <= input(35);
output(2, 16) <= input(3);
output(2, 17) <= input(4);
output(2, 18) <= input(5);
output(2, 19) <= input(6);
output(2, 20) <= input(7);
output(2, 21) <= input(8);
output(2, 22) <= input(9);
output(2, 23) <= input(10);
output(2, 24) <= input(11);
output(2, 25) <= input(12);
output(2, 26) <= input(13);
output(2, 27) <= input(14);
output(2, 28) <= input(15);
output(2, 29) <= input(32);
output(2, 30) <= input(34);
output(2, 31) <= input(36);
output(2, 32) <= input(4);
output(2, 33) <= input(5);
output(2, 34) <= input(6);
output(2, 35) <= input(7);
output(2, 36) <= input(8);
output(2, 37) <= input(9);
output(2, 38) <= input(10);
output(2, 39) <= input(11);
output(2, 40) <= input(12);
output(2, 41) <= input(13);
output(2, 42) <= input(14);
output(2, 43) <= input(15);
output(2, 44) <= input(32);
output(2, 45) <= input(34);
output(2, 46) <= input(36);
output(2, 47) <= input(37);
output(2, 48) <= input(20);
output(2, 49) <= input(21);
output(2, 50) <= input(22);
output(2, 51) <= input(23);
output(2, 52) <= input(24);
output(2, 53) <= input(25);
output(2, 54) <= input(26);
output(2, 55) <= input(27);
output(2, 56) <= input(28);
output(2, 57) <= input(29);
output(2, 58) <= input(30);
output(2, 59) <= input(31);
output(2, 60) <= input(33);
output(2, 61) <= input(35);
output(2, 62) <= input(38);
output(2, 63) <= input(39);
output(2, 64) <= input(21);
output(2, 65) <= input(22);
output(2, 66) <= input(23);
output(2, 67) <= input(24);
output(2, 68) <= input(25);
output(2, 69) <= input(26);
output(2, 70) <= input(27);
output(2, 71) <= input(28);
output(2, 72) <= input(29);
output(2, 73) <= input(30);
output(2, 74) <= input(31);
output(2, 75) <= input(33);
output(2, 76) <= input(35);
output(2, 77) <= input(38);
output(2, 78) <= input(39);
output(2, 79) <= input(41);
output(2, 80) <= input(6);
output(2, 81) <= input(7);
output(2, 82) <= input(8);
output(2, 83) <= input(9);
output(2, 84) <= input(10);
output(2, 85) <= input(11);
output(2, 86) <= input(12);
output(2, 87) <= input(13);
output(2, 88) <= input(14);
output(2, 89) <= input(15);
output(2, 90) <= input(32);
output(2, 91) <= input(34);
output(2, 92) <= input(36);
output(2, 93) <= input(37);
output(2, 94) <= input(40);
output(2, 95) <= input(42);
output(2, 96) <= input(7);
output(2, 97) <= input(8);
output(2, 98) <= input(9);
output(2, 99) <= input(10);
output(2, 100) <= input(11);
output(2, 101) <= input(12);
output(2, 102) <= input(13);
output(2, 103) <= input(14);
output(2, 104) <= input(15);
output(2, 105) <= input(32);
output(2, 106) <= input(34);
output(2, 107) <= input(36);
output(2, 108) <= input(37);
output(2, 109) <= input(40);
output(2, 110) <= input(42);
output(2, 111) <= input(44);
output(2, 112) <= input(23);
output(2, 113) <= input(24);
output(2, 114) <= input(25);
output(2, 115) <= input(26);
output(2, 116) <= input(27);
output(2, 117) <= input(28);
output(2, 118) <= input(29);
output(2, 119) <= input(30);
output(2, 120) <= input(31);
output(2, 121) <= input(33);
output(2, 122) <= input(35);
output(2, 123) <= input(38);
output(2, 124) <= input(39);
output(2, 125) <= input(41);
output(2, 126) <= input(43);
output(2, 127) <= input(45);
output(2, 128) <= input(8);
output(2, 129) <= input(9);
output(2, 130) <= input(10);
output(2, 131) <= input(11);
output(2, 132) <= input(12);
output(2, 133) <= input(13);
output(2, 134) <= input(14);
output(2, 135) <= input(15);
output(2, 136) <= input(32);
output(2, 137) <= input(34);
output(2, 138) <= input(36);
output(2, 139) <= input(37);
output(2, 140) <= input(40);
output(2, 141) <= input(42);
output(2, 142) <= input(44);
output(2, 143) <= input(47);
output(2, 144) <= input(9);
output(2, 145) <= input(10);
output(2, 146) <= input(11);
output(2, 147) <= input(12);
output(2, 148) <= input(13);
output(2, 149) <= input(14);
output(2, 150) <= input(15);
output(2, 151) <= input(32);
output(2, 152) <= input(34);
output(2, 153) <= input(36);
output(2, 154) <= input(37);
output(2, 155) <= input(40);
output(2, 156) <= input(42);
output(2, 157) <= input(44);
output(2, 158) <= input(47);
output(2, 159) <= input(48);
output(2, 160) <= input(25);
output(2, 161) <= input(26);
output(2, 162) <= input(27);
output(2, 163) <= input(28);
output(2, 164) <= input(29);
output(2, 165) <= input(30);
output(2, 166) <= input(31);
output(2, 167) <= input(33);
output(2, 168) <= input(35);
output(2, 169) <= input(38);
output(2, 170) <= input(39);
output(2, 171) <= input(41);
output(2, 172) <= input(43);
output(2, 173) <= input(45);
output(2, 174) <= input(46);
output(2, 175) <= input(49);
output(2, 176) <= input(26);
output(2, 177) <= input(27);
output(2, 178) <= input(28);
output(2, 179) <= input(29);
output(2, 180) <= input(30);
output(2, 181) <= input(31);
output(2, 182) <= input(33);
output(2, 183) <= input(35);
output(2, 184) <= input(38);
output(2, 185) <= input(39);
output(2, 186) <= input(41);
output(2, 187) <= input(43);
output(2, 188) <= input(45);
output(2, 189) <= input(46);
output(2, 190) <= input(49);
output(2, 191) <= input(50);
output(2, 192) <= input(11);
output(2, 193) <= input(12);
output(2, 194) <= input(13);
output(2, 195) <= input(14);
output(2, 196) <= input(15);
output(2, 197) <= input(32);
output(2, 198) <= input(34);
output(2, 199) <= input(36);
output(2, 200) <= input(37);
output(2, 201) <= input(40);
output(2, 202) <= input(42);
output(2, 203) <= input(44);
output(2, 204) <= input(47);
output(2, 205) <= input(48);
output(2, 206) <= input(51);
output(2, 207) <= input(52);
output(2, 208) <= input(12);
output(2, 209) <= input(13);
output(2, 210) <= input(14);
output(2, 211) <= input(15);
output(2, 212) <= input(32);
output(2, 213) <= input(34);
output(2, 214) <= input(36);
output(2, 215) <= input(37);
output(2, 216) <= input(40);
output(2, 217) <= input(42);
output(2, 218) <= input(44);
output(2, 219) <= input(47);
output(2, 220) <= input(48);
output(2, 221) <= input(51);
output(2, 222) <= input(52);
output(2, 223) <= input(53);
output(2, 224) <= input(28);
output(2, 225) <= input(29);
output(2, 226) <= input(30);
output(2, 227) <= input(31);
output(2, 228) <= input(33);
output(2, 229) <= input(35);
output(2, 230) <= input(38);
output(2, 231) <= input(39);
output(2, 232) <= input(41);
output(2, 233) <= input(43);
output(2, 234) <= input(45);
output(2, 235) <= input(46);
output(2, 236) <= input(49);
output(2, 237) <= input(50);
output(2, 238) <= input(54);
output(2, 239) <= input(55);
output(2, 240) <= input(29);
output(2, 241) <= input(30);
output(2, 242) <= input(31);
output(2, 243) <= input(33);
output(2, 244) <= input(35);
output(2, 245) <= input(38);
output(2, 246) <= input(39);
output(2, 247) <= input(41);
output(2, 248) <= input(43);
output(2, 249) <= input(45);
output(2, 250) <= input(46);
output(2, 251) <= input(49);
output(2, 252) <= input(50);
output(2, 253) <= input(54);
output(2, 254) <= input(55);
output(2, 255) <= input(56);
output(3, 0) <= input(4);
output(3, 1) <= input(5);
output(3, 2) <= input(6);
output(3, 3) <= input(7);
output(3, 4) <= input(8);
output(3, 5) <= input(9);
output(3, 6) <= input(10);
output(3, 7) <= input(11);
output(3, 8) <= input(12);
output(3, 9) <= input(13);
output(3, 10) <= input(14);
output(3, 11) <= input(15);
output(3, 12) <= input(32);
output(3, 13) <= input(34);
output(3, 14) <= input(36);
output(3, 15) <= input(37);
output(3, 16) <= input(5);
output(3, 17) <= input(6);
output(3, 18) <= input(7);
output(3, 19) <= input(8);
output(3, 20) <= input(9);
output(3, 21) <= input(10);
output(3, 22) <= input(11);
output(3, 23) <= input(12);
output(3, 24) <= input(13);
output(3, 25) <= input(14);
output(3, 26) <= input(15);
output(3, 27) <= input(32);
output(3, 28) <= input(34);
output(3, 29) <= input(36);
output(3, 30) <= input(37);
output(3, 31) <= input(40);
output(3, 32) <= input(21);
output(3, 33) <= input(22);
output(3, 34) <= input(23);
output(3, 35) <= input(24);
output(3, 36) <= input(25);
output(3, 37) <= input(26);
output(3, 38) <= input(27);
output(3, 39) <= input(28);
output(3, 40) <= input(29);
output(3, 41) <= input(30);
output(3, 42) <= input(31);
output(3, 43) <= input(33);
output(3, 44) <= input(35);
output(3, 45) <= input(38);
output(3, 46) <= input(39);
output(3, 47) <= input(41);
output(3, 48) <= input(22);
output(3, 49) <= input(23);
output(3, 50) <= input(24);
output(3, 51) <= input(25);
output(3, 52) <= input(26);
output(3, 53) <= input(27);
output(3, 54) <= input(28);
output(3, 55) <= input(29);
output(3, 56) <= input(30);
output(3, 57) <= input(31);
output(3, 58) <= input(33);
output(3, 59) <= input(35);
output(3, 60) <= input(38);
output(3, 61) <= input(39);
output(3, 62) <= input(41);
output(3, 63) <= input(43);
output(3, 64) <= input(23);
output(3, 65) <= input(24);
output(3, 66) <= input(25);
output(3, 67) <= input(26);
output(3, 68) <= input(27);
output(3, 69) <= input(28);
output(3, 70) <= input(29);
output(3, 71) <= input(30);
output(3, 72) <= input(31);
output(3, 73) <= input(33);
output(3, 74) <= input(35);
output(3, 75) <= input(38);
output(3, 76) <= input(39);
output(3, 77) <= input(41);
output(3, 78) <= input(43);
output(3, 79) <= input(45);
output(3, 80) <= input(8);
output(3, 81) <= input(9);
output(3, 82) <= input(10);
output(3, 83) <= input(11);
output(3, 84) <= input(12);
output(3, 85) <= input(13);
output(3, 86) <= input(14);
output(3, 87) <= input(15);
output(3, 88) <= input(32);
output(3, 89) <= input(34);
output(3, 90) <= input(36);
output(3, 91) <= input(37);
output(3, 92) <= input(40);
output(3, 93) <= input(42);
output(3, 94) <= input(44);
output(3, 95) <= input(47);
output(3, 96) <= input(9);
output(3, 97) <= input(10);
output(3, 98) <= input(11);
output(3, 99) <= input(12);
output(3, 100) <= input(13);
output(3, 101) <= input(14);
output(3, 102) <= input(15);
output(3, 103) <= input(32);
output(3, 104) <= input(34);
output(3, 105) <= input(36);
output(3, 106) <= input(37);
output(3, 107) <= input(40);
output(3, 108) <= input(42);
output(3, 109) <= input(44);
output(3, 110) <= input(47);
output(3, 111) <= input(48);
output(3, 112) <= input(10);
output(3, 113) <= input(11);
output(3, 114) <= input(12);
output(3, 115) <= input(13);
output(3, 116) <= input(14);
output(3, 117) <= input(15);
output(3, 118) <= input(32);
output(3, 119) <= input(34);
output(3, 120) <= input(36);
output(3, 121) <= input(37);
output(3, 122) <= input(40);
output(3, 123) <= input(42);
output(3, 124) <= input(44);
output(3, 125) <= input(47);
output(3, 126) <= input(48);
output(3, 127) <= input(51);
output(3, 128) <= input(26);
output(3, 129) <= input(27);
output(3, 130) <= input(28);
output(3, 131) <= input(29);
output(3, 132) <= input(30);
output(3, 133) <= input(31);
output(3, 134) <= input(33);
output(3, 135) <= input(35);
output(3, 136) <= input(38);
output(3, 137) <= input(39);
output(3, 138) <= input(41);
output(3, 139) <= input(43);
output(3, 140) <= input(45);
output(3, 141) <= input(46);
output(3, 142) <= input(49);
output(3, 143) <= input(50);
output(3, 144) <= input(27);
output(3, 145) <= input(28);
output(3, 146) <= input(29);
output(3, 147) <= input(30);
output(3, 148) <= input(31);
output(3, 149) <= input(33);
output(3, 150) <= input(35);
output(3, 151) <= input(38);
output(3, 152) <= input(39);
output(3, 153) <= input(41);
output(3, 154) <= input(43);
output(3, 155) <= input(45);
output(3, 156) <= input(46);
output(3, 157) <= input(49);
output(3, 158) <= input(50);
output(3, 159) <= input(54);
output(3, 160) <= input(12);
output(3, 161) <= input(13);
output(3, 162) <= input(14);
output(3, 163) <= input(15);
output(3, 164) <= input(32);
output(3, 165) <= input(34);
output(3, 166) <= input(36);
output(3, 167) <= input(37);
output(3, 168) <= input(40);
output(3, 169) <= input(42);
output(3, 170) <= input(44);
output(3, 171) <= input(47);
output(3, 172) <= input(48);
output(3, 173) <= input(51);
output(3, 174) <= input(52);
output(3, 175) <= input(53);
output(3, 176) <= input(13);
output(3, 177) <= input(14);
output(3, 178) <= input(15);
output(3, 179) <= input(32);
output(3, 180) <= input(34);
output(3, 181) <= input(36);
output(3, 182) <= input(37);
output(3, 183) <= input(40);
output(3, 184) <= input(42);
output(3, 185) <= input(44);
output(3, 186) <= input(47);
output(3, 187) <= input(48);
output(3, 188) <= input(51);
output(3, 189) <= input(52);
output(3, 190) <= input(53);
output(3, 191) <= input(57);
output(3, 192) <= input(14);
output(3, 193) <= input(15);
output(3, 194) <= input(32);
output(3, 195) <= input(34);
output(3, 196) <= input(36);
output(3, 197) <= input(37);
output(3, 198) <= input(40);
output(3, 199) <= input(42);
output(3, 200) <= input(44);
output(3, 201) <= input(47);
output(3, 202) <= input(48);
output(3, 203) <= input(51);
output(3, 204) <= input(52);
output(3, 205) <= input(53);
output(3, 206) <= input(57);
output(3, 207) <= input(58);
output(3, 208) <= input(30);
output(3, 209) <= input(31);
output(3, 210) <= input(33);
output(3, 211) <= input(35);
output(3, 212) <= input(38);
output(3, 213) <= input(39);
output(3, 214) <= input(41);
output(3, 215) <= input(43);
output(3, 216) <= input(45);
output(3, 217) <= input(46);
output(3, 218) <= input(49);
output(3, 219) <= input(50);
output(3, 220) <= input(54);
output(3, 221) <= input(55);
output(3, 222) <= input(56);
output(3, 223) <= input(59);
output(3, 224) <= input(31);
output(3, 225) <= input(33);
output(3, 226) <= input(35);
output(3, 227) <= input(38);
output(3, 228) <= input(39);
output(3, 229) <= input(41);
output(3, 230) <= input(43);
output(3, 231) <= input(45);
output(3, 232) <= input(46);
output(3, 233) <= input(49);
output(3, 234) <= input(50);
output(3, 235) <= input(54);
output(3, 236) <= input(55);
output(3, 237) <= input(56);
output(3, 238) <= input(59);
output(3, 239) <= input(60);
output(3, 240) <= input(33);
output(3, 241) <= input(35);
output(3, 242) <= input(38);
output(3, 243) <= input(39);
output(3, 244) <= input(41);
output(3, 245) <= input(43);
output(3, 246) <= input(45);
output(3, 247) <= input(46);
output(3, 248) <= input(49);
output(3, 249) <= input(50);
output(3, 250) <= input(54);
output(3, 251) <= input(55);
output(3, 252) <= input(56);
output(3, 253) <= input(59);
output(3, 254) <= input(60);
output(3, 255) <= input(61);
output(4, 0) <= input(21);
output(4, 1) <= input(22);
output(4, 2) <= input(23);
output(4, 3) <= input(24);
output(4, 4) <= input(25);
output(4, 5) <= input(26);
output(4, 6) <= input(27);
output(4, 7) <= input(28);
output(4, 8) <= input(29);
output(4, 9) <= input(30);
output(4, 10) <= input(31);
output(4, 11) <= input(33);
output(4, 12) <= input(35);
output(4, 13) <= input(38);
output(4, 14) <= input(39);
output(4, 15) <= input(41);
output(4, 16) <= input(22);
output(4, 17) <= input(23);
output(4, 18) <= input(24);
output(4, 19) <= input(25);
output(4, 20) <= input(26);
output(4, 21) <= input(27);
output(4, 22) <= input(28);
output(4, 23) <= input(29);
output(4, 24) <= input(30);
output(4, 25) <= input(31);
output(4, 26) <= input(33);
output(4, 27) <= input(35);
output(4, 28) <= input(38);
output(4, 29) <= input(39);
output(4, 30) <= input(41);
output(4, 31) <= input(43);
output(4, 32) <= input(23);
output(4, 33) <= input(24);
output(4, 34) <= input(25);
output(4, 35) <= input(26);
output(4, 36) <= input(27);
output(4, 37) <= input(28);
output(4, 38) <= input(29);
output(4, 39) <= input(30);
output(4, 40) <= input(31);
output(4, 41) <= input(33);
output(4, 42) <= input(35);
output(4, 43) <= input(38);
output(4, 44) <= input(39);
output(4, 45) <= input(41);
output(4, 46) <= input(43);
output(4, 47) <= input(45);
output(4, 48) <= input(24);
output(4, 49) <= input(25);
output(4, 50) <= input(26);
output(4, 51) <= input(27);
output(4, 52) <= input(28);
output(4, 53) <= input(29);
output(4, 54) <= input(30);
output(4, 55) <= input(31);
output(4, 56) <= input(33);
output(4, 57) <= input(35);
output(4, 58) <= input(38);
output(4, 59) <= input(39);
output(4, 60) <= input(41);
output(4, 61) <= input(43);
output(4, 62) <= input(45);
output(4, 63) <= input(46);
output(4, 64) <= input(25);
output(4, 65) <= input(26);
output(4, 66) <= input(27);
output(4, 67) <= input(28);
output(4, 68) <= input(29);
output(4, 69) <= input(30);
output(4, 70) <= input(31);
output(4, 71) <= input(33);
output(4, 72) <= input(35);
output(4, 73) <= input(38);
output(4, 74) <= input(39);
output(4, 75) <= input(41);
output(4, 76) <= input(43);
output(4, 77) <= input(45);
output(4, 78) <= input(46);
output(4, 79) <= input(49);
output(4, 80) <= input(10);
output(4, 81) <= input(11);
output(4, 82) <= input(12);
output(4, 83) <= input(13);
output(4, 84) <= input(14);
output(4, 85) <= input(15);
output(4, 86) <= input(32);
output(4, 87) <= input(34);
output(4, 88) <= input(36);
output(4, 89) <= input(37);
output(4, 90) <= input(40);
output(4, 91) <= input(42);
output(4, 92) <= input(44);
output(4, 93) <= input(47);
output(4, 94) <= input(48);
output(4, 95) <= input(51);
output(4, 96) <= input(11);
output(4, 97) <= input(12);
output(4, 98) <= input(13);
output(4, 99) <= input(14);
output(4, 100) <= input(15);
output(4, 101) <= input(32);
output(4, 102) <= input(34);
output(4, 103) <= input(36);
output(4, 104) <= input(37);
output(4, 105) <= input(40);
output(4, 106) <= input(42);
output(4, 107) <= input(44);
output(4, 108) <= input(47);
output(4, 109) <= input(48);
output(4, 110) <= input(51);
output(4, 111) <= input(52);
output(4, 112) <= input(12);
output(4, 113) <= input(13);
output(4, 114) <= input(14);
output(4, 115) <= input(15);
output(4, 116) <= input(32);
output(4, 117) <= input(34);
output(4, 118) <= input(36);
output(4, 119) <= input(37);
output(4, 120) <= input(40);
output(4, 121) <= input(42);
output(4, 122) <= input(44);
output(4, 123) <= input(47);
output(4, 124) <= input(48);
output(4, 125) <= input(51);
output(4, 126) <= input(52);
output(4, 127) <= input(53);
output(4, 128) <= input(13);
output(4, 129) <= input(14);
output(4, 130) <= input(15);
output(4, 131) <= input(32);
output(4, 132) <= input(34);
output(4, 133) <= input(36);
output(4, 134) <= input(37);
output(4, 135) <= input(40);
output(4, 136) <= input(42);
output(4, 137) <= input(44);
output(4, 138) <= input(47);
output(4, 139) <= input(48);
output(4, 140) <= input(51);
output(4, 141) <= input(52);
output(4, 142) <= input(53);
output(4, 143) <= input(57);
output(4, 144) <= input(14);
output(4, 145) <= input(15);
output(4, 146) <= input(32);
output(4, 147) <= input(34);
output(4, 148) <= input(36);
output(4, 149) <= input(37);
output(4, 150) <= input(40);
output(4, 151) <= input(42);
output(4, 152) <= input(44);
output(4, 153) <= input(47);
output(4, 154) <= input(48);
output(4, 155) <= input(51);
output(4, 156) <= input(52);
output(4, 157) <= input(53);
output(4, 158) <= input(57);
output(4, 159) <= input(58);
output(4, 160) <= input(30);
output(4, 161) <= input(31);
output(4, 162) <= input(33);
output(4, 163) <= input(35);
output(4, 164) <= input(38);
output(4, 165) <= input(39);
output(4, 166) <= input(41);
output(4, 167) <= input(43);
output(4, 168) <= input(45);
output(4, 169) <= input(46);
output(4, 170) <= input(49);
output(4, 171) <= input(50);
output(4, 172) <= input(54);
output(4, 173) <= input(55);
output(4, 174) <= input(56);
output(4, 175) <= input(59);
output(4, 176) <= input(31);
output(4, 177) <= input(33);
output(4, 178) <= input(35);
output(4, 179) <= input(38);
output(4, 180) <= input(39);
output(4, 181) <= input(41);
output(4, 182) <= input(43);
output(4, 183) <= input(45);
output(4, 184) <= input(46);
output(4, 185) <= input(49);
output(4, 186) <= input(50);
output(4, 187) <= input(54);
output(4, 188) <= input(55);
output(4, 189) <= input(56);
output(4, 190) <= input(59);
output(4, 191) <= input(60);
output(4, 192) <= input(33);
output(4, 193) <= input(35);
output(4, 194) <= input(38);
output(4, 195) <= input(39);
output(4, 196) <= input(41);
output(4, 197) <= input(43);
output(4, 198) <= input(45);
output(4, 199) <= input(46);
output(4, 200) <= input(49);
output(4, 201) <= input(50);
output(4, 202) <= input(54);
output(4, 203) <= input(55);
output(4, 204) <= input(56);
output(4, 205) <= input(59);
output(4, 206) <= input(60);
output(4, 207) <= input(61);
output(4, 208) <= input(35);
output(4, 209) <= input(38);
output(4, 210) <= input(39);
output(4, 211) <= input(41);
output(4, 212) <= input(43);
output(4, 213) <= input(45);
output(4, 214) <= input(46);
output(4, 215) <= input(49);
output(4, 216) <= input(50);
output(4, 217) <= input(54);
output(4, 218) <= input(55);
output(4, 219) <= input(56);
output(4, 220) <= input(59);
output(4, 221) <= input(60);
output(4, 222) <= input(61);
output(4, 223) <= input(62);
output(4, 224) <= input(38);
output(4, 225) <= input(39);
output(4, 226) <= input(41);
output(4, 227) <= input(43);
output(4, 228) <= input(45);
output(4, 229) <= input(46);
output(4, 230) <= input(49);
output(4, 231) <= input(50);
output(4, 232) <= input(54);
output(4, 233) <= input(55);
output(4, 234) <= input(56);
output(4, 235) <= input(59);
output(4, 236) <= input(60);
output(4, 237) <= input(61);
output(4, 238) <= input(62);
output(4, 239) <= input(63);
output(4, 240) <= input(39);
output(4, 241) <= input(41);
output(4, 242) <= input(43);
output(4, 243) <= input(45);
output(4, 244) <= input(46);
output(4, 245) <= input(49);
output(4, 246) <= input(50);
output(4, 247) <= input(54);
output(4, 248) <= input(55);
output(4, 249) <= input(56);
output(4, 250) <= input(59);
output(4, 251) <= input(60);
output(4, 252) <= input(61);
output(4, 253) <= input(62);
output(4, 254) <= input(63);
output(4, 255) <= input(64);
output(5, 0) <= input(23);
output(5, 1) <= input(24);
output(5, 2) <= input(25);
output(5, 3) <= input(26);
output(5, 4) <= input(27);
output(5, 5) <= input(28);
output(5, 6) <= input(29);
output(5, 7) <= input(30);
output(5, 8) <= input(31);
output(5, 9) <= input(33);
output(5, 10) <= input(35);
output(5, 11) <= input(38);
output(5, 12) <= input(39);
output(5, 13) <= input(41);
output(5, 14) <= input(43);
output(5, 15) <= input(45);
output(5, 16) <= input(24);
output(5, 17) <= input(25);
output(5, 18) <= input(26);
output(5, 19) <= input(27);
output(5, 20) <= input(28);
output(5, 21) <= input(29);
output(5, 22) <= input(30);
output(5, 23) <= input(31);
output(5, 24) <= input(33);
output(5, 25) <= input(35);
output(5, 26) <= input(38);
output(5, 27) <= input(39);
output(5, 28) <= input(41);
output(5, 29) <= input(43);
output(5, 30) <= input(45);
output(5, 31) <= input(46);
output(5, 32) <= input(25);
output(5, 33) <= input(26);
output(5, 34) <= input(27);
output(5, 35) <= input(28);
output(5, 36) <= input(29);
output(5, 37) <= input(30);
output(5, 38) <= input(31);
output(5, 39) <= input(33);
output(5, 40) <= input(35);
output(5, 41) <= input(38);
output(5, 42) <= input(39);
output(5, 43) <= input(41);
output(5, 44) <= input(43);
output(5, 45) <= input(45);
output(5, 46) <= input(46);
output(5, 47) <= input(49);
output(5, 48) <= input(26);
output(5, 49) <= input(27);
output(5, 50) <= input(28);
output(5, 51) <= input(29);
output(5, 52) <= input(30);
output(5, 53) <= input(31);
output(5, 54) <= input(33);
output(5, 55) <= input(35);
output(5, 56) <= input(38);
output(5, 57) <= input(39);
output(5, 58) <= input(41);
output(5, 59) <= input(43);
output(5, 60) <= input(45);
output(5, 61) <= input(46);
output(5, 62) <= input(49);
output(5, 63) <= input(50);
output(5, 64) <= input(27);
output(5, 65) <= input(28);
output(5, 66) <= input(29);
output(5, 67) <= input(30);
output(5, 68) <= input(31);
output(5, 69) <= input(33);
output(5, 70) <= input(35);
output(5, 71) <= input(38);
output(5, 72) <= input(39);
output(5, 73) <= input(41);
output(5, 74) <= input(43);
output(5, 75) <= input(45);
output(5, 76) <= input(46);
output(5, 77) <= input(49);
output(5, 78) <= input(50);
output(5, 79) <= input(54);
output(5, 80) <= input(28);
output(5, 81) <= input(29);
output(5, 82) <= input(30);
output(5, 83) <= input(31);
output(5, 84) <= input(33);
output(5, 85) <= input(35);
output(5, 86) <= input(38);
output(5, 87) <= input(39);
output(5, 88) <= input(41);
output(5, 89) <= input(43);
output(5, 90) <= input(45);
output(5, 91) <= input(46);
output(5, 92) <= input(49);
output(5, 93) <= input(50);
output(5, 94) <= input(54);
output(5, 95) <= input(55);
output(5, 96) <= input(29);
output(5, 97) <= input(30);
output(5, 98) <= input(31);
output(5, 99) <= input(33);
output(5, 100) <= input(35);
output(5, 101) <= input(38);
output(5, 102) <= input(39);
output(5, 103) <= input(41);
output(5, 104) <= input(43);
output(5, 105) <= input(45);
output(5, 106) <= input(46);
output(5, 107) <= input(49);
output(5, 108) <= input(50);
output(5, 109) <= input(54);
output(5, 110) <= input(55);
output(5, 111) <= input(56);
output(5, 112) <= input(30);
output(5, 113) <= input(31);
output(5, 114) <= input(33);
output(5, 115) <= input(35);
output(5, 116) <= input(38);
output(5, 117) <= input(39);
output(5, 118) <= input(41);
output(5, 119) <= input(43);
output(5, 120) <= input(45);
output(5, 121) <= input(46);
output(5, 122) <= input(49);
output(5, 123) <= input(50);
output(5, 124) <= input(54);
output(5, 125) <= input(55);
output(5, 126) <= input(56);
output(5, 127) <= input(59);
output(5, 128) <= input(31);
output(5, 129) <= input(33);
output(5, 130) <= input(35);
output(5, 131) <= input(38);
output(5, 132) <= input(39);
output(5, 133) <= input(41);
output(5, 134) <= input(43);
output(5, 135) <= input(45);
output(5, 136) <= input(46);
output(5, 137) <= input(49);
output(5, 138) <= input(50);
output(5, 139) <= input(54);
output(5, 140) <= input(55);
output(5, 141) <= input(56);
output(5, 142) <= input(59);
output(5, 143) <= input(60);
output(5, 144) <= input(33);
output(5, 145) <= input(35);
output(5, 146) <= input(38);
output(5, 147) <= input(39);
output(5, 148) <= input(41);
output(5, 149) <= input(43);
output(5, 150) <= input(45);
output(5, 151) <= input(46);
output(5, 152) <= input(49);
output(5, 153) <= input(50);
output(5, 154) <= input(54);
output(5, 155) <= input(55);
output(5, 156) <= input(56);
output(5, 157) <= input(59);
output(5, 158) <= input(60);
output(5, 159) <= input(61);
output(5, 160) <= input(35);
output(5, 161) <= input(38);
output(5, 162) <= input(39);
output(5, 163) <= input(41);
output(5, 164) <= input(43);
output(5, 165) <= input(45);
output(5, 166) <= input(46);
output(5, 167) <= input(49);
output(5, 168) <= input(50);
output(5, 169) <= input(54);
output(5, 170) <= input(55);
output(5, 171) <= input(56);
output(5, 172) <= input(59);
output(5, 173) <= input(60);
output(5, 174) <= input(61);
output(5, 175) <= input(62);
output(5, 176) <= input(38);
output(5, 177) <= input(39);
output(5, 178) <= input(41);
output(5, 179) <= input(43);
output(5, 180) <= input(45);
output(5, 181) <= input(46);
output(5, 182) <= input(49);
output(5, 183) <= input(50);
output(5, 184) <= input(54);
output(5, 185) <= input(55);
output(5, 186) <= input(56);
output(5, 187) <= input(59);
output(5, 188) <= input(60);
output(5, 189) <= input(61);
output(5, 190) <= input(62);
output(5, 191) <= input(63);
output(5, 192) <= input(39);
output(5, 193) <= input(41);
output(5, 194) <= input(43);
output(5, 195) <= input(45);
output(5, 196) <= input(46);
output(5, 197) <= input(49);
output(5, 198) <= input(50);
output(5, 199) <= input(54);
output(5, 200) <= input(55);
output(5, 201) <= input(56);
output(5, 202) <= input(59);
output(5, 203) <= input(60);
output(5, 204) <= input(61);
output(5, 205) <= input(62);
output(5, 206) <= input(63);
output(5, 207) <= input(64);
output(5, 208) <= input(41);
output(5, 209) <= input(43);
output(5, 210) <= input(45);
output(5, 211) <= input(46);
output(5, 212) <= input(49);
output(5, 213) <= input(50);
output(5, 214) <= input(54);
output(5, 215) <= input(55);
output(5, 216) <= input(56);
output(5, 217) <= input(59);
output(5, 218) <= input(60);
output(5, 219) <= input(61);
output(5, 220) <= input(62);
output(5, 221) <= input(63);
output(5, 222) <= input(64);
output(5, 223) <= input(65);
output(5, 224) <= input(43);
output(5, 225) <= input(45);
output(5, 226) <= input(46);
output(5, 227) <= input(49);
output(5, 228) <= input(50);
output(5, 229) <= input(54);
output(5, 230) <= input(55);
output(5, 231) <= input(56);
output(5, 232) <= input(59);
output(5, 233) <= input(60);
output(5, 234) <= input(61);
output(5, 235) <= input(62);
output(5, 236) <= input(63);
output(5, 237) <= input(64);
output(5, 238) <= input(65);
output(5, 239) <= input(66);
output(5, 240) <= input(45);
output(5, 241) <= input(46);
output(5, 242) <= input(49);
output(5, 243) <= input(50);
output(5, 244) <= input(54);
output(5, 245) <= input(55);
output(5, 246) <= input(56);
output(5, 247) <= input(59);
output(5, 248) <= input(60);
output(5, 249) <= input(61);
output(5, 250) <= input(62);
output(5, 251) <= input(63);
output(5, 252) <= input(64);
output(5, 253) <= input(65);
output(5, 254) <= input(66);
output(5, 255) <= input(67);
when others => for i in 0 to 7 loop for j in 0 to 255 loop output(i,j) <= "00000000"; end loop; end loop;
end case;
elsif control = "111" then 
case iteration_control is
when "0000" =>
output(0, 0) <= input(0);
output(0, 1) <= input(1);
output(0, 2) <= input(2);
output(0, 3) <= input(3);
output(0, 4) <= input(4);
output(0, 5) <= input(5);
output(0, 6) <= input(6);
output(0, 7) <= input(7);
output(0, 8) <= input(8);
output(0, 9) <= input(9);
output(0, 10) <= input(10);
output(0, 11) <= input(11);
output(0, 12) <= input(12);
output(0, 13) <= input(13);
output(0, 14) <= input(14);
output(0, 15) <= input(15);
output(0, 16) <= input(1);
output(0, 17) <= input(2);
output(0, 18) <= input(3);
output(0, 19) <= input(4);
output(0, 20) <= input(5);
output(0, 21) <= input(6);
output(0, 22) <= input(7);
output(0, 23) <= input(8);
output(0, 24) <= input(9);
output(0, 25) <= input(10);
output(0, 26) <= input(11);
output(0, 27) <= input(12);
output(0, 28) <= input(13);
output(0, 29) <= input(14);
output(0, 30) <= input(15);
output(0, 31) <= input(16);
output(0, 32) <= input(2);
output(0, 33) <= input(3);
output(0, 34) <= input(4);
output(0, 35) <= input(5);
output(0, 36) <= input(6);
output(0, 37) <= input(7);
output(0, 38) <= input(8);
output(0, 39) <= input(9);
output(0, 40) <= input(10);
output(0, 41) <= input(11);
output(0, 42) <= input(12);
output(0, 43) <= input(13);
output(0, 44) <= input(14);
output(0, 45) <= input(15);
output(0, 46) <= input(16);
output(0, 47) <= input(17);
output(0, 48) <= input(3);
output(0, 49) <= input(4);
output(0, 50) <= input(5);
output(0, 51) <= input(6);
output(0, 52) <= input(7);
output(0, 53) <= input(8);
output(0, 54) <= input(9);
output(0, 55) <= input(10);
output(0, 56) <= input(11);
output(0, 57) <= input(12);
output(0, 58) <= input(13);
output(0, 59) <= input(14);
output(0, 60) <= input(15);
output(0, 61) <= input(16);
output(0, 62) <= input(17);
output(0, 63) <= input(18);
output(0, 64) <= input(4);
output(0, 65) <= input(5);
output(0, 66) <= input(6);
output(0, 67) <= input(7);
output(0, 68) <= input(8);
output(0, 69) <= input(9);
output(0, 70) <= input(10);
output(0, 71) <= input(11);
output(0, 72) <= input(12);
output(0, 73) <= input(13);
output(0, 74) <= input(14);
output(0, 75) <= input(15);
output(0, 76) <= input(16);
output(0, 77) <= input(17);
output(0, 78) <= input(18);
output(0, 79) <= input(19);
output(0, 80) <= input(5);
output(0, 81) <= input(6);
output(0, 82) <= input(7);
output(0, 83) <= input(8);
output(0, 84) <= input(9);
output(0, 85) <= input(10);
output(0, 86) <= input(11);
output(0, 87) <= input(12);
output(0, 88) <= input(13);
output(0, 89) <= input(14);
output(0, 90) <= input(15);
output(0, 91) <= input(16);
output(0, 92) <= input(17);
output(0, 93) <= input(18);
output(0, 94) <= input(19);
output(0, 95) <= input(20);
output(0, 96) <= input(6);
output(0, 97) <= input(7);
output(0, 98) <= input(8);
output(0, 99) <= input(9);
output(0, 100) <= input(10);
output(0, 101) <= input(11);
output(0, 102) <= input(12);
output(0, 103) <= input(13);
output(0, 104) <= input(14);
output(0, 105) <= input(15);
output(0, 106) <= input(16);
output(0, 107) <= input(17);
output(0, 108) <= input(18);
output(0, 109) <= input(19);
output(0, 110) <= input(20);
output(0, 111) <= input(21);
output(0, 112) <= input(7);
output(0, 113) <= input(8);
output(0, 114) <= input(9);
output(0, 115) <= input(10);
output(0, 116) <= input(11);
output(0, 117) <= input(12);
output(0, 118) <= input(13);
output(0, 119) <= input(14);
output(0, 120) <= input(15);
output(0, 121) <= input(16);
output(0, 122) <= input(17);
output(0, 123) <= input(18);
output(0, 124) <= input(19);
output(0, 125) <= input(20);
output(0, 126) <= input(21);
output(0, 127) <= input(22);
output(0, 128) <= input(8);
output(0, 129) <= input(9);
output(0, 130) <= input(10);
output(0, 131) <= input(11);
output(0, 132) <= input(12);
output(0, 133) <= input(13);
output(0, 134) <= input(14);
output(0, 135) <= input(15);
output(0, 136) <= input(16);
output(0, 137) <= input(17);
output(0, 138) <= input(18);
output(0, 139) <= input(19);
output(0, 140) <= input(20);
output(0, 141) <= input(21);
output(0, 142) <= input(22);
output(0, 143) <= input(23);
output(0, 144) <= input(9);
output(0, 145) <= input(10);
output(0, 146) <= input(11);
output(0, 147) <= input(12);
output(0, 148) <= input(13);
output(0, 149) <= input(14);
output(0, 150) <= input(15);
output(0, 151) <= input(16);
output(0, 152) <= input(17);
output(0, 153) <= input(18);
output(0, 154) <= input(19);
output(0, 155) <= input(20);
output(0, 156) <= input(21);
output(0, 157) <= input(22);
output(0, 158) <= input(23);
output(0, 159) <= input(24);
output(0, 160) <= input(10);
output(0, 161) <= input(11);
output(0, 162) <= input(12);
output(0, 163) <= input(13);
output(0, 164) <= input(14);
output(0, 165) <= input(15);
output(0, 166) <= input(16);
output(0, 167) <= input(17);
output(0, 168) <= input(18);
output(0, 169) <= input(19);
output(0, 170) <= input(20);
output(0, 171) <= input(21);
output(0, 172) <= input(22);
output(0, 173) <= input(23);
output(0, 174) <= input(24);
output(0, 175) <= input(25);
output(0, 176) <= input(11);
output(0, 177) <= input(12);
output(0, 178) <= input(13);
output(0, 179) <= input(14);
output(0, 180) <= input(15);
output(0, 181) <= input(16);
output(0, 182) <= input(17);
output(0, 183) <= input(18);
output(0, 184) <= input(19);
output(0, 185) <= input(20);
output(0, 186) <= input(21);
output(0, 187) <= input(22);
output(0, 188) <= input(23);
output(0, 189) <= input(24);
output(0, 190) <= input(25);
output(0, 191) <= input(26);
output(0, 192) <= input(12);
output(0, 193) <= input(13);
output(0, 194) <= input(14);
output(0, 195) <= input(15);
output(0, 196) <= input(16);
output(0, 197) <= input(17);
output(0, 198) <= input(18);
output(0, 199) <= input(19);
output(0, 200) <= input(20);
output(0, 201) <= input(21);
output(0, 202) <= input(22);
output(0, 203) <= input(23);
output(0, 204) <= input(24);
output(0, 205) <= input(25);
output(0, 206) <= input(26);
output(0, 207) <= input(27);
output(0, 208) <= input(13);
output(0, 209) <= input(14);
output(0, 210) <= input(15);
output(0, 211) <= input(16);
output(0, 212) <= input(17);
output(0, 213) <= input(18);
output(0, 214) <= input(19);
output(0, 215) <= input(20);
output(0, 216) <= input(21);
output(0, 217) <= input(22);
output(0, 218) <= input(23);
output(0, 219) <= input(24);
output(0, 220) <= input(25);
output(0, 221) <= input(26);
output(0, 222) <= input(27);
output(0, 223) <= input(28);
output(0, 224) <= input(14);
output(0, 225) <= input(15);
output(0, 226) <= input(16);
output(0, 227) <= input(17);
output(0, 228) <= input(18);
output(0, 229) <= input(19);
output(0, 230) <= input(20);
output(0, 231) <= input(21);
output(0, 232) <= input(22);
output(0, 233) <= input(23);
output(0, 234) <= input(24);
output(0, 235) <= input(25);
output(0, 236) <= input(26);
output(0, 237) <= input(27);
output(0, 238) <= input(28);
output(0, 239) <= input(29);
output(0, 240) <= input(15);
output(0, 241) <= input(16);
output(0, 242) <= input(17);
output(0, 243) <= input(18);
output(0, 244) <= input(19);
output(0, 245) <= input(20);
output(0, 246) <= input(21);
output(0, 247) <= input(22);
output(0, 248) <= input(23);
output(0, 249) <= input(24);
output(0, 250) <= input(25);
output(0, 251) <= input(26);
output(0, 252) <= input(27);
output(0, 253) <= input(28);
output(0, 254) <= input(29);
output(0, 255) <= input(30);
output(1, 0) <= input(31);
output(1, 1) <= input(32);
output(1, 2) <= input(0);
output(1, 3) <= input(1);
output(1, 4) <= input(2);
output(1, 5) <= input(3);
output(1, 6) <= input(4);
output(1, 7) <= input(5);
output(1, 8) <= input(6);
output(1, 9) <= input(7);
output(1, 10) <= input(8);
output(1, 11) <= input(9);
output(1, 12) <= input(10);
output(1, 13) <= input(11);
output(1, 14) <= input(12);
output(1, 15) <= input(13);
output(1, 16) <= input(32);
output(1, 17) <= input(0);
output(1, 18) <= input(1);
output(1, 19) <= input(2);
output(1, 20) <= input(3);
output(1, 21) <= input(4);
output(1, 22) <= input(5);
output(1, 23) <= input(6);
output(1, 24) <= input(7);
output(1, 25) <= input(8);
output(1, 26) <= input(9);
output(1, 27) <= input(10);
output(1, 28) <= input(11);
output(1, 29) <= input(12);
output(1, 30) <= input(13);
output(1, 31) <= input(14);
output(1, 32) <= input(0);
output(1, 33) <= input(1);
output(1, 34) <= input(2);
output(1, 35) <= input(3);
output(1, 36) <= input(4);
output(1, 37) <= input(5);
output(1, 38) <= input(6);
output(1, 39) <= input(7);
output(1, 40) <= input(8);
output(1, 41) <= input(9);
output(1, 42) <= input(10);
output(1, 43) <= input(11);
output(1, 44) <= input(12);
output(1, 45) <= input(13);
output(1, 46) <= input(14);
output(1, 47) <= input(15);
output(1, 48) <= input(1);
output(1, 49) <= input(2);
output(1, 50) <= input(3);
output(1, 51) <= input(4);
output(1, 52) <= input(5);
output(1, 53) <= input(6);
output(1, 54) <= input(7);
output(1, 55) <= input(8);
output(1, 56) <= input(9);
output(1, 57) <= input(10);
output(1, 58) <= input(11);
output(1, 59) <= input(12);
output(1, 60) <= input(13);
output(1, 61) <= input(14);
output(1, 62) <= input(15);
output(1, 63) <= input(16);
output(1, 64) <= input(2);
output(1, 65) <= input(3);
output(1, 66) <= input(4);
output(1, 67) <= input(5);
output(1, 68) <= input(6);
output(1, 69) <= input(7);
output(1, 70) <= input(8);
output(1, 71) <= input(9);
output(1, 72) <= input(10);
output(1, 73) <= input(11);
output(1, 74) <= input(12);
output(1, 75) <= input(13);
output(1, 76) <= input(14);
output(1, 77) <= input(15);
output(1, 78) <= input(16);
output(1, 79) <= input(17);
output(1, 80) <= input(33);
output(1, 81) <= input(34);
output(1, 82) <= input(35);
output(1, 83) <= input(36);
output(1, 84) <= input(37);
output(1, 85) <= input(38);
output(1, 86) <= input(39);
output(1, 87) <= input(40);
output(1, 88) <= input(41);
output(1, 89) <= input(42);
output(1, 90) <= input(43);
output(1, 91) <= input(44);
output(1, 92) <= input(45);
output(1, 93) <= input(46);
output(1, 94) <= input(47);
output(1, 95) <= input(48);
output(1, 96) <= input(34);
output(1, 97) <= input(35);
output(1, 98) <= input(36);
output(1, 99) <= input(37);
output(1, 100) <= input(38);
output(1, 101) <= input(39);
output(1, 102) <= input(40);
output(1, 103) <= input(41);
output(1, 104) <= input(42);
output(1, 105) <= input(43);
output(1, 106) <= input(44);
output(1, 107) <= input(45);
output(1, 108) <= input(46);
output(1, 109) <= input(47);
output(1, 110) <= input(48);
output(1, 111) <= input(49);
output(1, 112) <= input(35);
output(1, 113) <= input(36);
output(1, 114) <= input(37);
output(1, 115) <= input(38);
output(1, 116) <= input(39);
output(1, 117) <= input(40);
output(1, 118) <= input(41);
output(1, 119) <= input(42);
output(1, 120) <= input(43);
output(1, 121) <= input(44);
output(1, 122) <= input(45);
output(1, 123) <= input(46);
output(1, 124) <= input(47);
output(1, 125) <= input(48);
output(1, 126) <= input(49);
output(1, 127) <= input(50);
output(1, 128) <= input(36);
output(1, 129) <= input(37);
output(1, 130) <= input(38);
output(1, 131) <= input(39);
output(1, 132) <= input(40);
output(1, 133) <= input(41);
output(1, 134) <= input(42);
output(1, 135) <= input(43);
output(1, 136) <= input(44);
output(1, 137) <= input(45);
output(1, 138) <= input(46);
output(1, 139) <= input(47);
output(1, 140) <= input(48);
output(1, 141) <= input(49);
output(1, 142) <= input(50);
output(1, 143) <= input(51);
output(1, 144) <= input(37);
output(1, 145) <= input(38);
output(1, 146) <= input(39);
output(1, 147) <= input(40);
output(1, 148) <= input(41);
output(1, 149) <= input(42);
output(1, 150) <= input(43);
output(1, 151) <= input(44);
output(1, 152) <= input(45);
output(1, 153) <= input(46);
output(1, 154) <= input(47);
output(1, 155) <= input(48);
output(1, 156) <= input(49);
output(1, 157) <= input(50);
output(1, 158) <= input(51);
output(1, 159) <= input(52);
output(1, 160) <= input(7);
output(1, 161) <= input(8);
output(1, 162) <= input(9);
output(1, 163) <= input(10);
output(1, 164) <= input(11);
output(1, 165) <= input(12);
output(1, 166) <= input(13);
output(1, 167) <= input(14);
output(1, 168) <= input(15);
output(1, 169) <= input(16);
output(1, 170) <= input(17);
output(1, 171) <= input(18);
output(1, 172) <= input(19);
output(1, 173) <= input(20);
output(1, 174) <= input(21);
output(1, 175) <= input(22);
output(1, 176) <= input(8);
output(1, 177) <= input(9);
output(1, 178) <= input(10);
output(1, 179) <= input(11);
output(1, 180) <= input(12);
output(1, 181) <= input(13);
output(1, 182) <= input(14);
output(1, 183) <= input(15);
output(1, 184) <= input(16);
output(1, 185) <= input(17);
output(1, 186) <= input(18);
output(1, 187) <= input(19);
output(1, 188) <= input(20);
output(1, 189) <= input(21);
output(1, 190) <= input(22);
output(1, 191) <= input(23);
output(1, 192) <= input(9);
output(1, 193) <= input(10);
output(1, 194) <= input(11);
output(1, 195) <= input(12);
output(1, 196) <= input(13);
output(1, 197) <= input(14);
output(1, 198) <= input(15);
output(1, 199) <= input(16);
output(1, 200) <= input(17);
output(1, 201) <= input(18);
output(1, 202) <= input(19);
output(1, 203) <= input(20);
output(1, 204) <= input(21);
output(1, 205) <= input(22);
output(1, 206) <= input(23);
output(1, 207) <= input(24);
output(1, 208) <= input(10);
output(1, 209) <= input(11);
output(1, 210) <= input(12);
output(1, 211) <= input(13);
output(1, 212) <= input(14);
output(1, 213) <= input(15);
output(1, 214) <= input(16);
output(1, 215) <= input(17);
output(1, 216) <= input(18);
output(1, 217) <= input(19);
output(1, 218) <= input(20);
output(1, 219) <= input(21);
output(1, 220) <= input(22);
output(1, 221) <= input(23);
output(1, 222) <= input(24);
output(1, 223) <= input(25);
output(1, 224) <= input(11);
output(1, 225) <= input(12);
output(1, 226) <= input(13);
output(1, 227) <= input(14);
output(1, 228) <= input(15);
output(1, 229) <= input(16);
output(1, 230) <= input(17);
output(1, 231) <= input(18);
output(1, 232) <= input(19);
output(1, 233) <= input(20);
output(1, 234) <= input(21);
output(1, 235) <= input(22);
output(1, 236) <= input(23);
output(1, 237) <= input(24);
output(1, 238) <= input(25);
output(1, 239) <= input(26);
output(1, 240) <= input(12);
output(1, 241) <= input(13);
output(1, 242) <= input(14);
output(1, 243) <= input(15);
output(1, 244) <= input(16);
output(1, 245) <= input(17);
output(1, 246) <= input(18);
output(1, 247) <= input(19);
output(1, 248) <= input(20);
output(1, 249) <= input(21);
output(1, 250) <= input(22);
output(1, 251) <= input(23);
output(1, 252) <= input(24);
output(1, 253) <= input(25);
output(1, 254) <= input(26);
output(1, 255) <= input(27);
output(2, 0) <= input(53);
output(2, 1) <= input(54);
output(2, 2) <= input(55);
output(2, 3) <= input(56);
output(2, 4) <= input(57);
output(2, 5) <= input(58);
output(2, 6) <= input(33);
output(2, 7) <= input(34);
output(2, 8) <= input(35);
output(2, 9) <= input(36);
output(2, 10) <= input(37);
output(2, 11) <= input(38);
output(2, 12) <= input(39);
output(2, 13) <= input(40);
output(2, 14) <= input(41);
output(2, 15) <= input(42);
output(2, 16) <= input(54);
output(2, 17) <= input(55);
output(2, 18) <= input(56);
output(2, 19) <= input(57);
output(2, 20) <= input(58);
output(2, 21) <= input(33);
output(2, 22) <= input(34);
output(2, 23) <= input(35);
output(2, 24) <= input(36);
output(2, 25) <= input(37);
output(2, 26) <= input(38);
output(2, 27) <= input(39);
output(2, 28) <= input(40);
output(2, 29) <= input(41);
output(2, 30) <= input(42);
output(2, 31) <= input(43);
output(2, 32) <= input(31);
output(2, 33) <= input(32);
output(2, 34) <= input(0);
output(2, 35) <= input(1);
output(2, 36) <= input(2);
output(2, 37) <= input(3);
output(2, 38) <= input(4);
output(2, 39) <= input(5);
output(2, 40) <= input(6);
output(2, 41) <= input(7);
output(2, 42) <= input(8);
output(2, 43) <= input(9);
output(2, 44) <= input(10);
output(2, 45) <= input(11);
output(2, 46) <= input(12);
output(2, 47) <= input(13);
output(2, 48) <= input(32);
output(2, 49) <= input(0);
output(2, 50) <= input(1);
output(2, 51) <= input(2);
output(2, 52) <= input(3);
output(2, 53) <= input(4);
output(2, 54) <= input(5);
output(2, 55) <= input(6);
output(2, 56) <= input(7);
output(2, 57) <= input(8);
output(2, 58) <= input(9);
output(2, 59) <= input(10);
output(2, 60) <= input(11);
output(2, 61) <= input(12);
output(2, 62) <= input(13);
output(2, 63) <= input(14);
output(2, 64) <= input(0);
output(2, 65) <= input(1);
output(2, 66) <= input(2);
output(2, 67) <= input(3);
output(2, 68) <= input(4);
output(2, 69) <= input(5);
output(2, 70) <= input(6);
output(2, 71) <= input(7);
output(2, 72) <= input(8);
output(2, 73) <= input(9);
output(2, 74) <= input(10);
output(2, 75) <= input(11);
output(2, 76) <= input(12);
output(2, 77) <= input(13);
output(2, 78) <= input(14);
output(2, 79) <= input(15);
output(2, 80) <= input(57);
output(2, 81) <= input(58);
output(2, 82) <= input(33);
output(2, 83) <= input(34);
output(2, 84) <= input(35);
output(2, 85) <= input(36);
output(2, 86) <= input(37);
output(2, 87) <= input(38);
output(2, 88) <= input(39);
output(2, 89) <= input(40);
output(2, 90) <= input(41);
output(2, 91) <= input(42);
output(2, 92) <= input(43);
output(2, 93) <= input(44);
output(2, 94) <= input(45);
output(2, 95) <= input(46);
output(2, 96) <= input(58);
output(2, 97) <= input(33);
output(2, 98) <= input(34);
output(2, 99) <= input(35);
output(2, 100) <= input(36);
output(2, 101) <= input(37);
output(2, 102) <= input(38);
output(2, 103) <= input(39);
output(2, 104) <= input(40);
output(2, 105) <= input(41);
output(2, 106) <= input(42);
output(2, 107) <= input(43);
output(2, 108) <= input(44);
output(2, 109) <= input(45);
output(2, 110) <= input(46);
output(2, 111) <= input(47);
output(2, 112) <= input(33);
output(2, 113) <= input(34);
output(2, 114) <= input(35);
output(2, 115) <= input(36);
output(2, 116) <= input(37);
output(2, 117) <= input(38);
output(2, 118) <= input(39);
output(2, 119) <= input(40);
output(2, 120) <= input(41);
output(2, 121) <= input(42);
output(2, 122) <= input(43);
output(2, 123) <= input(44);
output(2, 124) <= input(45);
output(2, 125) <= input(46);
output(2, 126) <= input(47);
output(2, 127) <= input(48);
output(2, 128) <= input(3);
output(2, 129) <= input(4);
output(2, 130) <= input(5);
output(2, 131) <= input(6);
output(2, 132) <= input(7);
output(2, 133) <= input(8);
output(2, 134) <= input(9);
output(2, 135) <= input(10);
output(2, 136) <= input(11);
output(2, 137) <= input(12);
output(2, 138) <= input(13);
output(2, 139) <= input(14);
output(2, 140) <= input(15);
output(2, 141) <= input(16);
output(2, 142) <= input(17);
output(2, 143) <= input(18);
output(2, 144) <= input(4);
output(2, 145) <= input(5);
output(2, 146) <= input(6);
output(2, 147) <= input(7);
output(2, 148) <= input(8);
output(2, 149) <= input(9);
output(2, 150) <= input(10);
output(2, 151) <= input(11);
output(2, 152) <= input(12);
output(2, 153) <= input(13);
output(2, 154) <= input(14);
output(2, 155) <= input(15);
output(2, 156) <= input(16);
output(2, 157) <= input(17);
output(2, 158) <= input(18);
output(2, 159) <= input(19);
output(2, 160) <= input(35);
output(2, 161) <= input(36);
output(2, 162) <= input(37);
output(2, 163) <= input(38);
output(2, 164) <= input(39);
output(2, 165) <= input(40);
output(2, 166) <= input(41);
output(2, 167) <= input(42);
output(2, 168) <= input(43);
output(2, 169) <= input(44);
output(2, 170) <= input(45);
output(2, 171) <= input(46);
output(2, 172) <= input(47);
output(2, 173) <= input(48);
output(2, 174) <= input(49);
output(2, 175) <= input(50);
output(2, 176) <= input(36);
output(2, 177) <= input(37);
output(2, 178) <= input(38);
output(2, 179) <= input(39);
output(2, 180) <= input(40);
output(2, 181) <= input(41);
output(2, 182) <= input(42);
output(2, 183) <= input(43);
output(2, 184) <= input(44);
output(2, 185) <= input(45);
output(2, 186) <= input(46);
output(2, 187) <= input(47);
output(2, 188) <= input(48);
output(2, 189) <= input(49);
output(2, 190) <= input(50);
output(2, 191) <= input(51);
output(2, 192) <= input(37);
output(2, 193) <= input(38);
output(2, 194) <= input(39);
output(2, 195) <= input(40);
output(2, 196) <= input(41);
output(2, 197) <= input(42);
output(2, 198) <= input(43);
output(2, 199) <= input(44);
output(2, 200) <= input(45);
output(2, 201) <= input(46);
output(2, 202) <= input(47);
output(2, 203) <= input(48);
output(2, 204) <= input(49);
output(2, 205) <= input(50);
output(2, 206) <= input(51);
output(2, 207) <= input(52);
output(2, 208) <= input(7);
output(2, 209) <= input(8);
output(2, 210) <= input(9);
output(2, 211) <= input(10);
output(2, 212) <= input(11);
output(2, 213) <= input(12);
output(2, 214) <= input(13);
output(2, 215) <= input(14);
output(2, 216) <= input(15);
output(2, 217) <= input(16);
output(2, 218) <= input(17);
output(2, 219) <= input(18);
output(2, 220) <= input(19);
output(2, 221) <= input(20);
output(2, 222) <= input(21);
output(2, 223) <= input(22);
output(2, 224) <= input(8);
output(2, 225) <= input(9);
output(2, 226) <= input(10);
output(2, 227) <= input(11);
output(2, 228) <= input(12);
output(2, 229) <= input(13);
output(2, 230) <= input(14);
output(2, 231) <= input(15);
output(2, 232) <= input(16);
output(2, 233) <= input(17);
output(2, 234) <= input(18);
output(2, 235) <= input(19);
output(2, 236) <= input(20);
output(2, 237) <= input(21);
output(2, 238) <= input(22);
output(2, 239) <= input(23);
output(2, 240) <= input(9);
output(2, 241) <= input(10);
output(2, 242) <= input(11);
output(2, 243) <= input(12);
output(2, 244) <= input(13);
output(2, 245) <= input(14);
output(2, 246) <= input(15);
output(2, 247) <= input(16);
output(2, 248) <= input(17);
output(2, 249) <= input(18);
output(2, 250) <= input(19);
output(2, 251) <= input(20);
output(2, 252) <= input(21);
output(2, 253) <= input(22);
output(2, 254) <= input(23);
output(2, 255) <= input(24);
output(3, 0) <= input(59);
output(3, 1) <= input(60);
output(3, 2) <= input(61);
output(3, 3) <= input(31);
output(3, 4) <= input(32);
output(3, 5) <= input(0);
output(3, 6) <= input(1);
output(3, 7) <= input(2);
output(3, 8) <= input(3);
output(3, 9) <= input(4);
output(3, 10) <= input(5);
output(3, 11) <= input(6);
output(3, 12) <= input(7);
output(3, 13) <= input(8);
output(3, 14) <= input(9);
output(3, 15) <= input(10);
output(3, 16) <= input(62);
output(3, 17) <= input(53);
output(3, 18) <= input(54);
output(3, 19) <= input(55);
output(3, 20) <= input(56);
output(3, 21) <= input(57);
output(3, 22) <= input(58);
output(3, 23) <= input(33);
output(3, 24) <= input(34);
output(3, 25) <= input(35);
output(3, 26) <= input(36);
output(3, 27) <= input(37);
output(3, 28) <= input(38);
output(3, 29) <= input(39);
output(3, 30) <= input(40);
output(3, 31) <= input(41);
output(3, 32) <= input(53);
output(3, 33) <= input(54);
output(3, 34) <= input(55);
output(3, 35) <= input(56);
output(3, 36) <= input(57);
output(3, 37) <= input(58);
output(3, 38) <= input(33);
output(3, 39) <= input(34);
output(3, 40) <= input(35);
output(3, 41) <= input(36);
output(3, 42) <= input(37);
output(3, 43) <= input(38);
output(3, 44) <= input(39);
output(3, 45) <= input(40);
output(3, 46) <= input(41);
output(3, 47) <= input(42);
output(3, 48) <= input(61);
output(3, 49) <= input(31);
output(3, 50) <= input(32);
output(3, 51) <= input(0);
output(3, 52) <= input(1);
output(3, 53) <= input(2);
output(3, 54) <= input(3);
output(3, 55) <= input(4);
output(3, 56) <= input(5);
output(3, 57) <= input(6);
output(3, 58) <= input(7);
output(3, 59) <= input(8);
output(3, 60) <= input(9);
output(3, 61) <= input(10);
output(3, 62) <= input(11);
output(3, 63) <= input(12);
output(3, 64) <= input(31);
output(3, 65) <= input(32);
output(3, 66) <= input(0);
output(3, 67) <= input(1);
output(3, 68) <= input(2);
output(3, 69) <= input(3);
output(3, 70) <= input(4);
output(3, 71) <= input(5);
output(3, 72) <= input(6);
output(3, 73) <= input(7);
output(3, 74) <= input(8);
output(3, 75) <= input(9);
output(3, 76) <= input(10);
output(3, 77) <= input(11);
output(3, 78) <= input(12);
output(3, 79) <= input(13);
output(3, 80) <= input(55);
output(3, 81) <= input(56);
output(3, 82) <= input(57);
output(3, 83) <= input(58);
output(3, 84) <= input(33);
output(3, 85) <= input(34);
output(3, 86) <= input(35);
output(3, 87) <= input(36);
output(3, 88) <= input(37);
output(3, 89) <= input(38);
output(3, 90) <= input(39);
output(3, 91) <= input(40);
output(3, 92) <= input(41);
output(3, 93) <= input(42);
output(3, 94) <= input(43);
output(3, 95) <= input(44);
output(3, 96) <= input(56);
output(3, 97) <= input(57);
output(3, 98) <= input(58);
output(3, 99) <= input(33);
output(3, 100) <= input(34);
output(3, 101) <= input(35);
output(3, 102) <= input(36);
output(3, 103) <= input(37);
output(3, 104) <= input(38);
output(3, 105) <= input(39);
output(3, 106) <= input(40);
output(3, 107) <= input(41);
output(3, 108) <= input(42);
output(3, 109) <= input(43);
output(3, 110) <= input(44);
output(3, 111) <= input(45);
output(3, 112) <= input(0);
output(3, 113) <= input(1);
output(3, 114) <= input(2);
output(3, 115) <= input(3);
output(3, 116) <= input(4);
output(3, 117) <= input(5);
output(3, 118) <= input(6);
output(3, 119) <= input(7);
output(3, 120) <= input(8);
output(3, 121) <= input(9);
output(3, 122) <= input(10);
output(3, 123) <= input(11);
output(3, 124) <= input(12);
output(3, 125) <= input(13);
output(3, 126) <= input(14);
output(3, 127) <= input(15);
output(3, 128) <= input(57);
output(3, 129) <= input(58);
output(3, 130) <= input(33);
output(3, 131) <= input(34);
output(3, 132) <= input(35);
output(3, 133) <= input(36);
output(3, 134) <= input(37);
output(3, 135) <= input(38);
output(3, 136) <= input(39);
output(3, 137) <= input(40);
output(3, 138) <= input(41);
output(3, 139) <= input(42);
output(3, 140) <= input(43);
output(3, 141) <= input(44);
output(3, 142) <= input(45);
output(3, 143) <= input(46);
output(3, 144) <= input(58);
output(3, 145) <= input(33);
output(3, 146) <= input(34);
output(3, 147) <= input(35);
output(3, 148) <= input(36);
output(3, 149) <= input(37);
output(3, 150) <= input(38);
output(3, 151) <= input(39);
output(3, 152) <= input(40);
output(3, 153) <= input(41);
output(3, 154) <= input(42);
output(3, 155) <= input(43);
output(3, 156) <= input(44);
output(3, 157) <= input(45);
output(3, 158) <= input(46);
output(3, 159) <= input(47);
output(3, 160) <= input(2);
output(3, 161) <= input(3);
output(3, 162) <= input(4);
output(3, 163) <= input(5);
output(3, 164) <= input(6);
output(3, 165) <= input(7);
output(3, 166) <= input(8);
output(3, 167) <= input(9);
output(3, 168) <= input(10);
output(3, 169) <= input(11);
output(3, 170) <= input(12);
output(3, 171) <= input(13);
output(3, 172) <= input(14);
output(3, 173) <= input(15);
output(3, 174) <= input(16);
output(3, 175) <= input(17);
output(3, 176) <= input(3);
output(3, 177) <= input(4);
output(3, 178) <= input(5);
output(3, 179) <= input(6);
output(3, 180) <= input(7);
output(3, 181) <= input(8);
output(3, 182) <= input(9);
output(3, 183) <= input(10);
output(3, 184) <= input(11);
output(3, 185) <= input(12);
output(3, 186) <= input(13);
output(3, 187) <= input(14);
output(3, 188) <= input(15);
output(3, 189) <= input(16);
output(3, 190) <= input(17);
output(3, 191) <= input(18);
output(3, 192) <= input(34);
output(3, 193) <= input(35);
output(3, 194) <= input(36);
output(3, 195) <= input(37);
output(3, 196) <= input(38);
output(3, 197) <= input(39);
output(3, 198) <= input(40);
output(3, 199) <= input(41);
output(3, 200) <= input(42);
output(3, 201) <= input(43);
output(3, 202) <= input(44);
output(3, 203) <= input(45);
output(3, 204) <= input(46);
output(3, 205) <= input(47);
output(3, 206) <= input(48);
output(3, 207) <= input(49);
output(3, 208) <= input(35);
output(3, 209) <= input(36);
output(3, 210) <= input(37);
output(3, 211) <= input(38);
output(3, 212) <= input(39);
output(3, 213) <= input(40);
output(3, 214) <= input(41);
output(3, 215) <= input(42);
output(3, 216) <= input(43);
output(3, 217) <= input(44);
output(3, 218) <= input(45);
output(3, 219) <= input(46);
output(3, 220) <= input(47);
output(3, 221) <= input(48);
output(3, 222) <= input(49);
output(3, 223) <= input(50);
output(3, 224) <= input(5);
output(3, 225) <= input(6);
output(3, 226) <= input(7);
output(3, 227) <= input(8);
output(3, 228) <= input(9);
output(3, 229) <= input(10);
output(3, 230) <= input(11);
output(3, 231) <= input(12);
output(3, 232) <= input(13);
output(3, 233) <= input(14);
output(3, 234) <= input(15);
output(3, 235) <= input(16);
output(3, 236) <= input(17);
output(3, 237) <= input(18);
output(3, 238) <= input(19);
output(3, 239) <= input(20);
output(3, 240) <= input(6);
output(3, 241) <= input(7);
output(3, 242) <= input(8);
output(3, 243) <= input(9);
output(3, 244) <= input(10);
output(3, 245) <= input(11);
output(3, 246) <= input(12);
output(3, 247) <= input(13);
output(3, 248) <= input(14);
output(3, 249) <= input(15);
output(3, 250) <= input(16);
output(3, 251) <= input(17);
output(3, 252) <= input(18);
output(3, 253) <= input(19);
output(3, 254) <= input(20);
output(3, 255) <= input(21);
output(4, 0) <= input(63);
output(4, 1) <= input(64);
output(4, 2) <= input(62);
output(4, 3) <= input(53);
output(4, 4) <= input(54);
output(4, 5) <= input(55);
output(4, 6) <= input(56);
output(4, 7) <= input(57);
output(4, 8) <= input(58);
output(4, 9) <= input(33);
output(4, 10) <= input(34);
output(4, 11) <= input(35);
output(4, 12) <= input(36);
output(4, 13) <= input(37);
output(4, 14) <= input(38);
output(4, 15) <= input(39);
output(4, 16) <= input(65);
output(4, 17) <= input(59);
output(4, 18) <= input(60);
output(4, 19) <= input(61);
output(4, 20) <= input(31);
output(4, 21) <= input(32);
output(4, 22) <= input(0);
output(4, 23) <= input(1);
output(4, 24) <= input(2);
output(4, 25) <= input(3);
output(4, 26) <= input(4);
output(4, 27) <= input(5);
output(4, 28) <= input(6);
output(4, 29) <= input(7);
output(4, 30) <= input(8);
output(4, 31) <= input(9);
output(4, 32) <= input(64);
output(4, 33) <= input(62);
output(4, 34) <= input(53);
output(4, 35) <= input(54);
output(4, 36) <= input(55);
output(4, 37) <= input(56);
output(4, 38) <= input(57);
output(4, 39) <= input(58);
output(4, 40) <= input(33);
output(4, 41) <= input(34);
output(4, 42) <= input(35);
output(4, 43) <= input(36);
output(4, 44) <= input(37);
output(4, 45) <= input(38);
output(4, 46) <= input(39);
output(4, 47) <= input(40);
output(4, 48) <= input(62);
output(4, 49) <= input(53);
output(4, 50) <= input(54);
output(4, 51) <= input(55);
output(4, 52) <= input(56);
output(4, 53) <= input(57);
output(4, 54) <= input(58);
output(4, 55) <= input(33);
output(4, 56) <= input(34);
output(4, 57) <= input(35);
output(4, 58) <= input(36);
output(4, 59) <= input(37);
output(4, 60) <= input(38);
output(4, 61) <= input(39);
output(4, 62) <= input(40);
output(4, 63) <= input(41);
output(4, 64) <= input(60);
output(4, 65) <= input(61);
output(4, 66) <= input(31);
output(4, 67) <= input(32);
output(4, 68) <= input(0);
output(4, 69) <= input(1);
output(4, 70) <= input(2);
output(4, 71) <= input(3);
output(4, 72) <= input(4);
output(4, 73) <= input(5);
output(4, 74) <= input(6);
output(4, 75) <= input(7);
output(4, 76) <= input(8);
output(4, 77) <= input(9);
output(4, 78) <= input(10);
output(4, 79) <= input(11);
output(4, 80) <= input(53);
output(4, 81) <= input(54);
output(4, 82) <= input(55);
output(4, 83) <= input(56);
output(4, 84) <= input(57);
output(4, 85) <= input(58);
output(4, 86) <= input(33);
output(4, 87) <= input(34);
output(4, 88) <= input(35);
output(4, 89) <= input(36);
output(4, 90) <= input(37);
output(4, 91) <= input(38);
output(4, 92) <= input(39);
output(4, 93) <= input(40);
output(4, 94) <= input(41);
output(4, 95) <= input(42);
output(4, 96) <= input(61);
output(4, 97) <= input(31);
output(4, 98) <= input(32);
output(4, 99) <= input(0);
output(4, 100) <= input(1);
output(4, 101) <= input(2);
output(4, 102) <= input(3);
output(4, 103) <= input(4);
output(4, 104) <= input(5);
output(4, 105) <= input(6);
output(4, 106) <= input(7);
output(4, 107) <= input(8);
output(4, 108) <= input(9);
output(4, 109) <= input(10);
output(4, 110) <= input(11);
output(4, 111) <= input(12);
output(4, 112) <= input(31);
output(4, 113) <= input(32);
output(4, 114) <= input(0);
output(4, 115) <= input(1);
output(4, 116) <= input(2);
output(4, 117) <= input(3);
output(4, 118) <= input(4);
output(4, 119) <= input(5);
output(4, 120) <= input(6);
output(4, 121) <= input(7);
output(4, 122) <= input(8);
output(4, 123) <= input(9);
output(4, 124) <= input(10);
output(4, 125) <= input(11);
output(4, 126) <= input(12);
output(4, 127) <= input(13);
output(4, 128) <= input(55);
output(4, 129) <= input(56);
output(4, 130) <= input(57);
output(4, 131) <= input(58);
output(4, 132) <= input(33);
output(4, 133) <= input(34);
output(4, 134) <= input(35);
output(4, 135) <= input(36);
output(4, 136) <= input(37);
output(4, 137) <= input(38);
output(4, 138) <= input(39);
output(4, 139) <= input(40);
output(4, 140) <= input(41);
output(4, 141) <= input(42);
output(4, 142) <= input(43);
output(4, 143) <= input(44);
output(4, 144) <= input(32);
output(4, 145) <= input(0);
output(4, 146) <= input(1);
output(4, 147) <= input(2);
output(4, 148) <= input(3);
output(4, 149) <= input(4);
output(4, 150) <= input(5);
output(4, 151) <= input(6);
output(4, 152) <= input(7);
output(4, 153) <= input(8);
output(4, 154) <= input(9);
output(4, 155) <= input(10);
output(4, 156) <= input(11);
output(4, 157) <= input(12);
output(4, 158) <= input(13);
output(4, 159) <= input(14);
output(4, 160) <= input(56);
output(4, 161) <= input(57);
output(4, 162) <= input(58);
output(4, 163) <= input(33);
output(4, 164) <= input(34);
output(4, 165) <= input(35);
output(4, 166) <= input(36);
output(4, 167) <= input(37);
output(4, 168) <= input(38);
output(4, 169) <= input(39);
output(4, 170) <= input(40);
output(4, 171) <= input(41);
output(4, 172) <= input(42);
output(4, 173) <= input(43);
output(4, 174) <= input(44);
output(4, 175) <= input(45);
output(4, 176) <= input(57);
output(4, 177) <= input(58);
output(4, 178) <= input(33);
output(4, 179) <= input(34);
output(4, 180) <= input(35);
output(4, 181) <= input(36);
output(4, 182) <= input(37);
output(4, 183) <= input(38);
output(4, 184) <= input(39);
output(4, 185) <= input(40);
output(4, 186) <= input(41);
output(4, 187) <= input(42);
output(4, 188) <= input(43);
output(4, 189) <= input(44);
output(4, 190) <= input(45);
output(4, 191) <= input(46);
output(4, 192) <= input(1);
output(4, 193) <= input(2);
output(4, 194) <= input(3);
output(4, 195) <= input(4);
output(4, 196) <= input(5);
output(4, 197) <= input(6);
output(4, 198) <= input(7);
output(4, 199) <= input(8);
output(4, 200) <= input(9);
output(4, 201) <= input(10);
output(4, 202) <= input(11);
output(4, 203) <= input(12);
output(4, 204) <= input(13);
output(4, 205) <= input(14);
output(4, 206) <= input(15);
output(4, 207) <= input(16);
output(4, 208) <= input(58);
output(4, 209) <= input(33);
output(4, 210) <= input(34);
output(4, 211) <= input(35);
output(4, 212) <= input(36);
output(4, 213) <= input(37);
output(4, 214) <= input(38);
output(4, 215) <= input(39);
output(4, 216) <= input(40);
output(4, 217) <= input(41);
output(4, 218) <= input(42);
output(4, 219) <= input(43);
output(4, 220) <= input(44);
output(4, 221) <= input(45);
output(4, 222) <= input(46);
output(4, 223) <= input(47);
output(4, 224) <= input(2);
output(4, 225) <= input(3);
output(4, 226) <= input(4);
output(4, 227) <= input(5);
output(4, 228) <= input(6);
output(4, 229) <= input(7);
output(4, 230) <= input(8);
output(4, 231) <= input(9);
output(4, 232) <= input(10);
output(4, 233) <= input(11);
output(4, 234) <= input(12);
output(4, 235) <= input(13);
output(4, 236) <= input(14);
output(4, 237) <= input(15);
output(4, 238) <= input(16);
output(4, 239) <= input(17);
output(4, 240) <= input(3);
output(4, 241) <= input(4);
output(4, 242) <= input(5);
output(4, 243) <= input(6);
output(4, 244) <= input(7);
output(4, 245) <= input(8);
output(4, 246) <= input(9);
output(4, 247) <= input(10);
output(4, 248) <= input(11);
output(4, 249) <= input(12);
output(4, 250) <= input(13);
output(4, 251) <= input(14);
output(4, 252) <= input(15);
output(4, 253) <= input(16);
output(4, 254) <= input(17);
output(4, 255) <= input(18);
output(5, 0) <= input(66);
output(5, 1) <= input(63);
output(5, 2) <= input(64);
output(5, 3) <= input(62);
output(5, 4) <= input(53);
output(5, 5) <= input(54);
output(5, 6) <= input(55);
output(5, 7) <= input(56);
output(5, 8) <= input(57);
output(5, 9) <= input(58);
output(5, 10) <= input(33);
output(5, 11) <= input(34);
output(5, 12) <= input(35);
output(5, 13) <= input(36);
output(5, 14) <= input(37);
output(5, 15) <= input(38);
output(5, 16) <= input(67);
output(5, 17) <= input(65);
output(5, 18) <= input(59);
output(5, 19) <= input(60);
output(5, 20) <= input(61);
output(5, 21) <= input(31);
output(5, 22) <= input(32);
output(5, 23) <= input(0);
output(5, 24) <= input(1);
output(5, 25) <= input(2);
output(5, 26) <= input(3);
output(5, 27) <= input(4);
output(5, 28) <= input(5);
output(5, 29) <= input(6);
output(5, 30) <= input(7);
output(5, 31) <= input(8);
output(5, 32) <= input(63);
output(5, 33) <= input(64);
output(5, 34) <= input(62);
output(5, 35) <= input(53);
output(5, 36) <= input(54);
output(5, 37) <= input(55);
output(5, 38) <= input(56);
output(5, 39) <= input(57);
output(5, 40) <= input(58);
output(5, 41) <= input(33);
output(5, 42) <= input(34);
output(5, 43) <= input(35);
output(5, 44) <= input(36);
output(5, 45) <= input(37);
output(5, 46) <= input(38);
output(5, 47) <= input(39);
output(5, 48) <= input(65);
output(5, 49) <= input(59);
output(5, 50) <= input(60);
output(5, 51) <= input(61);
output(5, 52) <= input(31);
output(5, 53) <= input(32);
output(5, 54) <= input(0);
output(5, 55) <= input(1);
output(5, 56) <= input(2);
output(5, 57) <= input(3);
output(5, 58) <= input(4);
output(5, 59) <= input(5);
output(5, 60) <= input(6);
output(5, 61) <= input(7);
output(5, 62) <= input(8);
output(5, 63) <= input(9);
output(5, 64) <= input(64);
output(5, 65) <= input(62);
output(5, 66) <= input(53);
output(5, 67) <= input(54);
output(5, 68) <= input(55);
output(5, 69) <= input(56);
output(5, 70) <= input(57);
output(5, 71) <= input(58);
output(5, 72) <= input(33);
output(5, 73) <= input(34);
output(5, 74) <= input(35);
output(5, 75) <= input(36);
output(5, 76) <= input(37);
output(5, 77) <= input(38);
output(5, 78) <= input(39);
output(5, 79) <= input(40);
output(5, 80) <= input(59);
output(5, 81) <= input(60);
output(5, 82) <= input(61);
output(5, 83) <= input(31);
output(5, 84) <= input(32);
output(5, 85) <= input(0);
output(5, 86) <= input(1);
output(5, 87) <= input(2);
output(5, 88) <= input(3);
output(5, 89) <= input(4);
output(5, 90) <= input(5);
output(5, 91) <= input(6);
output(5, 92) <= input(7);
output(5, 93) <= input(8);
output(5, 94) <= input(9);
output(5, 95) <= input(10);
output(5, 96) <= input(62);
output(5, 97) <= input(53);
output(5, 98) <= input(54);
output(5, 99) <= input(55);
output(5, 100) <= input(56);
output(5, 101) <= input(57);
output(5, 102) <= input(58);
output(5, 103) <= input(33);
output(5, 104) <= input(34);
output(5, 105) <= input(35);
output(5, 106) <= input(36);
output(5, 107) <= input(37);
output(5, 108) <= input(38);
output(5, 109) <= input(39);
output(5, 110) <= input(40);
output(5, 111) <= input(41);
output(5, 112) <= input(53);
output(5, 113) <= input(54);
output(5, 114) <= input(55);
output(5, 115) <= input(56);
output(5, 116) <= input(57);
output(5, 117) <= input(58);
output(5, 118) <= input(33);
output(5, 119) <= input(34);
output(5, 120) <= input(35);
output(5, 121) <= input(36);
output(5, 122) <= input(37);
output(5, 123) <= input(38);
output(5, 124) <= input(39);
output(5, 125) <= input(40);
output(5, 126) <= input(41);
output(5, 127) <= input(42);
output(5, 128) <= input(61);
output(5, 129) <= input(31);
output(5, 130) <= input(32);
output(5, 131) <= input(0);
output(5, 132) <= input(1);
output(5, 133) <= input(2);
output(5, 134) <= input(3);
output(5, 135) <= input(4);
output(5, 136) <= input(5);
output(5, 137) <= input(6);
output(5, 138) <= input(7);
output(5, 139) <= input(8);
output(5, 140) <= input(9);
output(5, 141) <= input(10);
output(5, 142) <= input(11);
output(5, 143) <= input(12);
output(5, 144) <= input(54);
output(5, 145) <= input(55);
output(5, 146) <= input(56);
output(5, 147) <= input(57);
output(5, 148) <= input(58);
output(5, 149) <= input(33);
output(5, 150) <= input(34);
output(5, 151) <= input(35);
output(5, 152) <= input(36);
output(5, 153) <= input(37);
output(5, 154) <= input(38);
output(5, 155) <= input(39);
output(5, 156) <= input(40);
output(5, 157) <= input(41);
output(5, 158) <= input(42);
output(5, 159) <= input(43);
output(5, 160) <= input(31);
output(5, 161) <= input(32);
output(5, 162) <= input(0);
output(5, 163) <= input(1);
output(5, 164) <= input(2);
output(5, 165) <= input(3);
output(5, 166) <= input(4);
output(5, 167) <= input(5);
output(5, 168) <= input(6);
output(5, 169) <= input(7);
output(5, 170) <= input(8);
output(5, 171) <= input(9);
output(5, 172) <= input(10);
output(5, 173) <= input(11);
output(5, 174) <= input(12);
output(5, 175) <= input(13);
output(5, 176) <= input(55);
output(5, 177) <= input(56);
output(5, 178) <= input(57);
output(5, 179) <= input(58);
output(5, 180) <= input(33);
output(5, 181) <= input(34);
output(5, 182) <= input(35);
output(5, 183) <= input(36);
output(5, 184) <= input(37);
output(5, 185) <= input(38);
output(5, 186) <= input(39);
output(5, 187) <= input(40);
output(5, 188) <= input(41);
output(5, 189) <= input(42);
output(5, 190) <= input(43);
output(5, 191) <= input(44);
output(5, 192) <= input(32);
output(5, 193) <= input(0);
output(5, 194) <= input(1);
output(5, 195) <= input(2);
output(5, 196) <= input(3);
output(5, 197) <= input(4);
output(5, 198) <= input(5);
output(5, 199) <= input(6);
output(5, 200) <= input(7);
output(5, 201) <= input(8);
output(5, 202) <= input(9);
output(5, 203) <= input(10);
output(5, 204) <= input(11);
output(5, 205) <= input(12);
output(5, 206) <= input(13);
output(5, 207) <= input(14);
output(5, 208) <= input(56);
output(5, 209) <= input(57);
output(5, 210) <= input(58);
output(5, 211) <= input(33);
output(5, 212) <= input(34);
output(5, 213) <= input(35);
output(5, 214) <= input(36);
output(5, 215) <= input(37);
output(5, 216) <= input(38);
output(5, 217) <= input(39);
output(5, 218) <= input(40);
output(5, 219) <= input(41);
output(5, 220) <= input(42);
output(5, 221) <= input(43);
output(5, 222) <= input(44);
output(5, 223) <= input(45);
output(5, 224) <= input(0);
output(5, 225) <= input(1);
output(5, 226) <= input(2);
output(5, 227) <= input(3);
output(5, 228) <= input(4);
output(5, 229) <= input(5);
output(5, 230) <= input(6);
output(5, 231) <= input(7);
output(5, 232) <= input(8);
output(5, 233) <= input(9);
output(5, 234) <= input(10);
output(5, 235) <= input(11);
output(5, 236) <= input(12);
output(5, 237) <= input(13);
output(5, 238) <= input(14);
output(5, 239) <= input(15);
output(5, 240) <= input(1);
output(5, 241) <= input(2);
output(5, 242) <= input(3);
output(5, 243) <= input(4);
output(5, 244) <= input(5);
output(5, 245) <= input(6);
output(5, 246) <= input(7);
output(5, 247) <= input(8);
output(5, 248) <= input(9);
output(5, 249) <= input(10);
output(5, 250) <= input(11);
output(5, 251) <= input(12);
output(5, 252) <= input(13);
output(5, 253) <= input(14);
output(5, 254) <= input(15);
output(5, 255) <= input(16);
when "0001" =>
output(0, 0) <= input(0);
output(0, 1) <= input(1);
output(0, 2) <= input(2);
output(0, 3) <= input(3);
output(0, 4) <= input(4);
output(0, 5) <= input(5);
output(0, 6) <= input(6);
output(0, 7) <= input(7);
output(0, 8) <= input(8);
output(0, 9) <= input(9);
output(0, 10) <= input(10);
output(0, 11) <= input(11);
output(0, 12) <= input(12);
output(0, 13) <= input(13);
output(0, 14) <= input(14);
output(0, 15) <= input(15);
output(0, 16) <= input(16);
output(0, 17) <= input(17);
output(0, 18) <= input(18);
output(0, 19) <= input(19);
output(0, 20) <= input(20);
output(0, 21) <= input(21);
output(0, 22) <= input(22);
output(0, 23) <= input(23);
output(0, 24) <= input(24);
output(0, 25) <= input(25);
output(0, 26) <= input(26);
output(0, 27) <= input(27);
output(0, 28) <= input(28);
output(0, 29) <= input(29);
output(0, 30) <= input(30);
output(0, 31) <= input(31);
output(0, 32) <= input(1);
output(0, 33) <= input(2);
output(0, 34) <= input(3);
output(0, 35) <= input(4);
output(0, 36) <= input(5);
output(0, 37) <= input(6);
output(0, 38) <= input(7);
output(0, 39) <= input(8);
output(0, 40) <= input(9);
output(0, 41) <= input(10);
output(0, 42) <= input(11);
output(0, 43) <= input(12);
output(0, 44) <= input(13);
output(0, 45) <= input(14);
output(0, 46) <= input(15);
output(0, 47) <= input(32);
output(0, 48) <= input(17);
output(0, 49) <= input(18);
output(0, 50) <= input(19);
output(0, 51) <= input(20);
output(0, 52) <= input(21);
output(0, 53) <= input(22);
output(0, 54) <= input(23);
output(0, 55) <= input(24);
output(0, 56) <= input(25);
output(0, 57) <= input(26);
output(0, 58) <= input(27);
output(0, 59) <= input(28);
output(0, 60) <= input(29);
output(0, 61) <= input(30);
output(0, 62) <= input(31);
output(0, 63) <= input(33);
output(0, 64) <= input(2);
output(0, 65) <= input(3);
output(0, 66) <= input(4);
output(0, 67) <= input(5);
output(0, 68) <= input(6);
output(0, 69) <= input(7);
output(0, 70) <= input(8);
output(0, 71) <= input(9);
output(0, 72) <= input(10);
output(0, 73) <= input(11);
output(0, 74) <= input(12);
output(0, 75) <= input(13);
output(0, 76) <= input(14);
output(0, 77) <= input(15);
output(0, 78) <= input(32);
output(0, 79) <= input(34);
output(0, 80) <= input(18);
output(0, 81) <= input(19);
output(0, 82) <= input(20);
output(0, 83) <= input(21);
output(0, 84) <= input(22);
output(0, 85) <= input(23);
output(0, 86) <= input(24);
output(0, 87) <= input(25);
output(0, 88) <= input(26);
output(0, 89) <= input(27);
output(0, 90) <= input(28);
output(0, 91) <= input(29);
output(0, 92) <= input(30);
output(0, 93) <= input(31);
output(0, 94) <= input(33);
output(0, 95) <= input(35);
output(0, 96) <= input(3);
output(0, 97) <= input(4);
output(0, 98) <= input(5);
output(0, 99) <= input(6);
output(0, 100) <= input(7);
output(0, 101) <= input(8);
output(0, 102) <= input(9);
output(0, 103) <= input(10);
output(0, 104) <= input(11);
output(0, 105) <= input(12);
output(0, 106) <= input(13);
output(0, 107) <= input(14);
output(0, 108) <= input(15);
output(0, 109) <= input(32);
output(0, 110) <= input(34);
output(0, 111) <= input(36);
output(0, 112) <= input(19);
output(0, 113) <= input(20);
output(0, 114) <= input(21);
output(0, 115) <= input(22);
output(0, 116) <= input(23);
output(0, 117) <= input(24);
output(0, 118) <= input(25);
output(0, 119) <= input(26);
output(0, 120) <= input(27);
output(0, 121) <= input(28);
output(0, 122) <= input(29);
output(0, 123) <= input(30);
output(0, 124) <= input(31);
output(0, 125) <= input(33);
output(0, 126) <= input(35);
output(0, 127) <= input(37);
output(0, 128) <= input(4);
output(0, 129) <= input(5);
output(0, 130) <= input(6);
output(0, 131) <= input(7);
output(0, 132) <= input(8);
output(0, 133) <= input(9);
output(0, 134) <= input(10);
output(0, 135) <= input(11);
output(0, 136) <= input(12);
output(0, 137) <= input(13);
output(0, 138) <= input(14);
output(0, 139) <= input(15);
output(0, 140) <= input(32);
output(0, 141) <= input(34);
output(0, 142) <= input(36);
output(0, 143) <= input(38);
output(0, 144) <= input(20);
output(0, 145) <= input(21);
output(0, 146) <= input(22);
output(0, 147) <= input(23);
output(0, 148) <= input(24);
output(0, 149) <= input(25);
output(0, 150) <= input(26);
output(0, 151) <= input(27);
output(0, 152) <= input(28);
output(0, 153) <= input(29);
output(0, 154) <= input(30);
output(0, 155) <= input(31);
output(0, 156) <= input(33);
output(0, 157) <= input(35);
output(0, 158) <= input(37);
output(0, 159) <= input(39);
output(0, 160) <= input(5);
output(0, 161) <= input(6);
output(0, 162) <= input(7);
output(0, 163) <= input(8);
output(0, 164) <= input(9);
output(0, 165) <= input(10);
output(0, 166) <= input(11);
output(0, 167) <= input(12);
output(0, 168) <= input(13);
output(0, 169) <= input(14);
output(0, 170) <= input(15);
output(0, 171) <= input(32);
output(0, 172) <= input(34);
output(0, 173) <= input(36);
output(0, 174) <= input(38);
output(0, 175) <= input(40);
output(0, 176) <= input(21);
output(0, 177) <= input(22);
output(0, 178) <= input(23);
output(0, 179) <= input(24);
output(0, 180) <= input(25);
output(0, 181) <= input(26);
output(0, 182) <= input(27);
output(0, 183) <= input(28);
output(0, 184) <= input(29);
output(0, 185) <= input(30);
output(0, 186) <= input(31);
output(0, 187) <= input(33);
output(0, 188) <= input(35);
output(0, 189) <= input(37);
output(0, 190) <= input(39);
output(0, 191) <= input(41);
output(0, 192) <= input(6);
output(0, 193) <= input(7);
output(0, 194) <= input(8);
output(0, 195) <= input(9);
output(0, 196) <= input(10);
output(0, 197) <= input(11);
output(0, 198) <= input(12);
output(0, 199) <= input(13);
output(0, 200) <= input(14);
output(0, 201) <= input(15);
output(0, 202) <= input(32);
output(0, 203) <= input(34);
output(0, 204) <= input(36);
output(0, 205) <= input(38);
output(0, 206) <= input(40);
output(0, 207) <= input(42);
output(0, 208) <= input(22);
output(0, 209) <= input(23);
output(0, 210) <= input(24);
output(0, 211) <= input(25);
output(0, 212) <= input(26);
output(0, 213) <= input(27);
output(0, 214) <= input(28);
output(0, 215) <= input(29);
output(0, 216) <= input(30);
output(0, 217) <= input(31);
output(0, 218) <= input(33);
output(0, 219) <= input(35);
output(0, 220) <= input(37);
output(0, 221) <= input(39);
output(0, 222) <= input(41);
output(0, 223) <= input(43);
output(0, 224) <= input(7);
output(0, 225) <= input(8);
output(0, 226) <= input(9);
output(0, 227) <= input(10);
output(0, 228) <= input(11);
output(0, 229) <= input(12);
output(0, 230) <= input(13);
output(0, 231) <= input(14);
output(0, 232) <= input(15);
output(0, 233) <= input(32);
output(0, 234) <= input(34);
output(0, 235) <= input(36);
output(0, 236) <= input(38);
output(0, 237) <= input(40);
output(0, 238) <= input(42);
output(0, 239) <= input(44);
output(0, 240) <= input(23);
output(0, 241) <= input(24);
output(0, 242) <= input(25);
output(0, 243) <= input(26);
output(0, 244) <= input(27);
output(0, 245) <= input(28);
output(0, 246) <= input(29);
output(0, 247) <= input(30);
output(0, 248) <= input(31);
output(0, 249) <= input(33);
output(0, 250) <= input(35);
output(0, 251) <= input(37);
output(0, 252) <= input(39);
output(0, 253) <= input(41);
output(0, 254) <= input(43);
output(0, 255) <= input(45);
output(1, 0) <= input(46);
output(1, 1) <= input(47);
output(1, 2) <= input(16);
output(1, 3) <= input(17);
output(1, 4) <= input(18);
output(1, 5) <= input(19);
output(1, 6) <= input(20);
output(1, 7) <= input(21);
output(1, 8) <= input(22);
output(1, 9) <= input(23);
output(1, 10) <= input(24);
output(1, 11) <= input(25);
output(1, 12) <= input(26);
output(1, 13) <= input(27);
output(1, 14) <= input(28);
output(1, 15) <= input(29);
output(1, 16) <= input(48);
output(1, 17) <= input(0);
output(1, 18) <= input(1);
output(1, 19) <= input(2);
output(1, 20) <= input(3);
output(1, 21) <= input(4);
output(1, 22) <= input(5);
output(1, 23) <= input(6);
output(1, 24) <= input(7);
output(1, 25) <= input(8);
output(1, 26) <= input(9);
output(1, 27) <= input(10);
output(1, 28) <= input(11);
output(1, 29) <= input(12);
output(1, 30) <= input(13);
output(1, 31) <= input(14);
output(1, 32) <= input(47);
output(1, 33) <= input(16);
output(1, 34) <= input(17);
output(1, 35) <= input(18);
output(1, 36) <= input(19);
output(1, 37) <= input(20);
output(1, 38) <= input(21);
output(1, 39) <= input(22);
output(1, 40) <= input(23);
output(1, 41) <= input(24);
output(1, 42) <= input(25);
output(1, 43) <= input(26);
output(1, 44) <= input(27);
output(1, 45) <= input(28);
output(1, 46) <= input(29);
output(1, 47) <= input(30);
output(1, 48) <= input(0);
output(1, 49) <= input(1);
output(1, 50) <= input(2);
output(1, 51) <= input(3);
output(1, 52) <= input(4);
output(1, 53) <= input(5);
output(1, 54) <= input(6);
output(1, 55) <= input(7);
output(1, 56) <= input(8);
output(1, 57) <= input(9);
output(1, 58) <= input(10);
output(1, 59) <= input(11);
output(1, 60) <= input(12);
output(1, 61) <= input(13);
output(1, 62) <= input(14);
output(1, 63) <= input(15);
output(1, 64) <= input(16);
output(1, 65) <= input(17);
output(1, 66) <= input(18);
output(1, 67) <= input(19);
output(1, 68) <= input(20);
output(1, 69) <= input(21);
output(1, 70) <= input(22);
output(1, 71) <= input(23);
output(1, 72) <= input(24);
output(1, 73) <= input(25);
output(1, 74) <= input(26);
output(1, 75) <= input(27);
output(1, 76) <= input(28);
output(1, 77) <= input(29);
output(1, 78) <= input(30);
output(1, 79) <= input(31);
output(1, 80) <= input(1);
output(1, 81) <= input(2);
output(1, 82) <= input(3);
output(1, 83) <= input(4);
output(1, 84) <= input(5);
output(1, 85) <= input(6);
output(1, 86) <= input(7);
output(1, 87) <= input(8);
output(1, 88) <= input(9);
output(1, 89) <= input(10);
output(1, 90) <= input(11);
output(1, 91) <= input(12);
output(1, 92) <= input(13);
output(1, 93) <= input(14);
output(1, 94) <= input(15);
output(1, 95) <= input(32);
output(1, 96) <= input(17);
output(1, 97) <= input(18);
output(1, 98) <= input(19);
output(1, 99) <= input(20);
output(1, 100) <= input(21);
output(1, 101) <= input(22);
output(1, 102) <= input(23);
output(1, 103) <= input(24);
output(1, 104) <= input(25);
output(1, 105) <= input(26);
output(1, 106) <= input(27);
output(1, 107) <= input(28);
output(1, 108) <= input(29);
output(1, 109) <= input(30);
output(1, 110) <= input(31);
output(1, 111) <= input(33);
output(1, 112) <= input(2);
output(1, 113) <= input(3);
output(1, 114) <= input(4);
output(1, 115) <= input(5);
output(1, 116) <= input(6);
output(1, 117) <= input(7);
output(1, 118) <= input(8);
output(1, 119) <= input(9);
output(1, 120) <= input(10);
output(1, 121) <= input(11);
output(1, 122) <= input(12);
output(1, 123) <= input(13);
output(1, 124) <= input(14);
output(1, 125) <= input(15);
output(1, 126) <= input(32);
output(1, 127) <= input(34);
output(1, 128) <= input(2);
output(1, 129) <= input(3);
output(1, 130) <= input(4);
output(1, 131) <= input(5);
output(1, 132) <= input(6);
output(1, 133) <= input(7);
output(1, 134) <= input(8);
output(1, 135) <= input(9);
output(1, 136) <= input(10);
output(1, 137) <= input(11);
output(1, 138) <= input(12);
output(1, 139) <= input(13);
output(1, 140) <= input(14);
output(1, 141) <= input(15);
output(1, 142) <= input(32);
output(1, 143) <= input(34);
output(1, 144) <= input(18);
output(1, 145) <= input(19);
output(1, 146) <= input(20);
output(1, 147) <= input(21);
output(1, 148) <= input(22);
output(1, 149) <= input(23);
output(1, 150) <= input(24);
output(1, 151) <= input(25);
output(1, 152) <= input(26);
output(1, 153) <= input(27);
output(1, 154) <= input(28);
output(1, 155) <= input(29);
output(1, 156) <= input(30);
output(1, 157) <= input(31);
output(1, 158) <= input(33);
output(1, 159) <= input(35);
output(1, 160) <= input(3);
output(1, 161) <= input(4);
output(1, 162) <= input(5);
output(1, 163) <= input(6);
output(1, 164) <= input(7);
output(1, 165) <= input(8);
output(1, 166) <= input(9);
output(1, 167) <= input(10);
output(1, 168) <= input(11);
output(1, 169) <= input(12);
output(1, 170) <= input(13);
output(1, 171) <= input(14);
output(1, 172) <= input(15);
output(1, 173) <= input(32);
output(1, 174) <= input(34);
output(1, 175) <= input(36);
output(1, 176) <= input(19);
output(1, 177) <= input(20);
output(1, 178) <= input(21);
output(1, 179) <= input(22);
output(1, 180) <= input(23);
output(1, 181) <= input(24);
output(1, 182) <= input(25);
output(1, 183) <= input(26);
output(1, 184) <= input(27);
output(1, 185) <= input(28);
output(1, 186) <= input(29);
output(1, 187) <= input(30);
output(1, 188) <= input(31);
output(1, 189) <= input(33);
output(1, 190) <= input(35);
output(1, 191) <= input(37);
output(1, 192) <= input(4);
output(1, 193) <= input(5);
output(1, 194) <= input(6);
output(1, 195) <= input(7);
output(1, 196) <= input(8);
output(1, 197) <= input(9);
output(1, 198) <= input(10);
output(1, 199) <= input(11);
output(1, 200) <= input(12);
output(1, 201) <= input(13);
output(1, 202) <= input(14);
output(1, 203) <= input(15);
output(1, 204) <= input(32);
output(1, 205) <= input(34);
output(1, 206) <= input(36);
output(1, 207) <= input(38);
output(1, 208) <= input(20);
output(1, 209) <= input(21);
output(1, 210) <= input(22);
output(1, 211) <= input(23);
output(1, 212) <= input(24);
output(1, 213) <= input(25);
output(1, 214) <= input(26);
output(1, 215) <= input(27);
output(1, 216) <= input(28);
output(1, 217) <= input(29);
output(1, 218) <= input(30);
output(1, 219) <= input(31);
output(1, 220) <= input(33);
output(1, 221) <= input(35);
output(1, 222) <= input(37);
output(1, 223) <= input(39);
output(1, 224) <= input(5);
output(1, 225) <= input(6);
output(1, 226) <= input(7);
output(1, 227) <= input(8);
output(1, 228) <= input(9);
output(1, 229) <= input(10);
output(1, 230) <= input(11);
output(1, 231) <= input(12);
output(1, 232) <= input(13);
output(1, 233) <= input(14);
output(1, 234) <= input(15);
output(1, 235) <= input(32);
output(1, 236) <= input(34);
output(1, 237) <= input(36);
output(1, 238) <= input(38);
output(1, 239) <= input(40);
output(1, 240) <= input(21);
output(1, 241) <= input(22);
output(1, 242) <= input(23);
output(1, 243) <= input(24);
output(1, 244) <= input(25);
output(1, 245) <= input(26);
output(1, 246) <= input(27);
output(1, 247) <= input(28);
output(1, 248) <= input(29);
output(1, 249) <= input(30);
output(1, 250) <= input(31);
output(1, 251) <= input(33);
output(1, 252) <= input(35);
output(1, 253) <= input(37);
output(1, 254) <= input(39);
output(1, 255) <= input(41);
output(2, 0) <= input(49);
output(2, 1) <= input(46);
output(2, 2) <= input(47);
output(2, 3) <= input(16);
output(2, 4) <= input(17);
output(2, 5) <= input(18);
output(2, 6) <= input(19);
output(2, 7) <= input(20);
output(2, 8) <= input(21);
output(2, 9) <= input(22);
output(2, 10) <= input(23);
output(2, 11) <= input(24);
output(2, 12) <= input(25);
output(2, 13) <= input(26);
output(2, 14) <= input(27);
output(2, 15) <= input(28);
output(2, 16) <= input(50);
output(2, 17) <= input(48);
output(2, 18) <= input(0);
output(2, 19) <= input(1);
output(2, 20) <= input(2);
output(2, 21) <= input(3);
output(2, 22) <= input(4);
output(2, 23) <= input(5);
output(2, 24) <= input(6);
output(2, 25) <= input(7);
output(2, 26) <= input(8);
output(2, 27) <= input(9);
output(2, 28) <= input(10);
output(2, 29) <= input(11);
output(2, 30) <= input(12);
output(2, 31) <= input(13);
output(2, 32) <= input(46);
output(2, 33) <= input(47);
output(2, 34) <= input(16);
output(2, 35) <= input(17);
output(2, 36) <= input(18);
output(2, 37) <= input(19);
output(2, 38) <= input(20);
output(2, 39) <= input(21);
output(2, 40) <= input(22);
output(2, 41) <= input(23);
output(2, 42) <= input(24);
output(2, 43) <= input(25);
output(2, 44) <= input(26);
output(2, 45) <= input(27);
output(2, 46) <= input(28);
output(2, 47) <= input(29);
output(2, 48) <= input(48);
output(2, 49) <= input(0);
output(2, 50) <= input(1);
output(2, 51) <= input(2);
output(2, 52) <= input(3);
output(2, 53) <= input(4);
output(2, 54) <= input(5);
output(2, 55) <= input(6);
output(2, 56) <= input(7);
output(2, 57) <= input(8);
output(2, 58) <= input(9);
output(2, 59) <= input(10);
output(2, 60) <= input(11);
output(2, 61) <= input(12);
output(2, 62) <= input(13);
output(2, 63) <= input(14);
output(2, 64) <= input(48);
output(2, 65) <= input(0);
output(2, 66) <= input(1);
output(2, 67) <= input(2);
output(2, 68) <= input(3);
output(2, 69) <= input(4);
output(2, 70) <= input(5);
output(2, 71) <= input(6);
output(2, 72) <= input(7);
output(2, 73) <= input(8);
output(2, 74) <= input(9);
output(2, 75) <= input(10);
output(2, 76) <= input(11);
output(2, 77) <= input(12);
output(2, 78) <= input(13);
output(2, 79) <= input(14);
output(2, 80) <= input(47);
output(2, 81) <= input(16);
output(2, 82) <= input(17);
output(2, 83) <= input(18);
output(2, 84) <= input(19);
output(2, 85) <= input(20);
output(2, 86) <= input(21);
output(2, 87) <= input(22);
output(2, 88) <= input(23);
output(2, 89) <= input(24);
output(2, 90) <= input(25);
output(2, 91) <= input(26);
output(2, 92) <= input(27);
output(2, 93) <= input(28);
output(2, 94) <= input(29);
output(2, 95) <= input(30);
output(2, 96) <= input(0);
output(2, 97) <= input(1);
output(2, 98) <= input(2);
output(2, 99) <= input(3);
output(2, 100) <= input(4);
output(2, 101) <= input(5);
output(2, 102) <= input(6);
output(2, 103) <= input(7);
output(2, 104) <= input(8);
output(2, 105) <= input(9);
output(2, 106) <= input(10);
output(2, 107) <= input(11);
output(2, 108) <= input(12);
output(2, 109) <= input(13);
output(2, 110) <= input(14);
output(2, 111) <= input(15);
output(2, 112) <= input(16);
output(2, 113) <= input(17);
output(2, 114) <= input(18);
output(2, 115) <= input(19);
output(2, 116) <= input(20);
output(2, 117) <= input(21);
output(2, 118) <= input(22);
output(2, 119) <= input(23);
output(2, 120) <= input(24);
output(2, 121) <= input(25);
output(2, 122) <= input(26);
output(2, 123) <= input(27);
output(2, 124) <= input(28);
output(2, 125) <= input(29);
output(2, 126) <= input(30);
output(2, 127) <= input(31);
output(2, 128) <= input(16);
output(2, 129) <= input(17);
output(2, 130) <= input(18);
output(2, 131) <= input(19);
output(2, 132) <= input(20);
output(2, 133) <= input(21);
output(2, 134) <= input(22);
output(2, 135) <= input(23);
output(2, 136) <= input(24);
output(2, 137) <= input(25);
output(2, 138) <= input(26);
output(2, 139) <= input(27);
output(2, 140) <= input(28);
output(2, 141) <= input(29);
output(2, 142) <= input(30);
output(2, 143) <= input(31);
output(2, 144) <= input(1);
output(2, 145) <= input(2);
output(2, 146) <= input(3);
output(2, 147) <= input(4);
output(2, 148) <= input(5);
output(2, 149) <= input(6);
output(2, 150) <= input(7);
output(2, 151) <= input(8);
output(2, 152) <= input(9);
output(2, 153) <= input(10);
output(2, 154) <= input(11);
output(2, 155) <= input(12);
output(2, 156) <= input(13);
output(2, 157) <= input(14);
output(2, 158) <= input(15);
output(2, 159) <= input(32);
output(2, 160) <= input(17);
output(2, 161) <= input(18);
output(2, 162) <= input(19);
output(2, 163) <= input(20);
output(2, 164) <= input(21);
output(2, 165) <= input(22);
output(2, 166) <= input(23);
output(2, 167) <= input(24);
output(2, 168) <= input(25);
output(2, 169) <= input(26);
output(2, 170) <= input(27);
output(2, 171) <= input(28);
output(2, 172) <= input(29);
output(2, 173) <= input(30);
output(2, 174) <= input(31);
output(2, 175) <= input(33);
output(2, 176) <= input(2);
output(2, 177) <= input(3);
output(2, 178) <= input(4);
output(2, 179) <= input(5);
output(2, 180) <= input(6);
output(2, 181) <= input(7);
output(2, 182) <= input(8);
output(2, 183) <= input(9);
output(2, 184) <= input(10);
output(2, 185) <= input(11);
output(2, 186) <= input(12);
output(2, 187) <= input(13);
output(2, 188) <= input(14);
output(2, 189) <= input(15);
output(2, 190) <= input(32);
output(2, 191) <= input(34);
output(2, 192) <= input(2);
output(2, 193) <= input(3);
output(2, 194) <= input(4);
output(2, 195) <= input(5);
output(2, 196) <= input(6);
output(2, 197) <= input(7);
output(2, 198) <= input(8);
output(2, 199) <= input(9);
output(2, 200) <= input(10);
output(2, 201) <= input(11);
output(2, 202) <= input(12);
output(2, 203) <= input(13);
output(2, 204) <= input(14);
output(2, 205) <= input(15);
output(2, 206) <= input(32);
output(2, 207) <= input(34);
output(2, 208) <= input(18);
output(2, 209) <= input(19);
output(2, 210) <= input(20);
output(2, 211) <= input(21);
output(2, 212) <= input(22);
output(2, 213) <= input(23);
output(2, 214) <= input(24);
output(2, 215) <= input(25);
output(2, 216) <= input(26);
output(2, 217) <= input(27);
output(2, 218) <= input(28);
output(2, 219) <= input(29);
output(2, 220) <= input(30);
output(2, 221) <= input(31);
output(2, 222) <= input(33);
output(2, 223) <= input(35);
output(2, 224) <= input(3);
output(2, 225) <= input(4);
output(2, 226) <= input(5);
output(2, 227) <= input(6);
output(2, 228) <= input(7);
output(2, 229) <= input(8);
output(2, 230) <= input(9);
output(2, 231) <= input(10);
output(2, 232) <= input(11);
output(2, 233) <= input(12);
output(2, 234) <= input(13);
output(2, 235) <= input(14);
output(2, 236) <= input(15);
output(2, 237) <= input(32);
output(2, 238) <= input(34);
output(2, 239) <= input(36);
output(2, 240) <= input(19);
output(2, 241) <= input(20);
output(2, 242) <= input(21);
output(2, 243) <= input(22);
output(2, 244) <= input(23);
output(2, 245) <= input(24);
output(2, 246) <= input(25);
output(2, 247) <= input(26);
output(2, 248) <= input(27);
output(2, 249) <= input(28);
output(2, 250) <= input(29);
output(2, 251) <= input(30);
output(2, 252) <= input(31);
output(2, 253) <= input(33);
output(2, 254) <= input(35);
output(2, 255) <= input(37);
output(3, 0) <= input(51);
output(3, 1) <= input(49);
output(3, 2) <= input(46);
output(3, 3) <= input(47);
output(3, 4) <= input(16);
output(3, 5) <= input(17);
output(3, 6) <= input(18);
output(3, 7) <= input(19);
output(3, 8) <= input(20);
output(3, 9) <= input(21);
output(3, 10) <= input(22);
output(3, 11) <= input(23);
output(3, 12) <= input(24);
output(3, 13) <= input(25);
output(3, 14) <= input(26);
output(3, 15) <= input(27);
output(3, 16) <= input(52);
output(3, 17) <= input(50);
output(3, 18) <= input(48);
output(3, 19) <= input(0);
output(3, 20) <= input(1);
output(3, 21) <= input(2);
output(3, 22) <= input(3);
output(3, 23) <= input(4);
output(3, 24) <= input(5);
output(3, 25) <= input(6);
output(3, 26) <= input(7);
output(3, 27) <= input(8);
output(3, 28) <= input(9);
output(3, 29) <= input(10);
output(3, 30) <= input(11);
output(3, 31) <= input(12);
output(3, 32) <= input(52);
output(3, 33) <= input(50);
output(3, 34) <= input(48);
output(3, 35) <= input(0);
output(3, 36) <= input(1);
output(3, 37) <= input(2);
output(3, 38) <= input(3);
output(3, 39) <= input(4);
output(3, 40) <= input(5);
output(3, 41) <= input(6);
output(3, 42) <= input(7);
output(3, 43) <= input(8);
output(3, 44) <= input(9);
output(3, 45) <= input(10);
output(3, 46) <= input(11);
output(3, 47) <= input(12);
output(3, 48) <= input(49);
output(3, 49) <= input(46);
output(3, 50) <= input(47);
output(3, 51) <= input(16);
output(3, 52) <= input(17);
output(3, 53) <= input(18);
output(3, 54) <= input(19);
output(3, 55) <= input(20);
output(3, 56) <= input(21);
output(3, 57) <= input(22);
output(3, 58) <= input(23);
output(3, 59) <= input(24);
output(3, 60) <= input(25);
output(3, 61) <= input(26);
output(3, 62) <= input(27);
output(3, 63) <= input(28);
output(3, 64) <= input(50);
output(3, 65) <= input(48);
output(3, 66) <= input(0);
output(3, 67) <= input(1);
output(3, 68) <= input(2);
output(3, 69) <= input(3);
output(3, 70) <= input(4);
output(3, 71) <= input(5);
output(3, 72) <= input(6);
output(3, 73) <= input(7);
output(3, 74) <= input(8);
output(3, 75) <= input(9);
output(3, 76) <= input(10);
output(3, 77) <= input(11);
output(3, 78) <= input(12);
output(3, 79) <= input(13);
output(3, 80) <= input(50);
output(3, 81) <= input(48);
output(3, 82) <= input(0);
output(3, 83) <= input(1);
output(3, 84) <= input(2);
output(3, 85) <= input(3);
output(3, 86) <= input(4);
output(3, 87) <= input(5);
output(3, 88) <= input(6);
output(3, 89) <= input(7);
output(3, 90) <= input(8);
output(3, 91) <= input(9);
output(3, 92) <= input(10);
output(3, 93) <= input(11);
output(3, 94) <= input(12);
output(3, 95) <= input(13);
output(3, 96) <= input(46);
output(3, 97) <= input(47);
output(3, 98) <= input(16);
output(3, 99) <= input(17);
output(3, 100) <= input(18);
output(3, 101) <= input(19);
output(3, 102) <= input(20);
output(3, 103) <= input(21);
output(3, 104) <= input(22);
output(3, 105) <= input(23);
output(3, 106) <= input(24);
output(3, 107) <= input(25);
output(3, 108) <= input(26);
output(3, 109) <= input(27);
output(3, 110) <= input(28);
output(3, 111) <= input(29);
output(3, 112) <= input(48);
output(3, 113) <= input(0);
output(3, 114) <= input(1);
output(3, 115) <= input(2);
output(3, 116) <= input(3);
output(3, 117) <= input(4);
output(3, 118) <= input(5);
output(3, 119) <= input(6);
output(3, 120) <= input(7);
output(3, 121) <= input(8);
output(3, 122) <= input(9);
output(3, 123) <= input(10);
output(3, 124) <= input(11);
output(3, 125) <= input(12);
output(3, 126) <= input(13);
output(3, 127) <= input(14);
output(3, 128) <= input(48);
output(3, 129) <= input(0);
output(3, 130) <= input(1);
output(3, 131) <= input(2);
output(3, 132) <= input(3);
output(3, 133) <= input(4);
output(3, 134) <= input(5);
output(3, 135) <= input(6);
output(3, 136) <= input(7);
output(3, 137) <= input(8);
output(3, 138) <= input(9);
output(3, 139) <= input(10);
output(3, 140) <= input(11);
output(3, 141) <= input(12);
output(3, 142) <= input(13);
output(3, 143) <= input(14);
output(3, 144) <= input(47);
output(3, 145) <= input(16);
output(3, 146) <= input(17);
output(3, 147) <= input(18);
output(3, 148) <= input(19);
output(3, 149) <= input(20);
output(3, 150) <= input(21);
output(3, 151) <= input(22);
output(3, 152) <= input(23);
output(3, 153) <= input(24);
output(3, 154) <= input(25);
output(3, 155) <= input(26);
output(3, 156) <= input(27);
output(3, 157) <= input(28);
output(3, 158) <= input(29);
output(3, 159) <= input(30);
output(3, 160) <= input(47);
output(3, 161) <= input(16);
output(3, 162) <= input(17);
output(3, 163) <= input(18);
output(3, 164) <= input(19);
output(3, 165) <= input(20);
output(3, 166) <= input(21);
output(3, 167) <= input(22);
output(3, 168) <= input(23);
output(3, 169) <= input(24);
output(3, 170) <= input(25);
output(3, 171) <= input(26);
output(3, 172) <= input(27);
output(3, 173) <= input(28);
output(3, 174) <= input(29);
output(3, 175) <= input(30);
output(3, 176) <= input(0);
output(3, 177) <= input(1);
output(3, 178) <= input(2);
output(3, 179) <= input(3);
output(3, 180) <= input(4);
output(3, 181) <= input(5);
output(3, 182) <= input(6);
output(3, 183) <= input(7);
output(3, 184) <= input(8);
output(3, 185) <= input(9);
output(3, 186) <= input(10);
output(3, 187) <= input(11);
output(3, 188) <= input(12);
output(3, 189) <= input(13);
output(3, 190) <= input(14);
output(3, 191) <= input(15);
output(3, 192) <= input(16);
output(3, 193) <= input(17);
output(3, 194) <= input(18);
output(3, 195) <= input(19);
output(3, 196) <= input(20);
output(3, 197) <= input(21);
output(3, 198) <= input(22);
output(3, 199) <= input(23);
output(3, 200) <= input(24);
output(3, 201) <= input(25);
output(3, 202) <= input(26);
output(3, 203) <= input(27);
output(3, 204) <= input(28);
output(3, 205) <= input(29);
output(3, 206) <= input(30);
output(3, 207) <= input(31);
output(3, 208) <= input(16);
output(3, 209) <= input(17);
output(3, 210) <= input(18);
output(3, 211) <= input(19);
output(3, 212) <= input(20);
output(3, 213) <= input(21);
output(3, 214) <= input(22);
output(3, 215) <= input(23);
output(3, 216) <= input(24);
output(3, 217) <= input(25);
output(3, 218) <= input(26);
output(3, 219) <= input(27);
output(3, 220) <= input(28);
output(3, 221) <= input(29);
output(3, 222) <= input(30);
output(3, 223) <= input(31);
output(3, 224) <= input(1);
output(3, 225) <= input(2);
output(3, 226) <= input(3);
output(3, 227) <= input(4);
output(3, 228) <= input(5);
output(3, 229) <= input(6);
output(3, 230) <= input(7);
output(3, 231) <= input(8);
output(3, 232) <= input(9);
output(3, 233) <= input(10);
output(3, 234) <= input(11);
output(3, 235) <= input(12);
output(3, 236) <= input(13);
output(3, 237) <= input(14);
output(3, 238) <= input(15);
output(3, 239) <= input(32);
output(3, 240) <= input(17);
output(3, 241) <= input(18);
output(3, 242) <= input(19);
output(3, 243) <= input(20);
output(3, 244) <= input(21);
output(3, 245) <= input(22);
output(3, 246) <= input(23);
output(3, 247) <= input(24);
output(3, 248) <= input(25);
output(3, 249) <= input(26);
output(3, 250) <= input(27);
output(3, 251) <= input(28);
output(3, 252) <= input(29);
output(3, 253) <= input(30);
output(3, 254) <= input(31);
output(3, 255) <= input(33);
output(4, 0) <= input(53);
output(4, 1) <= input(51);
output(4, 2) <= input(49);
output(4, 3) <= input(46);
output(4, 4) <= input(47);
output(4, 5) <= input(16);
output(4, 6) <= input(17);
output(4, 7) <= input(18);
output(4, 8) <= input(19);
output(4, 9) <= input(20);
output(4, 10) <= input(21);
output(4, 11) <= input(22);
output(4, 12) <= input(23);
output(4, 13) <= input(24);
output(4, 14) <= input(25);
output(4, 15) <= input(26);
output(4, 16) <= input(54);
output(4, 17) <= input(52);
output(4, 18) <= input(50);
output(4, 19) <= input(48);
output(4, 20) <= input(0);
output(4, 21) <= input(1);
output(4, 22) <= input(2);
output(4, 23) <= input(3);
output(4, 24) <= input(4);
output(4, 25) <= input(5);
output(4, 26) <= input(6);
output(4, 27) <= input(7);
output(4, 28) <= input(8);
output(4, 29) <= input(9);
output(4, 30) <= input(10);
output(4, 31) <= input(11);
output(4, 32) <= input(54);
output(4, 33) <= input(52);
output(4, 34) <= input(50);
output(4, 35) <= input(48);
output(4, 36) <= input(0);
output(4, 37) <= input(1);
output(4, 38) <= input(2);
output(4, 39) <= input(3);
output(4, 40) <= input(4);
output(4, 41) <= input(5);
output(4, 42) <= input(6);
output(4, 43) <= input(7);
output(4, 44) <= input(8);
output(4, 45) <= input(9);
output(4, 46) <= input(10);
output(4, 47) <= input(11);
output(4, 48) <= input(51);
output(4, 49) <= input(49);
output(4, 50) <= input(46);
output(4, 51) <= input(47);
output(4, 52) <= input(16);
output(4, 53) <= input(17);
output(4, 54) <= input(18);
output(4, 55) <= input(19);
output(4, 56) <= input(20);
output(4, 57) <= input(21);
output(4, 58) <= input(22);
output(4, 59) <= input(23);
output(4, 60) <= input(24);
output(4, 61) <= input(25);
output(4, 62) <= input(26);
output(4, 63) <= input(27);
output(4, 64) <= input(51);
output(4, 65) <= input(49);
output(4, 66) <= input(46);
output(4, 67) <= input(47);
output(4, 68) <= input(16);
output(4, 69) <= input(17);
output(4, 70) <= input(18);
output(4, 71) <= input(19);
output(4, 72) <= input(20);
output(4, 73) <= input(21);
output(4, 74) <= input(22);
output(4, 75) <= input(23);
output(4, 76) <= input(24);
output(4, 77) <= input(25);
output(4, 78) <= input(26);
output(4, 79) <= input(27);
output(4, 80) <= input(52);
output(4, 81) <= input(50);
output(4, 82) <= input(48);
output(4, 83) <= input(0);
output(4, 84) <= input(1);
output(4, 85) <= input(2);
output(4, 86) <= input(3);
output(4, 87) <= input(4);
output(4, 88) <= input(5);
output(4, 89) <= input(6);
output(4, 90) <= input(7);
output(4, 91) <= input(8);
output(4, 92) <= input(9);
output(4, 93) <= input(10);
output(4, 94) <= input(11);
output(4, 95) <= input(12);
output(4, 96) <= input(52);
output(4, 97) <= input(50);
output(4, 98) <= input(48);
output(4, 99) <= input(0);
output(4, 100) <= input(1);
output(4, 101) <= input(2);
output(4, 102) <= input(3);
output(4, 103) <= input(4);
output(4, 104) <= input(5);
output(4, 105) <= input(6);
output(4, 106) <= input(7);
output(4, 107) <= input(8);
output(4, 108) <= input(9);
output(4, 109) <= input(10);
output(4, 110) <= input(11);
output(4, 111) <= input(12);
output(4, 112) <= input(49);
output(4, 113) <= input(46);
output(4, 114) <= input(47);
output(4, 115) <= input(16);
output(4, 116) <= input(17);
output(4, 117) <= input(18);
output(4, 118) <= input(19);
output(4, 119) <= input(20);
output(4, 120) <= input(21);
output(4, 121) <= input(22);
output(4, 122) <= input(23);
output(4, 123) <= input(24);
output(4, 124) <= input(25);
output(4, 125) <= input(26);
output(4, 126) <= input(27);
output(4, 127) <= input(28);
output(4, 128) <= input(49);
output(4, 129) <= input(46);
output(4, 130) <= input(47);
output(4, 131) <= input(16);
output(4, 132) <= input(17);
output(4, 133) <= input(18);
output(4, 134) <= input(19);
output(4, 135) <= input(20);
output(4, 136) <= input(21);
output(4, 137) <= input(22);
output(4, 138) <= input(23);
output(4, 139) <= input(24);
output(4, 140) <= input(25);
output(4, 141) <= input(26);
output(4, 142) <= input(27);
output(4, 143) <= input(28);
output(4, 144) <= input(50);
output(4, 145) <= input(48);
output(4, 146) <= input(0);
output(4, 147) <= input(1);
output(4, 148) <= input(2);
output(4, 149) <= input(3);
output(4, 150) <= input(4);
output(4, 151) <= input(5);
output(4, 152) <= input(6);
output(4, 153) <= input(7);
output(4, 154) <= input(8);
output(4, 155) <= input(9);
output(4, 156) <= input(10);
output(4, 157) <= input(11);
output(4, 158) <= input(12);
output(4, 159) <= input(13);
output(4, 160) <= input(50);
output(4, 161) <= input(48);
output(4, 162) <= input(0);
output(4, 163) <= input(1);
output(4, 164) <= input(2);
output(4, 165) <= input(3);
output(4, 166) <= input(4);
output(4, 167) <= input(5);
output(4, 168) <= input(6);
output(4, 169) <= input(7);
output(4, 170) <= input(8);
output(4, 171) <= input(9);
output(4, 172) <= input(10);
output(4, 173) <= input(11);
output(4, 174) <= input(12);
output(4, 175) <= input(13);
output(4, 176) <= input(46);
output(4, 177) <= input(47);
output(4, 178) <= input(16);
output(4, 179) <= input(17);
output(4, 180) <= input(18);
output(4, 181) <= input(19);
output(4, 182) <= input(20);
output(4, 183) <= input(21);
output(4, 184) <= input(22);
output(4, 185) <= input(23);
output(4, 186) <= input(24);
output(4, 187) <= input(25);
output(4, 188) <= input(26);
output(4, 189) <= input(27);
output(4, 190) <= input(28);
output(4, 191) <= input(29);
output(4, 192) <= input(46);
output(4, 193) <= input(47);
output(4, 194) <= input(16);
output(4, 195) <= input(17);
output(4, 196) <= input(18);
output(4, 197) <= input(19);
output(4, 198) <= input(20);
output(4, 199) <= input(21);
output(4, 200) <= input(22);
output(4, 201) <= input(23);
output(4, 202) <= input(24);
output(4, 203) <= input(25);
output(4, 204) <= input(26);
output(4, 205) <= input(27);
output(4, 206) <= input(28);
output(4, 207) <= input(29);
output(4, 208) <= input(48);
output(4, 209) <= input(0);
output(4, 210) <= input(1);
output(4, 211) <= input(2);
output(4, 212) <= input(3);
output(4, 213) <= input(4);
output(4, 214) <= input(5);
output(4, 215) <= input(6);
output(4, 216) <= input(7);
output(4, 217) <= input(8);
output(4, 218) <= input(9);
output(4, 219) <= input(10);
output(4, 220) <= input(11);
output(4, 221) <= input(12);
output(4, 222) <= input(13);
output(4, 223) <= input(14);
output(4, 224) <= input(48);
output(4, 225) <= input(0);
output(4, 226) <= input(1);
output(4, 227) <= input(2);
output(4, 228) <= input(3);
output(4, 229) <= input(4);
output(4, 230) <= input(5);
output(4, 231) <= input(6);
output(4, 232) <= input(7);
output(4, 233) <= input(8);
output(4, 234) <= input(9);
output(4, 235) <= input(10);
output(4, 236) <= input(11);
output(4, 237) <= input(12);
output(4, 238) <= input(13);
output(4, 239) <= input(14);
output(4, 240) <= input(47);
output(4, 241) <= input(16);
output(4, 242) <= input(17);
output(4, 243) <= input(18);
output(4, 244) <= input(19);
output(4, 245) <= input(20);
output(4, 246) <= input(21);
output(4, 247) <= input(22);
output(4, 248) <= input(23);
output(4, 249) <= input(24);
output(4, 250) <= input(25);
output(4, 251) <= input(26);
output(4, 252) <= input(27);
output(4, 253) <= input(28);
output(4, 254) <= input(29);
output(4, 255) <= input(30);
output(5, 0) <= input(55);
output(5, 1) <= input(53);
output(5, 2) <= input(51);
output(5, 3) <= input(49);
output(5, 4) <= input(46);
output(5, 5) <= input(47);
output(5, 6) <= input(16);
output(5, 7) <= input(17);
output(5, 8) <= input(18);
output(5, 9) <= input(19);
output(5, 10) <= input(20);
output(5, 11) <= input(21);
output(5, 12) <= input(22);
output(5, 13) <= input(23);
output(5, 14) <= input(24);
output(5, 15) <= input(25);
output(5, 16) <= input(55);
output(5, 17) <= input(53);
output(5, 18) <= input(51);
output(5, 19) <= input(49);
output(5, 20) <= input(46);
output(5, 21) <= input(47);
output(5, 22) <= input(16);
output(5, 23) <= input(17);
output(5, 24) <= input(18);
output(5, 25) <= input(19);
output(5, 26) <= input(20);
output(5, 27) <= input(21);
output(5, 28) <= input(22);
output(5, 29) <= input(23);
output(5, 30) <= input(24);
output(5, 31) <= input(25);
output(5, 32) <= input(56);
output(5, 33) <= input(54);
output(5, 34) <= input(52);
output(5, 35) <= input(50);
output(5, 36) <= input(48);
output(5, 37) <= input(0);
output(5, 38) <= input(1);
output(5, 39) <= input(2);
output(5, 40) <= input(3);
output(5, 41) <= input(4);
output(5, 42) <= input(5);
output(5, 43) <= input(6);
output(5, 44) <= input(7);
output(5, 45) <= input(8);
output(5, 46) <= input(9);
output(5, 47) <= input(10);
output(5, 48) <= input(56);
output(5, 49) <= input(54);
output(5, 50) <= input(52);
output(5, 51) <= input(50);
output(5, 52) <= input(48);
output(5, 53) <= input(0);
output(5, 54) <= input(1);
output(5, 55) <= input(2);
output(5, 56) <= input(3);
output(5, 57) <= input(4);
output(5, 58) <= input(5);
output(5, 59) <= input(6);
output(5, 60) <= input(7);
output(5, 61) <= input(8);
output(5, 62) <= input(9);
output(5, 63) <= input(10);
output(5, 64) <= input(56);
output(5, 65) <= input(54);
output(5, 66) <= input(52);
output(5, 67) <= input(50);
output(5, 68) <= input(48);
output(5, 69) <= input(0);
output(5, 70) <= input(1);
output(5, 71) <= input(2);
output(5, 72) <= input(3);
output(5, 73) <= input(4);
output(5, 74) <= input(5);
output(5, 75) <= input(6);
output(5, 76) <= input(7);
output(5, 77) <= input(8);
output(5, 78) <= input(9);
output(5, 79) <= input(10);
output(5, 80) <= input(53);
output(5, 81) <= input(51);
output(5, 82) <= input(49);
output(5, 83) <= input(46);
output(5, 84) <= input(47);
output(5, 85) <= input(16);
output(5, 86) <= input(17);
output(5, 87) <= input(18);
output(5, 88) <= input(19);
output(5, 89) <= input(20);
output(5, 90) <= input(21);
output(5, 91) <= input(22);
output(5, 92) <= input(23);
output(5, 93) <= input(24);
output(5, 94) <= input(25);
output(5, 95) <= input(26);
output(5, 96) <= input(53);
output(5, 97) <= input(51);
output(5, 98) <= input(49);
output(5, 99) <= input(46);
output(5, 100) <= input(47);
output(5, 101) <= input(16);
output(5, 102) <= input(17);
output(5, 103) <= input(18);
output(5, 104) <= input(19);
output(5, 105) <= input(20);
output(5, 106) <= input(21);
output(5, 107) <= input(22);
output(5, 108) <= input(23);
output(5, 109) <= input(24);
output(5, 110) <= input(25);
output(5, 111) <= input(26);
output(5, 112) <= input(54);
output(5, 113) <= input(52);
output(5, 114) <= input(50);
output(5, 115) <= input(48);
output(5, 116) <= input(0);
output(5, 117) <= input(1);
output(5, 118) <= input(2);
output(5, 119) <= input(3);
output(5, 120) <= input(4);
output(5, 121) <= input(5);
output(5, 122) <= input(6);
output(5, 123) <= input(7);
output(5, 124) <= input(8);
output(5, 125) <= input(9);
output(5, 126) <= input(10);
output(5, 127) <= input(11);
output(5, 128) <= input(54);
output(5, 129) <= input(52);
output(5, 130) <= input(50);
output(5, 131) <= input(48);
output(5, 132) <= input(0);
output(5, 133) <= input(1);
output(5, 134) <= input(2);
output(5, 135) <= input(3);
output(5, 136) <= input(4);
output(5, 137) <= input(5);
output(5, 138) <= input(6);
output(5, 139) <= input(7);
output(5, 140) <= input(8);
output(5, 141) <= input(9);
output(5, 142) <= input(10);
output(5, 143) <= input(11);
output(5, 144) <= input(54);
output(5, 145) <= input(52);
output(5, 146) <= input(50);
output(5, 147) <= input(48);
output(5, 148) <= input(0);
output(5, 149) <= input(1);
output(5, 150) <= input(2);
output(5, 151) <= input(3);
output(5, 152) <= input(4);
output(5, 153) <= input(5);
output(5, 154) <= input(6);
output(5, 155) <= input(7);
output(5, 156) <= input(8);
output(5, 157) <= input(9);
output(5, 158) <= input(10);
output(5, 159) <= input(11);
output(5, 160) <= input(51);
output(5, 161) <= input(49);
output(5, 162) <= input(46);
output(5, 163) <= input(47);
output(5, 164) <= input(16);
output(5, 165) <= input(17);
output(5, 166) <= input(18);
output(5, 167) <= input(19);
output(5, 168) <= input(20);
output(5, 169) <= input(21);
output(5, 170) <= input(22);
output(5, 171) <= input(23);
output(5, 172) <= input(24);
output(5, 173) <= input(25);
output(5, 174) <= input(26);
output(5, 175) <= input(27);
output(5, 176) <= input(51);
output(5, 177) <= input(49);
output(5, 178) <= input(46);
output(5, 179) <= input(47);
output(5, 180) <= input(16);
output(5, 181) <= input(17);
output(5, 182) <= input(18);
output(5, 183) <= input(19);
output(5, 184) <= input(20);
output(5, 185) <= input(21);
output(5, 186) <= input(22);
output(5, 187) <= input(23);
output(5, 188) <= input(24);
output(5, 189) <= input(25);
output(5, 190) <= input(26);
output(5, 191) <= input(27);
output(5, 192) <= input(51);
output(5, 193) <= input(49);
output(5, 194) <= input(46);
output(5, 195) <= input(47);
output(5, 196) <= input(16);
output(5, 197) <= input(17);
output(5, 198) <= input(18);
output(5, 199) <= input(19);
output(5, 200) <= input(20);
output(5, 201) <= input(21);
output(5, 202) <= input(22);
output(5, 203) <= input(23);
output(5, 204) <= input(24);
output(5, 205) <= input(25);
output(5, 206) <= input(26);
output(5, 207) <= input(27);
output(5, 208) <= input(52);
output(5, 209) <= input(50);
output(5, 210) <= input(48);
output(5, 211) <= input(0);
output(5, 212) <= input(1);
output(5, 213) <= input(2);
output(5, 214) <= input(3);
output(5, 215) <= input(4);
output(5, 216) <= input(5);
output(5, 217) <= input(6);
output(5, 218) <= input(7);
output(5, 219) <= input(8);
output(5, 220) <= input(9);
output(5, 221) <= input(10);
output(5, 222) <= input(11);
output(5, 223) <= input(12);
output(5, 224) <= input(52);
output(5, 225) <= input(50);
output(5, 226) <= input(48);
output(5, 227) <= input(0);
output(5, 228) <= input(1);
output(5, 229) <= input(2);
output(5, 230) <= input(3);
output(5, 231) <= input(4);
output(5, 232) <= input(5);
output(5, 233) <= input(6);
output(5, 234) <= input(7);
output(5, 235) <= input(8);
output(5, 236) <= input(9);
output(5, 237) <= input(10);
output(5, 238) <= input(11);
output(5, 239) <= input(12);
output(5, 240) <= input(49);
output(5, 241) <= input(46);
output(5, 242) <= input(47);
output(5, 243) <= input(16);
output(5, 244) <= input(17);
output(5, 245) <= input(18);
output(5, 246) <= input(19);
output(5, 247) <= input(20);
output(5, 248) <= input(21);
output(5, 249) <= input(22);
output(5, 250) <= input(23);
output(5, 251) <= input(24);
output(5, 252) <= input(25);
output(5, 253) <= input(26);
output(5, 254) <= input(27);
output(5, 255) <= input(28);
when "0010" =>
output(0, 0) <= input(0);
output(0, 1) <= input(1);
output(0, 2) <= input(2);
output(0, 3) <= input(3);
output(0, 4) <= input(4);
output(0, 5) <= input(5);
output(0, 6) <= input(6);
output(0, 7) <= input(7);
output(0, 8) <= input(8);
output(0, 9) <= input(9);
output(0, 10) <= input(10);
output(0, 11) <= input(11);
output(0, 12) <= input(12);
output(0, 13) <= input(13);
output(0, 14) <= input(14);
output(0, 15) <= input(15);
output(0, 16) <= input(0);
output(0, 17) <= input(1);
output(0, 18) <= input(2);
output(0, 19) <= input(3);
output(0, 20) <= input(4);
output(0, 21) <= input(5);
output(0, 22) <= input(6);
output(0, 23) <= input(7);
output(0, 24) <= input(8);
output(0, 25) <= input(9);
output(0, 26) <= input(10);
output(0, 27) <= input(11);
output(0, 28) <= input(12);
output(0, 29) <= input(13);
output(0, 30) <= input(14);
output(0, 31) <= input(15);
output(0, 32) <= input(0);
output(0, 33) <= input(1);
output(0, 34) <= input(2);
output(0, 35) <= input(3);
output(0, 36) <= input(4);
output(0, 37) <= input(5);
output(0, 38) <= input(6);
output(0, 39) <= input(7);
output(0, 40) <= input(8);
output(0, 41) <= input(9);
output(0, 42) <= input(10);
output(0, 43) <= input(11);
output(0, 44) <= input(12);
output(0, 45) <= input(13);
output(0, 46) <= input(14);
output(0, 47) <= input(15);
output(0, 48) <= input(16);
output(0, 49) <= input(17);
output(0, 50) <= input(18);
output(0, 51) <= input(19);
output(0, 52) <= input(20);
output(0, 53) <= input(21);
output(0, 54) <= input(22);
output(0, 55) <= input(23);
output(0, 56) <= input(24);
output(0, 57) <= input(25);
output(0, 58) <= input(26);
output(0, 59) <= input(27);
output(0, 60) <= input(28);
output(0, 61) <= input(29);
output(0, 62) <= input(30);
output(0, 63) <= input(31);
output(0, 64) <= input(16);
output(0, 65) <= input(17);
output(0, 66) <= input(18);
output(0, 67) <= input(19);
output(0, 68) <= input(20);
output(0, 69) <= input(21);
output(0, 70) <= input(22);
output(0, 71) <= input(23);
output(0, 72) <= input(24);
output(0, 73) <= input(25);
output(0, 74) <= input(26);
output(0, 75) <= input(27);
output(0, 76) <= input(28);
output(0, 77) <= input(29);
output(0, 78) <= input(30);
output(0, 79) <= input(31);
output(0, 80) <= input(16);
output(0, 81) <= input(17);
output(0, 82) <= input(18);
output(0, 83) <= input(19);
output(0, 84) <= input(20);
output(0, 85) <= input(21);
output(0, 86) <= input(22);
output(0, 87) <= input(23);
output(0, 88) <= input(24);
output(0, 89) <= input(25);
output(0, 90) <= input(26);
output(0, 91) <= input(27);
output(0, 92) <= input(28);
output(0, 93) <= input(29);
output(0, 94) <= input(30);
output(0, 95) <= input(31);
output(0, 96) <= input(16);
output(0, 97) <= input(17);
output(0, 98) <= input(18);
output(0, 99) <= input(19);
output(0, 100) <= input(20);
output(0, 101) <= input(21);
output(0, 102) <= input(22);
output(0, 103) <= input(23);
output(0, 104) <= input(24);
output(0, 105) <= input(25);
output(0, 106) <= input(26);
output(0, 107) <= input(27);
output(0, 108) <= input(28);
output(0, 109) <= input(29);
output(0, 110) <= input(30);
output(0, 111) <= input(31);
output(0, 112) <= input(1);
output(0, 113) <= input(2);
output(0, 114) <= input(3);
output(0, 115) <= input(4);
output(0, 116) <= input(5);
output(0, 117) <= input(6);
output(0, 118) <= input(7);
output(0, 119) <= input(8);
output(0, 120) <= input(9);
output(0, 121) <= input(10);
output(0, 122) <= input(11);
output(0, 123) <= input(12);
output(0, 124) <= input(13);
output(0, 125) <= input(14);
output(0, 126) <= input(15);
output(0, 127) <= input(32);
output(0, 128) <= input(1);
output(0, 129) <= input(2);
output(0, 130) <= input(3);
output(0, 131) <= input(4);
output(0, 132) <= input(5);
output(0, 133) <= input(6);
output(0, 134) <= input(7);
output(0, 135) <= input(8);
output(0, 136) <= input(9);
output(0, 137) <= input(10);
output(0, 138) <= input(11);
output(0, 139) <= input(12);
output(0, 140) <= input(13);
output(0, 141) <= input(14);
output(0, 142) <= input(15);
output(0, 143) <= input(32);
output(0, 144) <= input(1);
output(0, 145) <= input(2);
output(0, 146) <= input(3);
output(0, 147) <= input(4);
output(0, 148) <= input(5);
output(0, 149) <= input(6);
output(0, 150) <= input(7);
output(0, 151) <= input(8);
output(0, 152) <= input(9);
output(0, 153) <= input(10);
output(0, 154) <= input(11);
output(0, 155) <= input(12);
output(0, 156) <= input(13);
output(0, 157) <= input(14);
output(0, 158) <= input(15);
output(0, 159) <= input(32);
output(0, 160) <= input(1);
output(0, 161) <= input(2);
output(0, 162) <= input(3);
output(0, 163) <= input(4);
output(0, 164) <= input(5);
output(0, 165) <= input(6);
output(0, 166) <= input(7);
output(0, 167) <= input(8);
output(0, 168) <= input(9);
output(0, 169) <= input(10);
output(0, 170) <= input(11);
output(0, 171) <= input(12);
output(0, 172) <= input(13);
output(0, 173) <= input(14);
output(0, 174) <= input(15);
output(0, 175) <= input(32);
output(0, 176) <= input(17);
output(0, 177) <= input(18);
output(0, 178) <= input(19);
output(0, 179) <= input(20);
output(0, 180) <= input(21);
output(0, 181) <= input(22);
output(0, 182) <= input(23);
output(0, 183) <= input(24);
output(0, 184) <= input(25);
output(0, 185) <= input(26);
output(0, 186) <= input(27);
output(0, 187) <= input(28);
output(0, 188) <= input(29);
output(0, 189) <= input(30);
output(0, 190) <= input(31);
output(0, 191) <= input(33);
output(0, 192) <= input(17);
output(0, 193) <= input(18);
output(0, 194) <= input(19);
output(0, 195) <= input(20);
output(0, 196) <= input(21);
output(0, 197) <= input(22);
output(0, 198) <= input(23);
output(0, 199) <= input(24);
output(0, 200) <= input(25);
output(0, 201) <= input(26);
output(0, 202) <= input(27);
output(0, 203) <= input(28);
output(0, 204) <= input(29);
output(0, 205) <= input(30);
output(0, 206) <= input(31);
output(0, 207) <= input(33);
output(0, 208) <= input(17);
output(0, 209) <= input(18);
output(0, 210) <= input(19);
output(0, 211) <= input(20);
output(0, 212) <= input(21);
output(0, 213) <= input(22);
output(0, 214) <= input(23);
output(0, 215) <= input(24);
output(0, 216) <= input(25);
output(0, 217) <= input(26);
output(0, 218) <= input(27);
output(0, 219) <= input(28);
output(0, 220) <= input(29);
output(0, 221) <= input(30);
output(0, 222) <= input(31);
output(0, 223) <= input(33);
output(0, 224) <= input(17);
output(0, 225) <= input(18);
output(0, 226) <= input(19);
output(0, 227) <= input(20);
output(0, 228) <= input(21);
output(0, 229) <= input(22);
output(0, 230) <= input(23);
output(0, 231) <= input(24);
output(0, 232) <= input(25);
output(0, 233) <= input(26);
output(0, 234) <= input(27);
output(0, 235) <= input(28);
output(0, 236) <= input(29);
output(0, 237) <= input(30);
output(0, 238) <= input(31);
output(0, 239) <= input(33);
output(0, 240) <= input(2);
output(0, 241) <= input(3);
output(0, 242) <= input(4);
output(0, 243) <= input(5);
output(0, 244) <= input(6);
output(0, 245) <= input(7);
output(0, 246) <= input(8);
output(0, 247) <= input(9);
output(0, 248) <= input(10);
output(0, 249) <= input(11);
output(0, 250) <= input(12);
output(0, 251) <= input(13);
output(0, 252) <= input(14);
output(0, 253) <= input(15);
output(0, 254) <= input(32);
output(0, 255) <= input(34);
output(1, 0) <= input(35);
output(1, 1) <= input(16);
output(1, 2) <= input(17);
output(1, 3) <= input(18);
output(1, 4) <= input(19);
output(1, 5) <= input(20);
output(1, 6) <= input(21);
output(1, 7) <= input(22);
output(1, 8) <= input(23);
output(1, 9) <= input(24);
output(1, 10) <= input(25);
output(1, 11) <= input(26);
output(1, 12) <= input(27);
output(1, 13) <= input(28);
output(1, 14) <= input(29);
output(1, 15) <= input(30);
output(1, 16) <= input(35);
output(1, 17) <= input(16);
output(1, 18) <= input(17);
output(1, 19) <= input(18);
output(1, 20) <= input(19);
output(1, 21) <= input(20);
output(1, 22) <= input(21);
output(1, 23) <= input(22);
output(1, 24) <= input(23);
output(1, 25) <= input(24);
output(1, 26) <= input(25);
output(1, 27) <= input(26);
output(1, 28) <= input(27);
output(1, 29) <= input(28);
output(1, 30) <= input(29);
output(1, 31) <= input(30);
output(1, 32) <= input(35);
output(1, 33) <= input(16);
output(1, 34) <= input(17);
output(1, 35) <= input(18);
output(1, 36) <= input(19);
output(1, 37) <= input(20);
output(1, 38) <= input(21);
output(1, 39) <= input(22);
output(1, 40) <= input(23);
output(1, 41) <= input(24);
output(1, 42) <= input(25);
output(1, 43) <= input(26);
output(1, 44) <= input(27);
output(1, 45) <= input(28);
output(1, 46) <= input(29);
output(1, 47) <= input(30);
output(1, 48) <= input(35);
output(1, 49) <= input(16);
output(1, 50) <= input(17);
output(1, 51) <= input(18);
output(1, 52) <= input(19);
output(1, 53) <= input(20);
output(1, 54) <= input(21);
output(1, 55) <= input(22);
output(1, 56) <= input(23);
output(1, 57) <= input(24);
output(1, 58) <= input(25);
output(1, 59) <= input(26);
output(1, 60) <= input(27);
output(1, 61) <= input(28);
output(1, 62) <= input(29);
output(1, 63) <= input(30);
output(1, 64) <= input(35);
output(1, 65) <= input(16);
output(1, 66) <= input(17);
output(1, 67) <= input(18);
output(1, 68) <= input(19);
output(1, 69) <= input(20);
output(1, 70) <= input(21);
output(1, 71) <= input(22);
output(1, 72) <= input(23);
output(1, 73) <= input(24);
output(1, 74) <= input(25);
output(1, 75) <= input(26);
output(1, 76) <= input(27);
output(1, 77) <= input(28);
output(1, 78) <= input(29);
output(1, 79) <= input(30);
output(1, 80) <= input(0);
output(1, 81) <= input(1);
output(1, 82) <= input(2);
output(1, 83) <= input(3);
output(1, 84) <= input(4);
output(1, 85) <= input(5);
output(1, 86) <= input(6);
output(1, 87) <= input(7);
output(1, 88) <= input(8);
output(1, 89) <= input(9);
output(1, 90) <= input(10);
output(1, 91) <= input(11);
output(1, 92) <= input(12);
output(1, 93) <= input(13);
output(1, 94) <= input(14);
output(1, 95) <= input(15);
output(1, 96) <= input(0);
output(1, 97) <= input(1);
output(1, 98) <= input(2);
output(1, 99) <= input(3);
output(1, 100) <= input(4);
output(1, 101) <= input(5);
output(1, 102) <= input(6);
output(1, 103) <= input(7);
output(1, 104) <= input(8);
output(1, 105) <= input(9);
output(1, 106) <= input(10);
output(1, 107) <= input(11);
output(1, 108) <= input(12);
output(1, 109) <= input(13);
output(1, 110) <= input(14);
output(1, 111) <= input(15);
output(1, 112) <= input(0);
output(1, 113) <= input(1);
output(1, 114) <= input(2);
output(1, 115) <= input(3);
output(1, 116) <= input(4);
output(1, 117) <= input(5);
output(1, 118) <= input(6);
output(1, 119) <= input(7);
output(1, 120) <= input(8);
output(1, 121) <= input(9);
output(1, 122) <= input(10);
output(1, 123) <= input(11);
output(1, 124) <= input(12);
output(1, 125) <= input(13);
output(1, 126) <= input(14);
output(1, 127) <= input(15);
output(1, 128) <= input(0);
output(1, 129) <= input(1);
output(1, 130) <= input(2);
output(1, 131) <= input(3);
output(1, 132) <= input(4);
output(1, 133) <= input(5);
output(1, 134) <= input(6);
output(1, 135) <= input(7);
output(1, 136) <= input(8);
output(1, 137) <= input(9);
output(1, 138) <= input(10);
output(1, 139) <= input(11);
output(1, 140) <= input(12);
output(1, 141) <= input(13);
output(1, 142) <= input(14);
output(1, 143) <= input(15);
output(1, 144) <= input(0);
output(1, 145) <= input(1);
output(1, 146) <= input(2);
output(1, 147) <= input(3);
output(1, 148) <= input(4);
output(1, 149) <= input(5);
output(1, 150) <= input(6);
output(1, 151) <= input(7);
output(1, 152) <= input(8);
output(1, 153) <= input(9);
output(1, 154) <= input(10);
output(1, 155) <= input(11);
output(1, 156) <= input(12);
output(1, 157) <= input(13);
output(1, 158) <= input(14);
output(1, 159) <= input(15);
output(1, 160) <= input(16);
output(1, 161) <= input(17);
output(1, 162) <= input(18);
output(1, 163) <= input(19);
output(1, 164) <= input(20);
output(1, 165) <= input(21);
output(1, 166) <= input(22);
output(1, 167) <= input(23);
output(1, 168) <= input(24);
output(1, 169) <= input(25);
output(1, 170) <= input(26);
output(1, 171) <= input(27);
output(1, 172) <= input(28);
output(1, 173) <= input(29);
output(1, 174) <= input(30);
output(1, 175) <= input(31);
output(1, 176) <= input(16);
output(1, 177) <= input(17);
output(1, 178) <= input(18);
output(1, 179) <= input(19);
output(1, 180) <= input(20);
output(1, 181) <= input(21);
output(1, 182) <= input(22);
output(1, 183) <= input(23);
output(1, 184) <= input(24);
output(1, 185) <= input(25);
output(1, 186) <= input(26);
output(1, 187) <= input(27);
output(1, 188) <= input(28);
output(1, 189) <= input(29);
output(1, 190) <= input(30);
output(1, 191) <= input(31);
output(1, 192) <= input(16);
output(1, 193) <= input(17);
output(1, 194) <= input(18);
output(1, 195) <= input(19);
output(1, 196) <= input(20);
output(1, 197) <= input(21);
output(1, 198) <= input(22);
output(1, 199) <= input(23);
output(1, 200) <= input(24);
output(1, 201) <= input(25);
output(1, 202) <= input(26);
output(1, 203) <= input(27);
output(1, 204) <= input(28);
output(1, 205) <= input(29);
output(1, 206) <= input(30);
output(1, 207) <= input(31);
output(1, 208) <= input(16);
output(1, 209) <= input(17);
output(1, 210) <= input(18);
output(1, 211) <= input(19);
output(1, 212) <= input(20);
output(1, 213) <= input(21);
output(1, 214) <= input(22);
output(1, 215) <= input(23);
output(1, 216) <= input(24);
output(1, 217) <= input(25);
output(1, 218) <= input(26);
output(1, 219) <= input(27);
output(1, 220) <= input(28);
output(1, 221) <= input(29);
output(1, 222) <= input(30);
output(1, 223) <= input(31);
output(1, 224) <= input(16);
output(1, 225) <= input(17);
output(1, 226) <= input(18);
output(1, 227) <= input(19);
output(1, 228) <= input(20);
output(1, 229) <= input(21);
output(1, 230) <= input(22);
output(1, 231) <= input(23);
output(1, 232) <= input(24);
output(1, 233) <= input(25);
output(1, 234) <= input(26);
output(1, 235) <= input(27);
output(1, 236) <= input(28);
output(1, 237) <= input(29);
output(1, 238) <= input(30);
output(1, 239) <= input(31);
output(1, 240) <= input(1);
output(1, 241) <= input(2);
output(1, 242) <= input(3);
output(1, 243) <= input(4);
output(1, 244) <= input(5);
output(1, 245) <= input(6);
output(1, 246) <= input(7);
output(1, 247) <= input(8);
output(1, 248) <= input(9);
output(1, 249) <= input(10);
output(1, 250) <= input(11);
output(1, 251) <= input(12);
output(1, 252) <= input(13);
output(1, 253) <= input(14);
output(1, 254) <= input(15);
output(1, 255) <= input(32);
output(2, 0) <= input(36);
output(2, 1) <= input(0);
output(2, 2) <= input(1);
output(2, 3) <= input(2);
output(2, 4) <= input(3);
output(2, 5) <= input(4);
output(2, 6) <= input(5);
output(2, 7) <= input(6);
output(2, 8) <= input(7);
output(2, 9) <= input(8);
output(2, 10) <= input(9);
output(2, 11) <= input(10);
output(2, 12) <= input(11);
output(2, 13) <= input(12);
output(2, 14) <= input(13);
output(2, 15) <= input(14);
output(2, 16) <= input(36);
output(2, 17) <= input(0);
output(2, 18) <= input(1);
output(2, 19) <= input(2);
output(2, 20) <= input(3);
output(2, 21) <= input(4);
output(2, 22) <= input(5);
output(2, 23) <= input(6);
output(2, 24) <= input(7);
output(2, 25) <= input(8);
output(2, 26) <= input(9);
output(2, 27) <= input(10);
output(2, 28) <= input(11);
output(2, 29) <= input(12);
output(2, 30) <= input(13);
output(2, 31) <= input(14);
output(2, 32) <= input(36);
output(2, 33) <= input(0);
output(2, 34) <= input(1);
output(2, 35) <= input(2);
output(2, 36) <= input(3);
output(2, 37) <= input(4);
output(2, 38) <= input(5);
output(2, 39) <= input(6);
output(2, 40) <= input(7);
output(2, 41) <= input(8);
output(2, 42) <= input(9);
output(2, 43) <= input(10);
output(2, 44) <= input(11);
output(2, 45) <= input(12);
output(2, 46) <= input(13);
output(2, 47) <= input(14);
output(2, 48) <= input(36);
output(2, 49) <= input(0);
output(2, 50) <= input(1);
output(2, 51) <= input(2);
output(2, 52) <= input(3);
output(2, 53) <= input(4);
output(2, 54) <= input(5);
output(2, 55) <= input(6);
output(2, 56) <= input(7);
output(2, 57) <= input(8);
output(2, 58) <= input(9);
output(2, 59) <= input(10);
output(2, 60) <= input(11);
output(2, 61) <= input(12);
output(2, 62) <= input(13);
output(2, 63) <= input(14);
output(2, 64) <= input(36);
output(2, 65) <= input(0);
output(2, 66) <= input(1);
output(2, 67) <= input(2);
output(2, 68) <= input(3);
output(2, 69) <= input(4);
output(2, 70) <= input(5);
output(2, 71) <= input(6);
output(2, 72) <= input(7);
output(2, 73) <= input(8);
output(2, 74) <= input(9);
output(2, 75) <= input(10);
output(2, 76) <= input(11);
output(2, 77) <= input(12);
output(2, 78) <= input(13);
output(2, 79) <= input(14);
output(2, 80) <= input(36);
output(2, 81) <= input(0);
output(2, 82) <= input(1);
output(2, 83) <= input(2);
output(2, 84) <= input(3);
output(2, 85) <= input(4);
output(2, 86) <= input(5);
output(2, 87) <= input(6);
output(2, 88) <= input(7);
output(2, 89) <= input(8);
output(2, 90) <= input(9);
output(2, 91) <= input(10);
output(2, 92) <= input(11);
output(2, 93) <= input(12);
output(2, 94) <= input(13);
output(2, 95) <= input(14);
output(2, 96) <= input(36);
output(2, 97) <= input(0);
output(2, 98) <= input(1);
output(2, 99) <= input(2);
output(2, 100) <= input(3);
output(2, 101) <= input(4);
output(2, 102) <= input(5);
output(2, 103) <= input(6);
output(2, 104) <= input(7);
output(2, 105) <= input(8);
output(2, 106) <= input(9);
output(2, 107) <= input(10);
output(2, 108) <= input(11);
output(2, 109) <= input(12);
output(2, 110) <= input(13);
output(2, 111) <= input(14);
output(2, 112) <= input(35);
output(2, 113) <= input(16);
output(2, 114) <= input(17);
output(2, 115) <= input(18);
output(2, 116) <= input(19);
output(2, 117) <= input(20);
output(2, 118) <= input(21);
output(2, 119) <= input(22);
output(2, 120) <= input(23);
output(2, 121) <= input(24);
output(2, 122) <= input(25);
output(2, 123) <= input(26);
output(2, 124) <= input(27);
output(2, 125) <= input(28);
output(2, 126) <= input(29);
output(2, 127) <= input(30);
output(2, 128) <= input(35);
output(2, 129) <= input(16);
output(2, 130) <= input(17);
output(2, 131) <= input(18);
output(2, 132) <= input(19);
output(2, 133) <= input(20);
output(2, 134) <= input(21);
output(2, 135) <= input(22);
output(2, 136) <= input(23);
output(2, 137) <= input(24);
output(2, 138) <= input(25);
output(2, 139) <= input(26);
output(2, 140) <= input(27);
output(2, 141) <= input(28);
output(2, 142) <= input(29);
output(2, 143) <= input(30);
output(2, 144) <= input(35);
output(2, 145) <= input(16);
output(2, 146) <= input(17);
output(2, 147) <= input(18);
output(2, 148) <= input(19);
output(2, 149) <= input(20);
output(2, 150) <= input(21);
output(2, 151) <= input(22);
output(2, 152) <= input(23);
output(2, 153) <= input(24);
output(2, 154) <= input(25);
output(2, 155) <= input(26);
output(2, 156) <= input(27);
output(2, 157) <= input(28);
output(2, 158) <= input(29);
output(2, 159) <= input(30);
output(2, 160) <= input(35);
output(2, 161) <= input(16);
output(2, 162) <= input(17);
output(2, 163) <= input(18);
output(2, 164) <= input(19);
output(2, 165) <= input(20);
output(2, 166) <= input(21);
output(2, 167) <= input(22);
output(2, 168) <= input(23);
output(2, 169) <= input(24);
output(2, 170) <= input(25);
output(2, 171) <= input(26);
output(2, 172) <= input(27);
output(2, 173) <= input(28);
output(2, 174) <= input(29);
output(2, 175) <= input(30);
output(2, 176) <= input(35);
output(2, 177) <= input(16);
output(2, 178) <= input(17);
output(2, 179) <= input(18);
output(2, 180) <= input(19);
output(2, 181) <= input(20);
output(2, 182) <= input(21);
output(2, 183) <= input(22);
output(2, 184) <= input(23);
output(2, 185) <= input(24);
output(2, 186) <= input(25);
output(2, 187) <= input(26);
output(2, 188) <= input(27);
output(2, 189) <= input(28);
output(2, 190) <= input(29);
output(2, 191) <= input(30);
output(2, 192) <= input(35);
output(2, 193) <= input(16);
output(2, 194) <= input(17);
output(2, 195) <= input(18);
output(2, 196) <= input(19);
output(2, 197) <= input(20);
output(2, 198) <= input(21);
output(2, 199) <= input(22);
output(2, 200) <= input(23);
output(2, 201) <= input(24);
output(2, 202) <= input(25);
output(2, 203) <= input(26);
output(2, 204) <= input(27);
output(2, 205) <= input(28);
output(2, 206) <= input(29);
output(2, 207) <= input(30);
output(2, 208) <= input(35);
output(2, 209) <= input(16);
output(2, 210) <= input(17);
output(2, 211) <= input(18);
output(2, 212) <= input(19);
output(2, 213) <= input(20);
output(2, 214) <= input(21);
output(2, 215) <= input(22);
output(2, 216) <= input(23);
output(2, 217) <= input(24);
output(2, 218) <= input(25);
output(2, 219) <= input(26);
output(2, 220) <= input(27);
output(2, 221) <= input(28);
output(2, 222) <= input(29);
output(2, 223) <= input(30);
output(2, 224) <= input(35);
output(2, 225) <= input(16);
output(2, 226) <= input(17);
output(2, 227) <= input(18);
output(2, 228) <= input(19);
output(2, 229) <= input(20);
output(2, 230) <= input(21);
output(2, 231) <= input(22);
output(2, 232) <= input(23);
output(2, 233) <= input(24);
output(2, 234) <= input(25);
output(2, 235) <= input(26);
output(2, 236) <= input(27);
output(2, 237) <= input(28);
output(2, 238) <= input(29);
output(2, 239) <= input(30);
output(2, 240) <= input(0);
output(2, 241) <= input(1);
output(2, 242) <= input(2);
output(2, 243) <= input(3);
output(2, 244) <= input(4);
output(2, 245) <= input(5);
output(2, 246) <= input(6);
output(2, 247) <= input(7);
output(2, 248) <= input(8);
output(2, 249) <= input(9);
output(2, 250) <= input(10);
output(2, 251) <= input(11);
output(2, 252) <= input(12);
output(2, 253) <= input(13);
output(2, 254) <= input(14);
output(2, 255) <= input(15);
output(3, 0) <= input(37);
output(3, 1) <= input(35);
output(3, 2) <= input(16);
output(3, 3) <= input(17);
output(3, 4) <= input(18);
output(3, 5) <= input(19);
output(3, 6) <= input(20);
output(3, 7) <= input(21);
output(3, 8) <= input(22);
output(3, 9) <= input(23);
output(3, 10) <= input(24);
output(3, 11) <= input(25);
output(3, 12) <= input(26);
output(3, 13) <= input(27);
output(3, 14) <= input(28);
output(3, 15) <= input(29);
output(3, 16) <= input(37);
output(3, 17) <= input(35);
output(3, 18) <= input(16);
output(3, 19) <= input(17);
output(3, 20) <= input(18);
output(3, 21) <= input(19);
output(3, 22) <= input(20);
output(3, 23) <= input(21);
output(3, 24) <= input(22);
output(3, 25) <= input(23);
output(3, 26) <= input(24);
output(3, 27) <= input(25);
output(3, 28) <= input(26);
output(3, 29) <= input(27);
output(3, 30) <= input(28);
output(3, 31) <= input(29);
output(3, 32) <= input(37);
output(3, 33) <= input(35);
output(3, 34) <= input(16);
output(3, 35) <= input(17);
output(3, 36) <= input(18);
output(3, 37) <= input(19);
output(3, 38) <= input(20);
output(3, 39) <= input(21);
output(3, 40) <= input(22);
output(3, 41) <= input(23);
output(3, 42) <= input(24);
output(3, 43) <= input(25);
output(3, 44) <= input(26);
output(3, 45) <= input(27);
output(3, 46) <= input(28);
output(3, 47) <= input(29);
output(3, 48) <= input(37);
output(3, 49) <= input(35);
output(3, 50) <= input(16);
output(3, 51) <= input(17);
output(3, 52) <= input(18);
output(3, 53) <= input(19);
output(3, 54) <= input(20);
output(3, 55) <= input(21);
output(3, 56) <= input(22);
output(3, 57) <= input(23);
output(3, 58) <= input(24);
output(3, 59) <= input(25);
output(3, 60) <= input(26);
output(3, 61) <= input(27);
output(3, 62) <= input(28);
output(3, 63) <= input(29);
output(3, 64) <= input(37);
output(3, 65) <= input(35);
output(3, 66) <= input(16);
output(3, 67) <= input(17);
output(3, 68) <= input(18);
output(3, 69) <= input(19);
output(3, 70) <= input(20);
output(3, 71) <= input(21);
output(3, 72) <= input(22);
output(3, 73) <= input(23);
output(3, 74) <= input(24);
output(3, 75) <= input(25);
output(3, 76) <= input(26);
output(3, 77) <= input(27);
output(3, 78) <= input(28);
output(3, 79) <= input(29);
output(3, 80) <= input(37);
output(3, 81) <= input(35);
output(3, 82) <= input(16);
output(3, 83) <= input(17);
output(3, 84) <= input(18);
output(3, 85) <= input(19);
output(3, 86) <= input(20);
output(3, 87) <= input(21);
output(3, 88) <= input(22);
output(3, 89) <= input(23);
output(3, 90) <= input(24);
output(3, 91) <= input(25);
output(3, 92) <= input(26);
output(3, 93) <= input(27);
output(3, 94) <= input(28);
output(3, 95) <= input(29);
output(3, 96) <= input(37);
output(3, 97) <= input(35);
output(3, 98) <= input(16);
output(3, 99) <= input(17);
output(3, 100) <= input(18);
output(3, 101) <= input(19);
output(3, 102) <= input(20);
output(3, 103) <= input(21);
output(3, 104) <= input(22);
output(3, 105) <= input(23);
output(3, 106) <= input(24);
output(3, 107) <= input(25);
output(3, 108) <= input(26);
output(3, 109) <= input(27);
output(3, 110) <= input(28);
output(3, 111) <= input(29);
output(3, 112) <= input(37);
output(3, 113) <= input(35);
output(3, 114) <= input(16);
output(3, 115) <= input(17);
output(3, 116) <= input(18);
output(3, 117) <= input(19);
output(3, 118) <= input(20);
output(3, 119) <= input(21);
output(3, 120) <= input(22);
output(3, 121) <= input(23);
output(3, 122) <= input(24);
output(3, 123) <= input(25);
output(3, 124) <= input(26);
output(3, 125) <= input(27);
output(3, 126) <= input(28);
output(3, 127) <= input(29);
output(3, 128) <= input(37);
output(3, 129) <= input(35);
output(3, 130) <= input(16);
output(3, 131) <= input(17);
output(3, 132) <= input(18);
output(3, 133) <= input(19);
output(3, 134) <= input(20);
output(3, 135) <= input(21);
output(3, 136) <= input(22);
output(3, 137) <= input(23);
output(3, 138) <= input(24);
output(3, 139) <= input(25);
output(3, 140) <= input(26);
output(3, 141) <= input(27);
output(3, 142) <= input(28);
output(3, 143) <= input(29);
output(3, 144) <= input(37);
output(3, 145) <= input(35);
output(3, 146) <= input(16);
output(3, 147) <= input(17);
output(3, 148) <= input(18);
output(3, 149) <= input(19);
output(3, 150) <= input(20);
output(3, 151) <= input(21);
output(3, 152) <= input(22);
output(3, 153) <= input(23);
output(3, 154) <= input(24);
output(3, 155) <= input(25);
output(3, 156) <= input(26);
output(3, 157) <= input(27);
output(3, 158) <= input(28);
output(3, 159) <= input(29);
output(3, 160) <= input(37);
output(3, 161) <= input(35);
output(3, 162) <= input(16);
output(3, 163) <= input(17);
output(3, 164) <= input(18);
output(3, 165) <= input(19);
output(3, 166) <= input(20);
output(3, 167) <= input(21);
output(3, 168) <= input(22);
output(3, 169) <= input(23);
output(3, 170) <= input(24);
output(3, 171) <= input(25);
output(3, 172) <= input(26);
output(3, 173) <= input(27);
output(3, 174) <= input(28);
output(3, 175) <= input(29);
output(3, 176) <= input(37);
output(3, 177) <= input(35);
output(3, 178) <= input(16);
output(3, 179) <= input(17);
output(3, 180) <= input(18);
output(3, 181) <= input(19);
output(3, 182) <= input(20);
output(3, 183) <= input(21);
output(3, 184) <= input(22);
output(3, 185) <= input(23);
output(3, 186) <= input(24);
output(3, 187) <= input(25);
output(3, 188) <= input(26);
output(3, 189) <= input(27);
output(3, 190) <= input(28);
output(3, 191) <= input(29);
output(3, 192) <= input(37);
output(3, 193) <= input(35);
output(3, 194) <= input(16);
output(3, 195) <= input(17);
output(3, 196) <= input(18);
output(3, 197) <= input(19);
output(3, 198) <= input(20);
output(3, 199) <= input(21);
output(3, 200) <= input(22);
output(3, 201) <= input(23);
output(3, 202) <= input(24);
output(3, 203) <= input(25);
output(3, 204) <= input(26);
output(3, 205) <= input(27);
output(3, 206) <= input(28);
output(3, 207) <= input(29);
output(3, 208) <= input(37);
output(3, 209) <= input(35);
output(3, 210) <= input(16);
output(3, 211) <= input(17);
output(3, 212) <= input(18);
output(3, 213) <= input(19);
output(3, 214) <= input(20);
output(3, 215) <= input(21);
output(3, 216) <= input(22);
output(3, 217) <= input(23);
output(3, 218) <= input(24);
output(3, 219) <= input(25);
output(3, 220) <= input(26);
output(3, 221) <= input(27);
output(3, 222) <= input(28);
output(3, 223) <= input(29);
output(3, 224) <= input(37);
output(3, 225) <= input(35);
output(3, 226) <= input(16);
output(3, 227) <= input(17);
output(3, 228) <= input(18);
output(3, 229) <= input(19);
output(3, 230) <= input(20);
output(3, 231) <= input(21);
output(3, 232) <= input(22);
output(3, 233) <= input(23);
output(3, 234) <= input(24);
output(3, 235) <= input(25);
output(3, 236) <= input(26);
output(3, 237) <= input(27);
output(3, 238) <= input(28);
output(3, 239) <= input(29);
output(3, 240) <= input(36);
output(3, 241) <= input(0);
output(3, 242) <= input(1);
output(3, 243) <= input(2);
output(3, 244) <= input(3);
output(3, 245) <= input(4);
output(3, 246) <= input(5);
output(3, 247) <= input(6);
output(3, 248) <= input(7);
output(3, 249) <= input(8);
output(3, 250) <= input(9);
output(3, 251) <= input(10);
output(3, 252) <= input(11);
output(3, 253) <= input(12);
output(3, 254) <= input(13);
output(3, 255) <= input(14);
output(4, 0) <= input(38);
output(4, 1) <= input(36);
output(4, 2) <= input(0);
output(4, 3) <= input(1);
output(4, 4) <= input(2);
output(4, 5) <= input(3);
output(4, 6) <= input(4);
output(4, 7) <= input(5);
output(4, 8) <= input(6);
output(4, 9) <= input(7);
output(4, 10) <= input(8);
output(4, 11) <= input(9);
output(4, 12) <= input(10);
output(4, 13) <= input(11);
output(4, 14) <= input(12);
output(4, 15) <= input(13);
output(4, 16) <= input(38);
output(4, 17) <= input(36);
output(4, 18) <= input(0);
output(4, 19) <= input(1);
output(4, 20) <= input(2);
output(4, 21) <= input(3);
output(4, 22) <= input(4);
output(4, 23) <= input(5);
output(4, 24) <= input(6);
output(4, 25) <= input(7);
output(4, 26) <= input(8);
output(4, 27) <= input(9);
output(4, 28) <= input(10);
output(4, 29) <= input(11);
output(4, 30) <= input(12);
output(4, 31) <= input(13);
output(4, 32) <= input(38);
output(4, 33) <= input(36);
output(4, 34) <= input(0);
output(4, 35) <= input(1);
output(4, 36) <= input(2);
output(4, 37) <= input(3);
output(4, 38) <= input(4);
output(4, 39) <= input(5);
output(4, 40) <= input(6);
output(4, 41) <= input(7);
output(4, 42) <= input(8);
output(4, 43) <= input(9);
output(4, 44) <= input(10);
output(4, 45) <= input(11);
output(4, 46) <= input(12);
output(4, 47) <= input(13);
output(4, 48) <= input(38);
output(4, 49) <= input(36);
output(4, 50) <= input(0);
output(4, 51) <= input(1);
output(4, 52) <= input(2);
output(4, 53) <= input(3);
output(4, 54) <= input(4);
output(4, 55) <= input(5);
output(4, 56) <= input(6);
output(4, 57) <= input(7);
output(4, 58) <= input(8);
output(4, 59) <= input(9);
output(4, 60) <= input(10);
output(4, 61) <= input(11);
output(4, 62) <= input(12);
output(4, 63) <= input(13);
output(4, 64) <= input(38);
output(4, 65) <= input(36);
output(4, 66) <= input(0);
output(4, 67) <= input(1);
output(4, 68) <= input(2);
output(4, 69) <= input(3);
output(4, 70) <= input(4);
output(4, 71) <= input(5);
output(4, 72) <= input(6);
output(4, 73) <= input(7);
output(4, 74) <= input(8);
output(4, 75) <= input(9);
output(4, 76) <= input(10);
output(4, 77) <= input(11);
output(4, 78) <= input(12);
output(4, 79) <= input(13);
output(4, 80) <= input(38);
output(4, 81) <= input(36);
output(4, 82) <= input(0);
output(4, 83) <= input(1);
output(4, 84) <= input(2);
output(4, 85) <= input(3);
output(4, 86) <= input(4);
output(4, 87) <= input(5);
output(4, 88) <= input(6);
output(4, 89) <= input(7);
output(4, 90) <= input(8);
output(4, 91) <= input(9);
output(4, 92) <= input(10);
output(4, 93) <= input(11);
output(4, 94) <= input(12);
output(4, 95) <= input(13);
output(4, 96) <= input(38);
output(4, 97) <= input(36);
output(4, 98) <= input(0);
output(4, 99) <= input(1);
output(4, 100) <= input(2);
output(4, 101) <= input(3);
output(4, 102) <= input(4);
output(4, 103) <= input(5);
output(4, 104) <= input(6);
output(4, 105) <= input(7);
output(4, 106) <= input(8);
output(4, 107) <= input(9);
output(4, 108) <= input(10);
output(4, 109) <= input(11);
output(4, 110) <= input(12);
output(4, 111) <= input(13);
output(4, 112) <= input(38);
output(4, 113) <= input(36);
output(4, 114) <= input(0);
output(4, 115) <= input(1);
output(4, 116) <= input(2);
output(4, 117) <= input(3);
output(4, 118) <= input(4);
output(4, 119) <= input(5);
output(4, 120) <= input(6);
output(4, 121) <= input(7);
output(4, 122) <= input(8);
output(4, 123) <= input(9);
output(4, 124) <= input(10);
output(4, 125) <= input(11);
output(4, 126) <= input(12);
output(4, 127) <= input(13);
output(4, 128) <= input(38);
output(4, 129) <= input(36);
output(4, 130) <= input(0);
output(4, 131) <= input(1);
output(4, 132) <= input(2);
output(4, 133) <= input(3);
output(4, 134) <= input(4);
output(4, 135) <= input(5);
output(4, 136) <= input(6);
output(4, 137) <= input(7);
output(4, 138) <= input(8);
output(4, 139) <= input(9);
output(4, 140) <= input(10);
output(4, 141) <= input(11);
output(4, 142) <= input(12);
output(4, 143) <= input(13);
output(4, 144) <= input(38);
output(4, 145) <= input(36);
output(4, 146) <= input(0);
output(4, 147) <= input(1);
output(4, 148) <= input(2);
output(4, 149) <= input(3);
output(4, 150) <= input(4);
output(4, 151) <= input(5);
output(4, 152) <= input(6);
output(4, 153) <= input(7);
output(4, 154) <= input(8);
output(4, 155) <= input(9);
output(4, 156) <= input(10);
output(4, 157) <= input(11);
output(4, 158) <= input(12);
output(4, 159) <= input(13);
output(4, 160) <= input(38);
output(4, 161) <= input(36);
output(4, 162) <= input(0);
output(4, 163) <= input(1);
output(4, 164) <= input(2);
output(4, 165) <= input(3);
output(4, 166) <= input(4);
output(4, 167) <= input(5);
output(4, 168) <= input(6);
output(4, 169) <= input(7);
output(4, 170) <= input(8);
output(4, 171) <= input(9);
output(4, 172) <= input(10);
output(4, 173) <= input(11);
output(4, 174) <= input(12);
output(4, 175) <= input(13);
output(4, 176) <= input(38);
output(4, 177) <= input(36);
output(4, 178) <= input(0);
output(4, 179) <= input(1);
output(4, 180) <= input(2);
output(4, 181) <= input(3);
output(4, 182) <= input(4);
output(4, 183) <= input(5);
output(4, 184) <= input(6);
output(4, 185) <= input(7);
output(4, 186) <= input(8);
output(4, 187) <= input(9);
output(4, 188) <= input(10);
output(4, 189) <= input(11);
output(4, 190) <= input(12);
output(4, 191) <= input(13);
output(4, 192) <= input(38);
output(4, 193) <= input(36);
output(4, 194) <= input(0);
output(4, 195) <= input(1);
output(4, 196) <= input(2);
output(4, 197) <= input(3);
output(4, 198) <= input(4);
output(4, 199) <= input(5);
output(4, 200) <= input(6);
output(4, 201) <= input(7);
output(4, 202) <= input(8);
output(4, 203) <= input(9);
output(4, 204) <= input(10);
output(4, 205) <= input(11);
output(4, 206) <= input(12);
output(4, 207) <= input(13);
output(4, 208) <= input(38);
output(4, 209) <= input(36);
output(4, 210) <= input(0);
output(4, 211) <= input(1);
output(4, 212) <= input(2);
output(4, 213) <= input(3);
output(4, 214) <= input(4);
output(4, 215) <= input(5);
output(4, 216) <= input(6);
output(4, 217) <= input(7);
output(4, 218) <= input(8);
output(4, 219) <= input(9);
output(4, 220) <= input(10);
output(4, 221) <= input(11);
output(4, 222) <= input(12);
output(4, 223) <= input(13);
output(4, 224) <= input(38);
output(4, 225) <= input(36);
output(4, 226) <= input(0);
output(4, 227) <= input(1);
output(4, 228) <= input(2);
output(4, 229) <= input(3);
output(4, 230) <= input(4);
output(4, 231) <= input(5);
output(4, 232) <= input(6);
output(4, 233) <= input(7);
output(4, 234) <= input(8);
output(4, 235) <= input(9);
output(4, 236) <= input(10);
output(4, 237) <= input(11);
output(4, 238) <= input(12);
output(4, 239) <= input(13);
output(4, 240) <= input(38);
output(4, 241) <= input(36);
output(4, 242) <= input(0);
output(4, 243) <= input(1);
output(4, 244) <= input(2);
output(4, 245) <= input(3);
output(4, 246) <= input(4);
output(4, 247) <= input(5);
output(4, 248) <= input(6);
output(4, 249) <= input(7);
output(4, 250) <= input(8);
output(4, 251) <= input(9);
output(4, 252) <= input(10);
output(4, 253) <= input(11);
output(4, 254) <= input(12);
output(4, 255) <= input(13);
output(5, 0) <= input(39);
output(5, 1) <= input(38);
output(5, 2) <= input(36);
output(5, 3) <= input(0);
output(5, 4) <= input(1);
output(5, 5) <= input(2);
output(5, 6) <= input(3);
output(5, 7) <= input(4);
output(5, 8) <= input(5);
output(5, 9) <= input(6);
output(5, 10) <= input(7);
output(5, 11) <= input(8);
output(5, 12) <= input(9);
output(5, 13) <= input(10);
output(5, 14) <= input(11);
output(5, 15) <= input(12);
output(5, 16) <= input(39);
output(5, 17) <= input(38);
output(5, 18) <= input(36);
output(5, 19) <= input(0);
output(5, 20) <= input(1);
output(5, 21) <= input(2);
output(5, 22) <= input(3);
output(5, 23) <= input(4);
output(5, 24) <= input(5);
output(5, 25) <= input(6);
output(5, 26) <= input(7);
output(5, 27) <= input(8);
output(5, 28) <= input(9);
output(5, 29) <= input(10);
output(5, 30) <= input(11);
output(5, 31) <= input(12);
output(5, 32) <= input(39);
output(5, 33) <= input(38);
output(5, 34) <= input(36);
output(5, 35) <= input(0);
output(5, 36) <= input(1);
output(5, 37) <= input(2);
output(5, 38) <= input(3);
output(5, 39) <= input(4);
output(5, 40) <= input(5);
output(5, 41) <= input(6);
output(5, 42) <= input(7);
output(5, 43) <= input(8);
output(5, 44) <= input(9);
output(5, 45) <= input(10);
output(5, 46) <= input(11);
output(5, 47) <= input(12);
output(5, 48) <= input(39);
output(5, 49) <= input(38);
output(5, 50) <= input(36);
output(5, 51) <= input(0);
output(5, 52) <= input(1);
output(5, 53) <= input(2);
output(5, 54) <= input(3);
output(5, 55) <= input(4);
output(5, 56) <= input(5);
output(5, 57) <= input(6);
output(5, 58) <= input(7);
output(5, 59) <= input(8);
output(5, 60) <= input(9);
output(5, 61) <= input(10);
output(5, 62) <= input(11);
output(5, 63) <= input(12);
output(5, 64) <= input(39);
output(5, 65) <= input(38);
output(5, 66) <= input(36);
output(5, 67) <= input(0);
output(5, 68) <= input(1);
output(5, 69) <= input(2);
output(5, 70) <= input(3);
output(5, 71) <= input(4);
output(5, 72) <= input(5);
output(5, 73) <= input(6);
output(5, 74) <= input(7);
output(5, 75) <= input(8);
output(5, 76) <= input(9);
output(5, 77) <= input(10);
output(5, 78) <= input(11);
output(5, 79) <= input(12);
output(5, 80) <= input(39);
output(5, 81) <= input(38);
output(5, 82) <= input(36);
output(5, 83) <= input(0);
output(5, 84) <= input(1);
output(5, 85) <= input(2);
output(5, 86) <= input(3);
output(5, 87) <= input(4);
output(5, 88) <= input(5);
output(5, 89) <= input(6);
output(5, 90) <= input(7);
output(5, 91) <= input(8);
output(5, 92) <= input(9);
output(5, 93) <= input(10);
output(5, 94) <= input(11);
output(5, 95) <= input(12);
output(5, 96) <= input(39);
output(5, 97) <= input(38);
output(5, 98) <= input(36);
output(5, 99) <= input(0);
output(5, 100) <= input(1);
output(5, 101) <= input(2);
output(5, 102) <= input(3);
output(5, 103) <= input(4);
output(5, 104) <= input(5);
output(5, 105) <= input(6);
output(5, 106) <= input(7);
output(5, 107) <= input(8);
output(5, 108) <= input(9);
output(5, 109) <= input(10);
output(5, 110) <= input(11);
output(5, 111) <= input(12);
output(5, 112) <= input(39);
output(5, 113) <= input(38);
output(5, 114) <= input(36);
output(5, 115) <= input(0);
output(5, 116) <= input(1);
output(5, 117) <= input(2);
output(5, 118) <= input(3);
output(5, 119) <= input(4);
output(5, 120) <= input(5);
output(5, 121) <= input(6);
output(5, 122) <= input(7);
output(5, 123) <= input(8);
output(5, 124) <= input(9);
output(5, 125) <= input(10);
output(5, 126) <= input(11);
output(5, 127) <= input(12);
output(5, 128) <= input(39);
output(5, 129) <= input(38);
output(5, 130) <= input(36);
output(5, 131) <= input(0);
output(5, 132) <= input(1);
output(5, 133) <= input(2);
output(5, 134) <= input(3);
output(5, 135) <= input(4);
output(5, 136) <= input(5);
output(5, 137) <= input(6);
output(5, 138) <= input(7);
output(5, 139) <= input(8);
output(5, 140) <= input(9);
output(5, 141) <= input(10);
output(5, 142) <= input(11);
output(5, 143) <= input(12);
output(5, 144) <= input(39);
output(5, 145) <= input(38);
output(5, 146) <= input(36);
output(5, 147) <= input(0);
output(5, 148) <= input(1);
output(5, 149) <= input(2);
output(5, 150) <= input(3);
output(5, 151) <= input(4);
output(5, 152) <= input(5);
output(5, 153) <= input(6);
output(5, 154) <= input(7);
output(5, 155) <= input(8);
output(5, 156) <= input(9);
output(5, 157) <= input(10);
output(5, 158) <= input(11);
output(5, 159) <= input(12);
output(5, 160) <= input(39);
output(5, 161) <= input(38);
output(5, 162) <= input(36);
output(5, 163) <= input(0);
output(5, 164) <= input(1);
output(5, 165) <= input(2);
output(5, 166) <= input(3);
output(5, 167) <= input(4);
output(5, 168) <= input(5);
output(5, 169) <= input(6);
output(5, 170) <= input(7);
output(5, 171) <= input(8);
output(5, 172) <= input(9);
output(5, 173) <= input(10);
output(5, 174) <= input(11);
output(5, 175) <= input(12);
output(5, 176) <= input(39);
output(5, 177) <= input(38);
output(5, 178) <= input(36);
output(5, 179) <= input(0);
output(5, 180) <= input(1);
output(5, 181) <= input(2);
output(5, 182) <= input(3);
output(5, 183) <= input(4);
output(5, 184) <= input(5);
output(5, 185) <= input(6);
output(5, 186) <= input(7);
output(5, 187) <= input(8);
output(5, 188) <= input(9);
output(5, 189) <= input(10);
output(5, 190) <= input(11);
output(5, 191) <= input(12);
output(5, 192) <= input(39);
output(5, 193) <= input(38);
output(5, 194) <= input(36);
output(5, 195) <= input(0);
output(5, 196) <= input(1);
output(5, 197) <= input(2);
output(5, 198) <= input(3);
output(5, 199) <= input(4);
output(5, 200) <= input(5);
output(5, 201) <= input(6);
output(5, 202) <= input(7);
output(5, 203) <= input(8);
output(5, 204) <= input(9);
output(5, 205) <= input(10);
output(5, 206) <= input(11);
output(5, 207) <= input(12);
output(5, 208) <= input(39);
output(5, 209) <= input(38);
output(5, 210) <= input(36);
output(5, 211) <= input(0);
output(5, 212) <= input(1);
output(5, 213) <= input(2);
output(5, 214) <= input(3);
output(5, 215) <= input(4);
output(5, 216) <= input(5);
output(5, 217) <= input(6);
output(5, 218) <= input(7);
output(5, 219) <= input(8);
output(5, 220) <= input(9);
output(5, 221) <= input(10);
output(5, 222) <= input(11);
output(5, 223) <= input(12);
output(5, 224) <= input(39);
output(5, 225) <= input(38);
output(5, 226) <= input(36);
output(5, 227) <= input(0);
output(5, 228) <= input(1);
output(5, 229) <= input(2);
output(5, 230) <= input(3);
output(5, 231) <= input(4);
output(5, 232) <= input(5);
output(5, 233) <= input(6);
output(5, 234) <= input(7);
output(5, 235) <= input(8);
output(5, 236) <= input(9);
output(5, 237) <= input(10);
output(5, 238) <= input(11);
output(5, 239) <= input(12);
output(5, 240) <= input(39);
output(5, 241) <= input(38);
output(5, 242) <= input(36);
output(5, 243) <= input(0);
output(5, 244) <= input(1);
output(5, 245) <= input(2);
output(5, 246) <= input(3);
output(5, 247) <= input(4);
output(5, 248) <= input(5);
output(5, 249) <= input(6);
output(5, 250) <= input(7);
output(5, 251) <= input(8);
output(5, 252) <= input(9);
output(5, 253) <= input(10);
output(5, 254) <= input(11);
output(5, 255) <= input(12);
output(6, 0) <= input(40);
output(6, 1) <= input(41);
output(6, 2) <= input(37);
output(6, 3) <= input(35);
output(6, 4) <= input(16);
output(6, 5) <= input(17);
output(6, 6) <= input(18);
output(6, 7) <= input(19);
output(6, 8) <= input(20);
output(6, 9) <= input(21);
output(6, 10) <= input(22);
output(6, 11) <= input(23);
output(6, 12) <= input(24);
output(6, 13) <= input(25);
output(6, 14) <= input(26);
output(6, 15) <= input(27);
output(6, 16) <= input(40);
output(6, 17) <= input(41);
output(6, 18) <= input(37);
output(6, 19) <= input(35);
output(6, 20) <= input(16);
output(6, 21) <= input(17);
output(6, 22) <= input(18);
output(6, 23) <= input(19);
output(6, 24) <= input(20);
output(6, 25) <= input(21);
output(6, 26) <= input(22);
output(6, 27) <= input(23);
output(6, 28) <= input(24);
output(6, 29) <= input(25);
output(6, 30) <= input(26);
output(6, 31) <= input(27);
output(6, 32) <= input(40);
output(6, 33) <= input(41);
output(6, 34) <= input(37);
output(6, 35) <= input(35);
output(6, 36) <= input(16);
output(6, 37) <= input(17);
output(6, 38) <= input(18);
output(6, 39) <= input(19);
output(6, 40) <= input(20);
output(6, 41) <= input(21);
output(6, 42) <= input(22);
output(6, 43) <= input(23);
output(6, 44) <= input(24);
output(6, 45) <= input(25);
output(6, 46) <= input(26);
output(6, 47) <= input(27);
output(6, 48) <= input(40);
output(6, 49) <= input(41);
output(6, 50) <= input(37);
output(6, 51) <= input(35);
output(6, 52) <= input(16);
output(6, 53) <= input(17);
output(6, 54) <= input(18);
output(6, 55) <= input(19);
output(6, 56) <= input(20);
output(6, 57) <= input(21);
output(6, 58) <= input(22);
output(6, 59) <= input(23);
output(6, 60) <= input(24);
output(6, 61) <= input(25);
output(6, 62) <= input(26);
output(6, 63) <= input(27);
output(6, 64) <= input(40);
output(6, 65) <= input(41);
output(6, 66) <= input(37);
output(6, 67) <= input(35);
output(6, 68) <= input(16);
output(6, 69) <= input(17);
output(6, 70) <= input(18);
output(6, 71) <= input(19);
output(6, 72) <= input(20);
output(6, 73) <= input(21);
output(6, 74) <= input(22);
output(6, 75) <= input(23);
output(6, 76) <= input(24);
output(6, 77) <= input(25);
output(6, 78) <= input(26);
output(6, 79) <= input(27);
output(6, 80) <= input(40);
output(6, 81) <= input(41);
output(6, 82) <= input(37);
output(6, 83) <= input(35);
output(6, 84) <= input(16);
output(6, 85) <= input(17);
output(6, 86) <= input(18);
output(6, 87) <= input(19);
output(6, 88) <= input(20);
output(6, 89) <= input(21);
output(6, 90) <= input(22);
output(6, 91) <= input(23);
output(6, 92) <= input(24);
output(6, 93) <= input(25);
output(6, 94) <= input(26);
output(6, 95) <= input(27);
output(6, 96) <= input(40);
output(6, 97) <= input(41);
output(6, 98) <= input(37);
output(6, 99) <= input(35);
output(6, 100) <= input(16);
output(6, 101) <= input(17);
output(6, 102) <= input(18);
output(6, 103) <= input(19);
output(6, 104) <= input(20);
output(6, 105) <= input(21);
output(6, 106) <= input(22);
output(6, 107) <= input(23);
output(6, 108) <= input(24);
output(6, 109) <= input(25);
output(6, 110) <= input(26);
output(6, 111) <= input(27);
output(6, 112) <= input(40);
output(6, 113) <= input(41);
output(6, 114) <= input(37);
output(6, 115) <= input(35);
output(6, 116) <= input(16);
output(6, 117) <= input(17);
output(6, 118) <= input(18);
output(6, 119) <= input(19);
output(6, 120) <= input(20);
output(6, 121) <= input(21);
output(6, 122) <= input(22);
output(6, 123) <= input(23);
output(6, 124) <= input(24);
output(6, 125) <= input(25);
output(6, 126) <= input(26);
output(6, 127) <= input(27);
output(6, 128) <= input(42);
output(6, 129) <= input(39);
output(6, 130) <= input(38);
output(6, 131) <= input(36);
output(6, 132) <= input(0);
output(6, 133) <= input(1);
output(6, 134) <= input(2);
output(6, 135) <= input(3);
output(6, 136) <= input(4);
output(6, 137) <= input(5);
output(6, 138) <= input(6);
output(6, 139) <= input(7);
output(6, 140) <= input(8);
output(6, 141) <= input(9);
output(6, 142) <= input(10);
output(6, 143) <= input(11);
output(6, 144) <= input(42);
output(6, 145) <= input(39);
output(6, 146) <= input(38);
output(6, 147) <= input(36);
output(6, 148) <= input(0);
output(6, 149) <= input(1);
output(6, 150) <= input(2);
output(6, 151) <= input(3);
output(6, 152) <= input(4);
output(6, 153) <= input(5);
output(6, 154) <= input(6);
output(6, 155) <= input(7);
output(6, 156) <= input(8);
output(6, 157) <= input(9);
output(6, 158) <= input(10);
output(6, 159) <= input(11);
output(6, 160) <= input(42);
output(6, 161) <= input(39);
output(6, 162) <= input(38);
output(6, 163) <= input(36);
output(6, 164) <= input(0);
output(6, 165) <= input(1);
output(6, 166) <= input(2);
output(6, 167) <= input(3);
output(6, 168) <= input(4);
output(6, 169) <= input(5);
output(6, 170) <= input(6);
output(6, 171) <= input(7);
output(6, 172) <= input(8);
output(6, 173) <= input(9);
output(6, 174) <= input(10);
output(6, 175) <= input(11);
output(6, 176) <= input(42);
output(6, 177) <= input(39);
output(6, 178) <= input(38);
output(6, 179) <= input(36);
output(6, 180) <= input(0);
output(6, 181) <= input(1);
output(6, 182) <= input(2);
output(6, 183) <= input(3);
output(6, 184) <= input(4);
output(6, 185) <= input(5);
output(6, 186) <= input(6);
output(6, 187) <= input(7);
output(6, 188) <= input(8);
output(6, 189) <= input(9);
output(6, 190) <= input(10);
output(6, 191) <= input(11);
output(6, 192) <= input(42);
output(6, 193) <= input(39);
output(6, 194) <= input(38);
output(6, 195) <= input(36);
output(6, 196) <= input(0);
output(6, 197) <= input(1);
output(6, 198) <= input(2);
output(6, 199) <= input(3);
output(6, 200) <= input(4);
output(6, 201) <= input(5);
output(6, 202) <= input(6);
output(6, 203) <= input(7);
output(6, 204) <= input(8);
output(6, 205) <= input(9);
output(6, 206) <= input(10);
output(6, 207) <= input(11);
output(6, 208) <= input(42);
output(6, 209) <= input(39);
output(6, 210) <= input(38);
output(6, 211) <= input(36);
output(6, 212) <= input(0);
output(6, 213) <= input(1);
output(6, 214) <= input(2);
output(6, 215) <= input(3);
output(6, 216) <= input(4);
output(6, 217) <= input(5);
output(6, 218) <= input(6);
output(6, 219) <= input(7);
output(6, 220) <= input(8);
output(6, 221) <= input(9);
output(6, 222) <= input(10);
output(6, 223) <= input(11);
output(6, 224) <= input(42);
output(6, 225) <= input(39);
output(6, 226) <= input(38);
output(6, 227) <= input(36);
output(6, 228) <= input(0);
output(6, 229) <= input(1);
output(6, 230) <= input(2);
output(6, 231) <= input(3);
output(6, 232) <= input(4);
output(6, 233) <= input(5);
output(6, 234) <= input(6);
output(6, 235) <= input(7);
output(6, 236) <= input(8);
output(6, 237) <= input(9);
output(6, 238) <= input(10);
output(6, 239) <= input(11);
output(6, 240) <= input(42);
output(6, 241) <= input(39);
output(6, 242) <= input(38);
output(6, 243) <= input(36);
output(6, 244) <= input(0);
output(6, 245) <= input(1);
output(6, 246) <= input(2);
output(6, 247) <= input(3);
output(6, 248) <= input(4);
output(6, 249) <= input(5);
output(6, 250) <= input(6);
output(6, 251) <= input(7);
output(6, 252) <= input(8);
output(6, 253) <= input(9);
output(6, 254) <= input(10);
output(6, 255) <= input(11);
output(7, 0) <= input(42);
output(7, 1) <= input(39);
output(7, 2) <= input(38);
output(7, 3) <= input(36);
output(7, 4) <= input(0);
output(7, 5) <= input(1);
output(7, 6) <= input(2);
output(7, 7) <= input(3);
output(7, 8) <= input(4);
output(7, 9) <= input(5);
output(7, 10) <= input(6);
output(7, 11) <= input(7);
output(7, 12) <= input(8);
output(7, 13) <= input(9);
output(7, 14) <= input(10);
output(7, 15) <= input(11);
output(7, 16) <= input(42);
output(7, 17) <= input(39);
output(7, 18) <= input(38);
output(7, 19) <= input(36);
output(7, 20) <= input(0);
output(7, 21) <= input(1);
output(7, 22) <= input(2);
output(7, 23) <= input(3);
output(7, 24) <= input(4);
output(7, 25) <= input(5);
output(7, 26) <= input(6);
output(7, 27) <= input(7);
output(7, 28) <= input(8);
output(7, 29) <= input(9);
output(7, 30) <= input(10);
output(7, 31) <= input(11);
output(7, 32) <= input(42);
output(7, 33) <= input(39);
output(7, 34) <= input(38);
output(7, 35) <= input(36);
output(7, 36) <= input(0);
output(7, 37) <= input(1);
output(7, 38) <= input(2);
output(7, 39) <= input(3);
output(7, 40) <= input(4);
output(7, 41) <= input(5);
output(7, 42) <= input(6);
output(7, 43) <= input(7);
output(7, 44) <= input(8);
output(7, 45) <= input(9);
output(7, 46) <= input(10);
output(7, 47) <= input(11);
output(7, 48) <= input(42);
output(7, 49) <= input(39);
output(7, 50) <= input(38);
output(7, 51) <= input(36);
output(7, 52) <= input(0);
output(7, 53) <= input(1);
output(7, 54) <= input(2);
output(7, 55) <= input(3);
output(7, 56) <= input(4);
output(7, 57) <= input(5);
output(7, 58) <= input(6);
output(7, 59) <= input(7);
output(7, 60) <= input(8);
output(7, 61) <= input(9);
output(7, 62) <= input(10);
output(7, 63) <= input(11);
output(7, 64) <= input(42);
output(7, 65) <= input(39);
output(7, 66) <= input(38);
output(7, 67) <= input(36);
output(7, 68) <= input(0);
output(7, 69) <= input(1);
output(7, 70) <= input(2);
output(7, 71) <= input(3);
output(7, 72) <= input(4);
output(7, 73) <= input(5);
output(7, 74) <= input(6);
output(7, 75) <= input(7);
output(7, 76) <= input(8);
output(7, 77) <= input(9);
output(7, 78) <= input(10);
output(7, 79) <= input(11);
output(7, 80) <= input(43);
output(7, 81) <= input(40);
output(7, 82) <= input(41);
output(7, 83) <= input(37);
output(7, 84) <= input(35);
output(7, 85) <= input(16);
output(7, 86) <= input(17);
output(7, 87) <= input(18);
output(7, 88) <= input(19);
output(7, 89) <= input(20);
output(7, 90) <= input(21);
output(7, 91) <= input(22);
output(7, 92) <= input(23);
output(7, 93) <= input(24);
output(7, 94) <= input(25);
output(7, 95) <= input(26);
output(7, 96) <= input(43);
output(7, 97) <= input(40);
output(7, 98) <= input(41);
output(7, 99) <= input(37);
output(7, 100) <= input(35);
output(7, 101) <= input(16);
output(7, 102) <= input(17);
output(7, 103) <= input(18);
output(7, 104) <= input(19);
output(7, 105) <= input(20);
output(7, 106) <= input(21);
output(7, 107) <= input(22);
output(7, 108) <= input(23);
output(7, 109) <= input(24);
output(7, 110) <= input(25);
output(7, 111) <= input(26);
output(7, 112) <= input(43);
output(7, 113) <= input(40);
output(7, 114) <= input(41);
output(7, 115) <= input(37);
output(7, 116) <= input(35);
output(7, 117) <= input(16);
output(7, 118) <= input(17);
output(7, 119) <= input(18);
output(7, 120) <= input(19);
output(7, 121) <= input(20);
output(7, 122) <= input(21);
output(7, 123) <= input(22);
output(7, 124) <= input(23);
output(7, 125) <= input(24);
output(7, 126) <= input(25);
output(7, 127) <= input(26);
output(7, 128) <= input(43);
output(7, 129) <= input(40);
output(7, 130) <= input(41);
output(7, 131) <= input(37);
output(7, 132) <= input(35);
output(7, 133) <= input(16);
output(7, 134) <= input(17);
output(7, 135) <= input(18);
output(7, 136) <= input(19);
output(7, 137) <= input(20);
output(7, 138) <= input(21);
output(7, 139) <= input(22);
output(7, 140) <= input(23);
output(7, 141) <= input(24);
output(7, 142) <= input(25);
output(7, 143) <= input(26);
output(7, 144) <= input(43);
output(7, 145) <= input(40);
output(7, 146) <= input(41);
output(7, 147) <= input(37);
output(7, 148) <= input(35);
output(7, 149) <= input(16);
output(7, 150) <= input(17);
output(7, 151) <= input(18);
output(7, 152) <= input(19);
output(7, 153) <= input(20);
output(7, 154) <= input(21);
output(7, 155) <= input(22);
output(7, 156) <= input(23);
output(7, 157) <= input(24);
output(7, 158) <= input(25);
output(7, 159) <= input(26);
output(7, 160) <= input(44);
output(7, 161) <= input(42);
output(7, 162) <= input(39);
output(7, 163) <= input(38);
output(7, 164) <= input(36);
output(7, 165) <= input(0);
output(7, 166) <= input(1);
output(7, 167) <= input(2);
output(7, 168) <= input(3);
output(7, 169) <= input(4);
output(7, 170) <= input(5);
output(7, 171) <= input(6);
output(7, 172) <= input(7);
output(7, 173) <= input(8);
output(7, 174) <= input(9);
output(7, 175) <= input(10);
output(7, 176) <= input(44);
output(7, 177) <= input(42);
output(7, 178) <= input(39);
output(7, 179) <= input(38);
output(7, 180) <= input(36);
output(7, 181) <= input(0);
output(7, 182) <= input(1);
output(7, 183) <= input(2);
output(7, 184) <= input(3);
output(7, 185) <= input(4);
output(7, 186) <= input(5);
output(7, 187) <= input(6);
output(7, 188) <= input(7);
output(7, 189) <= input(8);
output(7, 190) <= input(9);
output(7, 191) <= input(10);
output(7, 192) <= input(44);
output(7, 193) <= input(42);
output(7, 194) <= input(39);
output(7, 195) <= input(38);
output(7, 196) <= input(36);
output(7, 197) <= input(0);
output(7, 198) <= input(1);
output(7, 199) <= input(2);
output(7, 200) <= input(3);
output(7, 201) <= input(4);
output(7, 202) <= input(5);
output(7, 203) <= input(6);
output(7, 204) <= input(7);
output(7, 205) <= input(8);
output(7, 206) <= input(9);
output(7, 207) <= input(10);
output(7, 208) <= input(44);
output(7, 209) <= input(42);
output(7, 210) <= input(39);
output(7, 211) <= input(38);
output(7, 212) <= input(36);
output(7, 213) <= input(0);
output(7, 214) <= input(1);
output(7, 215) <= input(2);
output(7, 216) <= input(3);
output(7, 217) <= input(4);
output(7, 218) <= input(5);
output(7, 219) <= input(6);
output(7, 220) <= input(7);
output(7, 221) <= input(8);
output(7, 222) <= input(9);
output(7, 223) <= input(10);
output(7, 224) <= input(44);
output(7, 225) <= input(42);
output(7, 226) <= input(39);
output(7, 227) <= input(38);
output(7, 228) <= input(36);
output(7, 229) <= input(0);
output(7, 230) <= input(1);
output(7, 231) <= input(2);
output(7, 232) <= input(3);
output(7, 233) <= input(4);
output(7, 234) <= input(5);
output(7, 235) <= input(6);
output(7, 236) <= input(7);
output(7, 237) <= input(8);
output(7, 238) <= input(9);
output(7, 239) <= input(10);
output(7, 240) <= input(44);
output(7, 241) <= input(42);
output(7, 242) <= input(39);
output(7, 243) <= input(38);
output(7, 244) <= input(36);
output(7, 245) <= input(0);
output(7, 246) <= input(1);
output(7, 247) <= input(2);
output(7, 248) <= input(3);
output(7, 249) <= input(4);
output(7, 250) <= input(5);
output(7, 251) <= input(6);
output(7, 252) <= input(7);
output(7, 253) <= input(8);
output(7, 254) <= input(9);
output(7, 255) <= input(10);
when "0011" =>
output(0, 0) <= input(0);
output(0, 1) <= input(1);
output(0, 2) <= input(2);
output(0, 3) <= input(3);
output(0, 4) <= input(4);
output(0, 5) <= input(5);
output(0, 6) <= input(6);
output(0, 7) <= input(7);
output(0, 8) <= input(8);
output(0, 9) <= input(9);
output(0, 10) <= input(10);
output(0, 11) <= input(11);
output(0, 12) <= input(12);
output(0, 13) <= input(13);
output(0, 14) <= input(14);
output(0, 15) <= input(15);
output(0, 16) <= input(0);
output(0, 17) <= input(1);
output(0, 18) <= input(2);
output(0, 19) <= input(3);
output(0, 20) <= input(4);
output(0, 21) <= input(5);
output(0, 22) <= input(6);
output(0, 23) <= input(7);
output(0, 24) <= input(8);
output(0, 25) <= input(9);
output(0, 26) <= input(10);
output(0, 27) <= input(11);
output(0, 28) <= input(12);
output(0, 29) <= input(13);
output(0, 30) <= input(14);
output(0, 31) <= input(15);
output(0, 32) <= input(0);
output(0, 33) <= input(1);
output(0, 34) <= input(2);
output(0, 35) <= input(3);
output(0, 36) <= input(4);
output(0, 37) <= input(5);
output(0, 38) <= input(6);
output(0, 39) <= input(7);
output(0, 40) <= input(8);
output(0, 41) <= input(9);
output(0, 42) <= input(10);
output(0, 43) <= input(11);
output(0, 44) <= input(12);
output(0, 45) <= input(13);
output(0, 46) <= input(14);
output(0, 47) <= input(15);
output(0, 48) <= input(0);
output(0, 49) <= input(1);
output(0, 50) <= input(2);
output(0, 51) <= input(3);
output(0, 52) <= input(4);
output(0, 53) <= input(5);
output(0, 54) <= input(6);
output(0, 55) <= input(7);
output(0, 56) <= input(8);
output(0, 57) <= input(9);
output(0, 58) <= input(10);
output(0, 59) <= input(11);
output(0, 60) <= input(12);
output(0, 61) <= input(13);
output(0, 62) <= input(14);
output(0, 63) <= input(15);
output(0, 64) <= input(16);
output(0, 65) <= input(17);
output(0, 66) <= input(18);
output(0, 67) <= input(19);
output(0, 68) <= input(20);
output(0, 69) <= input(21);
output(0, 70) <= input(22);
output(0, 71) <= input(23);
output(0, 72) <= input(24);
output(0, 73) <= input(25);
output(0, 74) <= input(26);
output(0, 75) <= input(27);
output(0, 76) <= input(28);
output(0, 77) <= input(29);
output(0, 78) <= input(30);
output(0, 79) <= input(31);
output(0, 80) <= input(16);
output(0, 81) <= input(17);
output(0, 82) <= input(18);
output(0, 83) <= input(19);
output(0, 84) <= input(20);
output(0, 85) <= input(21);
output(0, 86) <= input(22);
output(0, 87) <= input(23);
output(0, 88) <= input(24);
output(0, 89) <= input(25);
output(0, 90) <= input(26);
output(0, 91) <= input(27);
output(0, 92) <= input(28);
output(0, 93) <= input(29);
output(0, 94) <= input(30);
output(0, 95) <= input(31);
output(0, 96) <= input(16);
output(0, 97) <= input(17);
output(0, 98) <= input(18);
output(0, 99) <= input(19);
output(0, 100) <= input(20);
output(0, 101) <= input(21);
output(0, 102) <= input(22);
output(0, 103) <= input(23);
output(0, 104) <= input(24);
output(0, 105) <= input(25);
output(0, 106) <= input(26);
output(0, 107) <= input(27);
output(0, 108) <= input(28);
output(0, 109) <= input(29);
output(0, 110) <= input(30);
output(0, 111) <= input(31);
output(0, 112) <= input(16);
output(0, 113) <= input(17);
output(0, 114) <= input(18);
output(0, 115) <= input(19);
output(0, 116) <= input(20);
output(0, 117) <= input(21);
output(0, 118) <= input(22);
output(0, 119) <= input(23);
output(0, 120) <= input(24);
output(0, 121) <= input(25);
output(0, 122) <= input(26);
output(0, 123) <= input(27);
output(0, 124) <= input(28);
output(0, 125) <= input(29);
output(0, 126) <= input(30);
output(0, 127) <= input(31);
output(0, 128) <= input(32);
output(0, 129) <= input(0);
output(0, 130) <= input(1);
output(0, 131) <= input(2);
output(0, 132) <= input(3);
output(0, 133) <= input(4);
output(0, 134) <= input(5);
output(0, 135) <= input(6);
output(0, 136) <= input(7);
output(0, 137) <= input(8);
output(0, 138) <= input(9);
output(0, 139) <= input(10);
output(0, 140) <= input(11);
output(0, 141) <= input(12);
output(0, 142) <= input(13);
output(0, 143) <= input(14);
output(0, 144) <= input(32);
output(0, 145) <= input(0);
output(0, 146) <= input(1);
output(0, 147) <= input(2);
output(0, 148) <= input(3);
output(0, 149) <= input(4);
output(0, 150) <= input(5);
output(0, 151) <= input(6);
output(0, 152) <= input(7);
output(0, 153) <= input(8);
output(0, 154) <= input(9);
output(0, 155) <= input(10);
output(0, 156) <= input(11);
output(0, 157) <= input(12);
output(0, 158) <= input(13);
output(0, 159) <= input(14);
output(0, 160) <= input(32);
output(0, 161) <= input(0);
output(0, 162) <= input(1);
output(0, 163) <= input(2);
output(0, 164) <= input(3);
output(0, 165) <= input(4);
output(0, 166) <= input(5);
output(0, 167) <= input(6);
output(0, 168) <= input(7);
output(0, 169) <= input(8);
output(0, 170) <= input(9);
output(0, 171) <= input(10);
output(0, 172) <= input(11);
output(0, 173) <= input(12);
output(0, 174) <= input(13);
output(0, 175) <= input(14);
output(0, 176) <= input(32);
output(0, 177) <= input(0);
output(0, 178) <= input(1);
output(0, 179) <= input(2);
output(0, 180) <= input(3);
output(0, 181) <= input(4);
output(0, 182) <= input(5);
output(0, 183) <= input(6);
output(0, 184) <= input(7);
output(0, 185) <= input(8);
output(0, 186) <= input(9);
output(0, 187) <= input(10);
output(0, 188) <= input(11);
output(0, 189) <= input(12);
output(0, 190) <= input(13);
output(0, 191) <= input(14);
output(0, 192) <= input(33);
output(0, 193) <= input(16);
output(0, 194) <= input(17);
output(0, 195) <= input(18);
output(0, 196) <= input(19);
output(0, 197) <= input(20);
output(0, 198) <= input(21);
output(0, 199) <= input(22);
output(0, 200) <= input(23);
output(0, 201) <= input(24);
output(0, 202) <= input(25);
output(0, 203) <= input(26);
output(0, 204) <= input(27);
output(0, 205) <= input(28);
output(0, 206) <= input(29);
output(0, 207) <= input(30);
output(0, 208) <= input(33);
output(0, 209) <= input(16);
output(0, 210) <= input(17);
output(0, 211) <= input(18);
output(0, 212) <= input(19);
output(0, 213) <= input(20);
output(0, 214) <= input(21);
output(0, 215) <= input(22);
output(0, 216) <= input(23);
output(0, 217) <= input(24);
output(0, 218) <= input(25);
output(0, 219) <= input(26);
output(0, 220) <= input(27);
output(0, 221) <= input(28);
output(0, 222) <= input(29);
output(0, 223) <= input(30);
output(0, 224) <= input(33);
output(0, 225) <= input(16);
output(0, 226) <= input(17);
output(0, 227) <= input(18);
output(0, 228) <= input(19);
output(0, 229) <= input(20);
output(0, 230) <= input(21);
output(0, 231) <= input(22);
output(0, 232) <= input(23);
output(0, 233) <= input(24);
output(0, 234) <= input(25);
output(0, 235) <= input(26);
output(0, 236) <= input(27);
output(0, 237) <= input(28);
output(0, 238) <= input(29);
output(0, 239) <= input(30);
output(0, 240) <= input(33);
output(0, 241) <= input(16);
output(0, 242) <= input(17);
output(0, 243) <= input(18);
output(0, 244) <= input(19);
output(0, 245) <= input(20);
output(0, 246) <= input(21);
output(0, 247) <= input(22);
output(0, 248) <= input(23);
output(0, 249) <= input(24);
output(0, 250) <= input(25);
output(0, 251) <= input(26);
output(0, 252) <= input(27);
output(0, 253) <= input(28);
output(0, 254) <= input(29);
output(0, 255) <= input(30);
output(1, 0) <= input(32);
output(1, 1) <= input(0);
output(1, 2) <= input(1);
output(1, 3) <= input(2);
output(1, 4) <= input(3);
output(1, 5) <= input(4);
output(1, 6) <= input(5);
output(1, 7) <= input(6);
output(1, 8) <= input(7);
output(1, 9) <= input(8);
output(1, 10) <= input(9);
output(1, 11) <= input(10);
output(1, 12) <= input(11);
output(1, 13) <= input(12);
output(1, 14) <= input(13);
output(1, 15) <= input(14);
output(1, 16) <= input(32);
output(1, 17) <= input(0);
output(1, 18) <= input(1);
output(1, 19) <= input(2);
output(1, 20) <= input(3);
output(1, 21) <= input(4);
output(1, 22) <= input(5);
output(1, 23) <= input(6);
output(1, 24) <= input(7);
output(1, 25) <= input(8);
output(1, 26) <= input(9);
output(1, 27) <= input(10);
output(1, 28) <= input(11);
output(1, 29) <= input(12);
output(1, 30) <= input(13);
output(1, 31) <= input(14);
output(1, 32) <= input(33);
output(1, 33) <= input(16);
output(1, 34) <= input(17);
output(1, 35) <= input(18);
output(1, 36) <= input(19);
output(1, 37) <= input(20);
output(1, 38) <= input(21);
output(1, 39) <= input(22);
output(1, 40) <= input(23);
output(1, 41) <= input(24);
output(1, 42) <= input(25);
output(1, 43) <= input(26);
output(1, 44) <= input(27);
output(1, 45) <= input(28);
output(1, 46) <= input(29);
output(1, 47) <= input(30);
output(1, 48) <= input(33);
output(1, 49) <= input(16);
output(1, 50) <= input(17);
output(1, 51) <= input(18);
output(1, 52) <= input(19);
output(1, 53) <= input(20);
output(1, 54) <= input(21);
output(1, 55) <= input(22);
output(1, 56) <= input(23);
output(1, 57) <= input(24);
output(1, 58) <= input(25);
output(1, 59) <= input(26);
output(1, 60) <= input(27);
output(1, 61) <= input(28);
output(1, 62) <= input(29);
output(1, 63) <= input(30);
output(1, 64) <= input(33);
output(1, 65) <= input(16);
output(1, 66) <= input(17);
output(1, 67) <= input(18);
output(1, 68) <= input(19);
output(1, 69) <= input(20);
output(1, 70) <= input(21);
output(1, 71) <= input(22);
output(1, 72) <= input(23);
output(1, 73) <= input(24);
output(1, 74) <= input(25);
output(1, 75) <= input(26);
output(1, 76) <= input(27);
output(1, 77) <= input(28);
output(1, 78) <= input(29);
output(1, 79) <= input(30);
output(1, 80) <= input(34);
output(1, 81) <= input(32);
output(1, 82) <= input(0);
output(1, 83) <= input(1);
output(1, 84) <= input(2);
output(1, 85) <= input(3);
output(1, 86) <= input(4);
output(1, 87) <= input(5);
output(1, 88) <= input(6);
output(1, 89) <= input(7);
output(1, 90) <= input(8);
output(1, 91) <= input(9);
output(1, 92) <= input(10);
output(1, 93) <= input(11);
output(1, 94) <= input(12);
output(1, 95) <= input(13);
output(1, 96) <= input(34);
output(1, 97) <= input(32);
output(1, 98) <= input(0);
output(1, 99) <= input(1);
output(1, 100) <= input(2);
output(1, 101) <= input(3);
output(1, 102) <= input(4);
output(1, 103) <= input(5);
output(1, 104) <= input(6);
output(1, 105) <= input(7);
output(1, 106) <= input(8);
output(1, 107) <= input(9);
output(1, 108) <= input(10);
output(1, 109) <= input(11);
output(1, 110) <= input(12);
output(1, 111) <= input(13);
output(1, 112) <= input(34);
output(1, 113) <= input(32);
output(1, 114) <= input(0);
output(1, 115) <= input(1);
output(1, 116) <= input(2);
output(1, 117) <= input(3);
output(1, 118) <= input(4);
output(1, 119) <= input(5);
output(1, 120) <= input(6);
output(1, 121) <= input(7);
output(1, 122) <= input(8);
output(1, 123) <= input(9);
output(1, 124) <= input(10);
output(1, 125) <= input(11);
output(1, 126) <= input(12);
output(1, 127) <= input(13);
output(1, 128) <= input(35);
output(1, 129) <= input(33);
output(1, 130) <= input(16);
output(1, 131) <= input(17);
output(1, 132) <= input(18);
output(1, 133) <= input(19);
output(1, 134) <= input(20);
output(1, 135) <= input(21);
output(1, 136) <= input(22);
output(1, 137) <= input(23);
output(1, 138) <= input(24);
output(1, 139) <= input(25);
output(1, 140) <= input(26);
output(1, 141) <= input(27);
output(1, 142) <= input(28);
output(1, 143) <= input(29);
output(1, 144) <= input(35);
output(1, 145) <= input(33);
output(1, 146) <= input(16);
output(1, 147) <= input(17);
output(1, 148) <= input(18);
output(1, 149) <= input(19);
output(1, 150) <= input(20);
output(1, 151) <= input(21);
output(1, 152) <= input(22);
output(1, 153) <= input(23);
output(1, 154) <= input(24);
output(1, 155) <= input(25);
output(1, 156) <= input(26);
output(1, 157) <= input(27);
output(1, 158) <= input(28);
output(1, 159) <= input(29);
output(1, 160) <= input(36);
output(1, 161) <= input(34);
output(1, 162) <= input(32);
output(1, 163) <= input(0);
output(1, 164) <= input(1);
output(1, 165) <= input(2);
output(1, 166) <= input(3);
output(1, 167) <= input(4);
output(1, 168) <= input(5);
output(1, 169) <= input(6);
output(1, 170) <= input(7);
output(1, 171) <= input(8);
output(1, 172) <= input(9);
output(1, 173) <= input(10);
output(1, 174) <= input(11);
output(1, 175) <= input(12);
output(1, 176) <= input(36);
output(1, 177) <= input(34);
output(1, 178) <= input(32);
output(1, 179) <= input(0);
output(1, 180) <= input(1);
output(1, 181) <= input(2);
output(1, 182) <= input(3);
output(1, 183) <= input(4);
output(1, 184) <= input(5);
output(1, 185) <= input(6);
output(1, 186) <= input(7);
output(1, 187) <= input(8);
output(1, 188) <= input(9);
output(1, 189) <= input(10);
output(1, 190) <= input(11);
output(1, 191) <= input(12);
output(1, 192) <= input(36);
output(1, 193) <= input(34);
output(1, 194) <= input(32);
output(1, 195) <= input(0);
output(1, 196) <= input(1);
output(1, 197) <= input(2);
output(1, 198) <= input(3);
output(1, 199) <= input(4);
output(1, 200) <= input(5);
output(1, 201) <= input(6);
output(1, 202) <= input(7);
output(1, 203) <= input(8);
output(1, 204) <= input(9);
output(1, 205) <= input(10);
output(1, 206) <= input(11);
output(1, 207) <= input(12);
output(1, 208) <= input(37);
output(1, 209) <= input(35);
output(1, 210) <= input(33);
output(1, 211) <= input(16);
output(1, 212) <= input(17);
output(1, 213) <= input(18);
output(1, 214) <= input(19);
output(1, 215) <= input(20);
output(1, 216) <= input(21);
output(1, 217) <= input(22);
output(1, 218) <= input(23);
output(1, 219) <= input(24);
output(1, 220) <= input(25);
output(1, 221) <= input(26);
output(1, 222) <= input(27);
output(1, 223) <= input(28);
output(1, 224) <= input(37);
output(1, 225) <= input(35);
output(1, 226) <= input(33);
output(1, 227) <= input(16);
output(1, 228) <= input(17);
output(1, 229) <= input(18);
output(1, 230) <= input(19);
output(1, 231) <= input(20);
output(1, 232) <= input(21);
output(1, 233) <= input(22);
output(1, 234) <= input(23);
output(1, 235) <= input(24);
output(1, 236) <= input(25);
output(1, 237) <= input(26);
output(1, 238) <= input(27);
output(1, 239) <= input(28);
output(1, 240) <= input(37);
output(1, 241) <= input(35);
output(1, 242) <= input(33);
output(1, 243) <= input(16);
output(1, 244) <= input(17);
output(1, 245) <= input(18);
output(1, 246) <= input(19);
output(1, 247) <= input(20);
output(1, 248) <= input(21);
output(1, 249) <= input(22);
output(1, 250) <= input(23);
output(1, 251) <= input(24);
output(1, 252) <= input(25);
output(1, 253) <= input(26);
output(1, 254) <= input(27);
output(1, 255) <= input(28);
output(2, 0) <= input(34);
output(2, 1) <= input(32);
output(2, 2) <= input(0);
output(2, 3) <= input(1);
output(2, 4) <= input(2);
output(2, 5) <= input(3);
output(2, 6) <= input(4);
output(2, 7) <= input(5);
output(2, 8) <= input(6);
output(2, 9) <= input(7);
output(2, 10) <= input(8);
output(2, 11) <= input(9);
output(2, 12) <= input(10);
output(2, 13) <= input(11);
output(2, 14) <= input(12);
output(2, 15) <= input(13);
output(2, 16) <= input(34);
output(2, 17) <= input(32);
output(2, 18) <= input(0);
output(2, 19) <= input(1);
output(2, 20) <= input(2);
output(2, 21) <= input(3);
output(2, 22) <= input(4);
output(2, 23) <= input(5);
output(2, 24) <= input(6);
output(2, 25) <= input(7);
output(2, 26) <= input(8);
output(2, 27) <= input(9);
output(2, 28) <= input(10);
output(2, 29) <= input(11);
output(2, 30) <= input(12);
output(2, 31) <= input(13);
output(2, 32) <= input(35);
output(2, 33) <= input(33);
output(2, 34) <= input(16);
output(2, 35) <= input(17);
output(2, 36) <= input(18);
output(2, 37) <= input(19);
output(2, 38) <= input(20);
output(2, 39) <= input(21);
output(2, 40) <= input(22);
output(2, 41) <= input(23);
output(2, 42) <= input(24);
output(2, 43) <= input(25);
output(2, 44) <= input(26);
output(2, 45) <= input(27);
output(2, 46) <= input(28);
output(2, 47) <= input(29);
output(2, 48) <= input(35);
output(2, 49) <= input(33);
output(2, 50) <= input(16);
output(2, 51) <= input(17);
output(2, 52) <= input(18);
output(2, 53) <= input(19);
output(2, 54) <= input(20);
output(2, 55) <= input(21);
output(2, 56) <= input(22);
output(2, 57) <= input(23);
output(2, 58) <= input(24);
output(2, 59) <= input(25);
output(2, 60) <= input(26);
output(2, 61) <= input(27);
output(2, 62) <= input(28);
output(2, 63) <= input(29);
output(2, 64) <= input(36);
output(2, 65) <= input(34);
output(2, 66) <= input(32);
output(2, 67) <= input(0);
output(2, 68) <= input(1);
output(2, 69) <= input(2);
output(2, 70) <= input(3);
output(2, 71) <= input(4);
output(2, 72) <= input(5);
output(2, 73) <= input(6);
output(2, 74) <= input(7);
output(2, 75) <= input(8);
output(2, 76) <= input(9);
output(2, 77) <= input(10);
output(2, 78) <= input(11);
output(2, 79) <= input(12);
output(2, 80) <= input(36);
output(2, 81) <= input(34);
output(2, 82) <= input(32);
output(2, 83) <= input(0);
output(2, 84) <= input(1);
output(2, 85) <= input(2);
output(2, 86) <= input(3);
output(2, 87) <= input(4);
output(2, 88) <= input(5);
output(2, 89) <= input(6);
output(2, 90) <= input(7);
output(2, 91) <= input(8);
output(2, 92) <= input(9);
output(2, 93) <= input(10);
output(2, 94) <= input(11);
output(2, 95) <= input(12);
output(2, 96) <= input(37);
output(2, 97) <= input(35);
output(2, 98) <= input(33);
output(2, 99) <= input(16);
output(2, 100) <= input(17);
output(2, 101) <= input(18);
output(2, 102) <= input(19);
output(2, 103) <= input(20);
output(2, 104) <= input(21);
output(2, 105) <= input(22);
output(2, 106) <= input(23);
output(2, 107) <= input(24);
output(2, 108) <= input(25);
output(2, 109) <= input(26);
output(2, 110) <= input(27);
output(2, 111) <= input(28);
output(2, 112) <= input(37);
output(2, 113) <= input(35);
output(2, 114) <= input(33);
output(2, 115) <= input(16);
output(2, 116) <= input(17);
output(2, 117) <= input(18);
output(2, 118) <= input(19);
output(2, 119) <= input(20);
output(2, 120) <= input(21);
output(2, 121) <= input(22);
output(2, 122) <= input(23);
output(2, 123) <= input(24);
output(2, 124) <= input(25);
output(2, 125) <= input(26);
output(2, 126) <= input(27);
output(2, 127) <= input(28);
output(2, 128) <= input(38);
output(2, 129) <= input(36);
output(2, 130) <= input(34);
output(2, 131) <= input(32);
output(2, 132) <= input(0);
output(2, 133) <= input(1);
output(2, 134) <= input(2);
output(2, 135) <= input(3);
output(2, 136) <= input(4);
output(2, 137) <= input(5);
output(2, 138) <= input(6);
output(2, 139) <= input(7);
output(2, 140) <= input(8);
output(2, 141) <= input(9);
output(2, 142) <= input(10);
output(2, 143) <= input(11);
output(2, 144) <= input(38);
output(2, 145) <= input(36);
output(2, 146) <= input(34);
output(2, 147) <= input(32);
output(2, 148) <= input(0);
output(2, 149) <= input(1);
output(2, 150) <= input(2);
output(2, 151) <= input(3);
output(2, 152) <= input(4);
output(2, 153) <= input(5);
output(2, 154) <= input(6);
output(2, 155) <= input(7);
output(2, 156) <= input(8);
output(2, 157) <= input(9);
output(2, 158) <= input(10);
output(2, 159) <= input(11);
output(2, 160) <= input(39);
output(2, 161) <= input(37);
output(2, 162) <= input(35);
output(2, 163) <= input(33);
output(2, 164) <= input(16);
output(2, 165) <= input(17);
output(2, 166) <= input(18);
output(2, 167) <= input(19);
output(2, 168) <= input(20);
output(2, 169) <= input(21);
output(2, 170) <= input(22);
output(2, 171) <= input(23);
output(2, 172) <= input(24);
output(2, 173) <= input(25);
output(2, 174) <= input(26);
output(2, 175) <= input(27);
output(2, 176) <= input(39);
output(2, 177) <= input(37);
output(2, 178) <= input(35);
output(2, 179) <= input(33);
output(2, 180) <= input(16);
output(2, 181) <= input(17);
output(2, 182) <= input(18);
output(2, 183) <= input(19);
output(2, 184) <= input(20);
output(2, 185) <= input(21);
output(2, 186) <= input(22);
output(2, 187) <= input(23);
output(2, 188) <= input(24);
output(2, 189) <= input(25);
output(2, 190) <= input(26);
output(2, 191) <= input(27);
output(2, 192) <= input(40);
output(2, 193) <= input(38);
output(2, 194) <= input(36);
output(2, 195) <= input(34);
output(2, 196) <= input(32);
output(2, 197) <= input(0);
output(2, 198) <= input(1);
output(2, 199) <= input(2);
output(2, 200) <= input(3);
output(2, 201) <= input(4);
output(2, 202) <= input(5);
output(2, 203) <= input(6);
output(2, 204) <= input(7);
output(2, 205) <= input(8);
output(2, 206) <= input(9);
output(2, 207) <= input(10);
output(2, 208) <= input(40);
output(2, 209) <= input(38);
output(2, 210) <= input(36);
output(2, 211) <= input(34);
output(2, 212) <= input(32);
output(2, 213) <= input(0);
output(2, 214) <= input(1);
output(2, 215) <= input(2);
output(2, 216) <= input(3);
output(2, 217) <= input(4);
output(2, 218) <= input(5);
output(2, 219) <= input(6);
output(2, 220) <= input(7);
output(2, 221) <= input(8);
output(2, 222) <= input(9);
output(2, 223) <= input(10);
output(2, 224) <= input(41);
output(2, 225) <= input(39);
output(2, 226) <= input(37);
output(2, 227) <= input(35);
output(2, 228) <= input(33);
output(2, 229) <= input(16);
output(2, 230) <= input(17);
output(2, 231) <= input(18);
output(2, 232) <= input(19);
output(2, 233) <= input(20);
output(2, 234) <= input(21);
output(2, 235) <= input(22);
output(2, 236) <= input(23);
output(2, 237) <= input(24);
output(2, 238) <= input(25);
output(2, 239) <= input(26);
output(2, 240) <= input(41);
output(2, 241) <= input(39);
output(2, 242) <= input(37);
output(2, 243) <= input(35);
output(2, 244) <= input(33);
output(2, 245) <= input(16);
output(2, 246) <= input(17);
output(2, 247) <= input(18);
output(2, 248) <= input(19);
output(2, 249) <= input(20);
output(2, 250) <= input(21);
output(2, 251) <= input(22);
output(2, 252) <= input(23);
output(2, 253) <= input(24);
output(2, 254) <= input(25);
output(2, 255) <= input(26);
when "0100" =>
output(0, 0) <= input(0);
output(0, 1) <= input(1);
output(0, 2) <= input(2);
output(0, 3) <= input(3);
output(0, 4) <= input(4);
output(0, 5) <= input(5);
output(0, 6) <= input(6);
output(0, 7) <= input(7);
output(0, 8) <= input(8);
output(0, 9) <= input(9);
output(0, 10) <= input(10);
output(0, 11) <= input(11);
output(0, 12) <= input(12);
output(0, 13) <= input(13);
output(0, 14) <= input(14);
output(0, 15) <= input(15);
output(0, 16) <= input(16);
output(0, 17) <= input(17);
output(0, 18) <= input(18);
output(0, 19) <= input(19);
output(0, 20) <= input(20);
output(0, 21) <= input(21);
output(0, 22) <= input(22);
output(0, 23) <= input(23);
output(0, 24) <= input(24);
output(0, 25) <= input(25);
output(0, 26) <= input(26);
output(0, 27) <= input(27);
output(0, 28) <= input(28);
output(0, 29) <= input(29);
output(0, 30) <= input(30);
output(0, 31) <= input(31);
output(0, 32) <= input(16);
output(0, 33) <= input(17);
output(0, 34) <= input(18);
output(0, 35) <= input(19);
output(0, 36) <= input(20);
output(0, 37) <= input(21);
output(0, 38) <= input(22);
output(0, 39) <= input(23);
output(0, 40) <= input(24);
output(0, 41) <= input(25);
output(0, 42) <= input(26);
output(0, 43) <= input(27);
output(0, 44) <= input(28);
output(0, 45) <= input(29);
output(0, 46) <= input(30);
output(0, 47) <= input(31);
output(0, 48) <= input(32);
output(0, 49) <= input(0);
output(0, 50) <= input(1);
output(0, 51) <= input(2);
output(0, 52) <= input(3);
output(0, 53) <= input(4);
output(0, 54) <= input(5);
output(0, 55) <= input(6);
output(0, 56) <= input(7);
output(0, 57) <= input(8);
output(0, 58) <= input(9);
output(0, 59) <= input(10);
output(0, 60) <= input(11);
output(0, 61) <= input(12);
output(0, 62) <= input(13);
output(0, 63) <= input(14);
output(0, 64) <= input(33);
output(0, 65) <= input(16);
output(0, 66) <= input(17);
output(0, 67) <= input(18);
output(0, 68) <= input(19);
output(0, 69) <= input(20);
output(0, 70) <= input(21);
output(0, 71) <= input(22);
output(0, 72) <= input(23);
output(0, 73) <= input(24);
output(0, 74) <= input(25);
output(0, 75) <= input(26);
output(0, 76) <= input(27);
output(0, 77) <= input(28);
output(0, 78) <= input(29);
output(0, 79) <= input(30);
output(0, 80) <= input(33);
output(0, 81) <= input(16);
output(0, 82) <= input(17);
output(0, 83) <= input(18);
output(0, 84) <= input(19);
output(0, 85) <= input(20);
output(0, 86) <= input(21);
output(0, 87) <= input(22);
output(0, 88) <= input(23);
output(0, 89) <= input(24);
output(0, 90) <= input(25);
output(0, 91) <= input(26);
output(0, 92) <= input(27);
output(0, 93) <= input(28);
output(0, 94) <= input(29);
output(0, 95) <= input(30);
output(0, 96) <= input(34);
output(0, 97) <= input(32);
output(0, 98) <= input(0);
output(0, 99) <= input(1);
output(0, 100) <= input(2);
output(0, 101) <= input(3);
output(0, 102) <= input(4);
output(0, 103) <= input(5);
output(0, 104) <= input(6);
output(0, 105) <= input(7);
output(0, 106) <= input(8);
output(0, 107) <= input(9);
output(0, 108) <= input(10);
output(0, 109) <= input(11);
output(0, 110) <= input(12);
output(0, 111) <= input(13);
output(0, 112) <= input(34);
output(0, 113) <= input(32);
output(0, 114) <= input(0);
output(0, 115) <= input(1);
output(0, 116) <= input(2);
output(0, 117) <= input(3);
output(0, 118) <= input(4);
output(0, 119) <= input(5);
output(0, 120) <= input(6);
output(0, 121) <= input(7);
output(0, 122) <= input(8);
output(0, 123) <= input(9);
output(0, 124) <= input(10);
output(0, 125) <= input(11);
output(0, 126) <= input(12);
output(0, 127) <= input(13);
output(0, 128) <= input(35);
output(0, 129) <= input(33);
output(0, 130) <= input(16);
output(0, 131) <= input(17);
output(0, 132) <= input(18);
output(0, 133) <= input(19);
output(0, 134) <= input(20);
output(0, 135) <= input(21);
output(0, 136) <= input(22);
output(0, 137) <= input(23);
output(0, 138) <= input(24);
output(0, 139) <= input(25);
output(0, 140) <= input(26);
output(0, 141) <= input(27);
output(0, 142) <= input(28);
output(0, 143) <= input(29);
output(0, 144) <= input(36);
output(0, 145) <= input(34);
output(0, 146) <= input(32);
output(0, 147) <= input(0);
output(0, 148) <= input(1);
output(0, 149) <= input(2);
output(0, 150) <= input(3);
output(0, 151) <= input(4);
output(0, 152) <= input(5);
output(0, 153) <= input(6);
output(0, 154) <= input(7);
output(0, 155) <= input(8);
output(0, 156) <= input(9);
output(0, 157) <= input(10);
output(0, 158) <= input(11);
output(0, 159) <= input(12);
output(0, 160) <= input(36);
output(0, 161) <= input(34);
output(0, 162) <= input(32);
output(0, 163) <= input(0);
output(0, 164) <= input(1);
output(0, 165) <= input(2);
output(0, 166) <= input(3);
output(0, 167) <= input(4);
output(0, 168) <= input(5);
output(0, 169) <= input(6);
output(0, 170) <= input(7);
output(0, 171) <= input(8);
output(0, 172) <= input(9);
output(0, 173) <= input(10);
output(0, 174) <= input(11);
output(0, 175) <= input(12);
output(0, 176) <= input(37);
output(0, 177) <= input(35);
output(0, 178) <= input(33);
output(0, 179) <= input(16);
output(0, 180) <= input(17);
output(0, 181) <= input(18);
output(0, 182) <= input(19);
output(0, 183) <= input(20);
output(0, 184) <= input(21);
output(0, 185) <= input(22);
output(0, 186) <= input(23);
output(0, 187) <= input(24);
output(0, 188) <= input(25);
output(0, 189) <= input(26);
output(0, 190) <= input(27);
output(0, 191) <= input(28);
output(0, 192) <= input(38);
output(0, 193) <= input(36);
output(0, 194) <= input(34);
output(0, 195) <= input(32);
output(0, 196) <= input(0);
output(0, 197) <= input(1);
output(0, 198) <= input(2);
output(0, 199) <= input(3);
output(0, 200) <= input(4);
output(0, 201) <= input(5);
output(0, 202) <= input(6);
output(0, 203) <= input(7);
output(0, 204) <= input(8);
output(0, 205) <= input(9);
output(0, 206) <= input(10);
output(0, 207) <= input(11);
output(0, 208) <= input(38);
output(0, 209) <= input(36);
output(0, 210) <= input(34);
output(0, 211) <= input(32);
output(0, 212) <= input(0);
output(0, 213) <= input(1);
output(0, 214) <= input(2);
output(0, 215) <= input(3);
output(0, 216) <= input(4);
output(0, 217) <= input(5);
output(0, 218) <= input(6);
output(0, 219) <= input(7);
output(0, 220) <= input(8);
output(0, 221) <= input(9);
output(0, 222) <= input(10);
output(0, 223) <= input(11);
output(0, 224) <= input(39);
output(0, 225) <= input(37);
output(0, 226) <= input(35);
output(0, 227) <= input(33);
output(0, 228) <= input(16);
output(0, 229) <= input(17);
output(0, 230) <= input(18);
output(0, 231) <= input(19);
output(0, 232) <= input(20);
output(0, 233) <= input(21);
output(0, 234) <= input(22);
output(0, 235) <= input(23);
output(0, 236) <= input(24);
output(0, 237) <= input(25);
output(0, 238) <= input(26);
output(0, 239) <= input(27);
output(0, 240) <= input(39);
output(0, 241) <= input(37);
output(0, 242) <= input(35);
output(0, 243) <= input(33);
output(0, 244) <= input(16);
output(0, 245) <= input(17);
output(0, 246) <= input(18);
output(0, 247) <= input(19);
output(0, 248) <= input(20);
output(0, 249) <= input(21);
output(0, 250) <= input(22);
output(0, 251) <= input(23);
output(0, 252) <= input(24);
output(0, 253) <= input(25);
output(0, 254) <= input(26);
output(0, 255) <= input(27);
output(1, 0) <= input(32);
output(1, 1) <= input(0);
output(1, 2) <= input(1);
output(1, 3) <= input(2);
output(1, 4) <= input(3);
output(1, 5) <= input(4);
output(1, 6) <= input(5);
output(1, 7) <= input(6);
output(1, 8) <= input(7);
output(1, 9) <= input(8);
output(1, 10) <= input(9);
output(1, 11) <= input(10);
output(1, 12) <= input(11);
output(1, 13) <= input(12);
output(1, 14) <= input(13);
output(1, 15) <= input(14);
output(1, 16) <= input(33);
output(1, 17) <= input(16);
output(1, 18) <= input(17);
output(1, 19) <= input(18);
output(1, 20) <= input(19);
output(1, 21) <= input(20);
output(1, 22) <= input(21);
output(1, 23) <= input(22);
output(1, 24) <= input(23);
output(1, 25) <= input(24);
output(1, 26) <= input(25);
output(1, 27) <= input(26);
output(1, 28) <= input(27);
output(1, 29) <= input(28);
output(1, 30) <= input(29);
output(1, 31) <= input(30);
output(1, 32) <= input(34);
output(1, 33) <= input(32);
output(1, 34) <= input(0);
output(1, 35) <= input(1);
output(1, 36) <= input(2);
output(1, 37) <= input(3);
output(1, 38) <= input(4);
output(1, 39) <= input(5);
output(1, 40) <= input(6);
output(1, 41) <= input(7);
output(1, 42) <= input(8);
output(1, 43) <= input(9);
output(1, 44) <= input(10);
output(1, 45) <= input(11);
output(1, 46) <= input(12);
output(1, 47) <= input(13);
output(1, 48) <= input(34);
output(1, 49) <= input(32);
output(1, 50) <= input(0);
output(1, 51) <= input(1);
output(1, 52) <= input(2);
output(1, 53) <= input(3);
output(1, 54) <= input(4);
output(1, 55) <= input(5);
output(1, 56) <= input(6);
output(1, 57) <= input(7);
output(1, 58) <= input(8);
output(1, 59) <= input(9);
output(1, 60) <= input(10);
output(1, 61) <= input(11);
output(1, 62) <= input(12);
output(1, 63) <= input(13);
output(1, 64) <= input(35);
output(1, 65) <= input(33);
output(1, 66) <= input(16);
output(1, 67) <= input(17);
output(1, 68) <= input(18);
output(1, 69) <= input(19);
output(1, 70) <= input(20);
output(1, 71) <= input(21);
output(1, 72) <= input(22);
output(1, 73) <= input(23);
output(1, 74) <= input(24);
output(1, 75) <= input(25);
output(1, 76) <= input(26);
output(1, 77) <= input(27);
output(1, 78) <= input(28);
output(1, 79) <= input(29);
output(1, 80) <= input(36);
output(1, 81) <= input(34);
output(1, 82) <= input(32);
output(1, 83) <= input(0);
output(1, 84) <= input(1);
output(1, 85) <= input(2);
output(1, 86) <= input(3);
output(1, 87) <= input(4);
output(1, 88) <= input(5);
output(1, 89) <= input(6);
output(1, 90) <= input(7);
output(1, 91) <= input(8);
output(1, 92) <= input(9);
output(1, 93) <= input(10);
output(1, 94) <= input(11);
output(1, 95) <= input(12);
output(1, 96) <= input(37);
output(1, 97) <= input(35);
output(1, 98) <= input(33);
output(1, 99) <= input(16);
output(1, 100) <= input(17);
output(1, 101) <= input(18);
output(1, 102) <= input(19);
output(1, 103) <= input(20);
output(1, 104) <= input(21);
output(1, 105) <= input(22);
output(1, 106) <= input(23);
output(1, 107) <= input(24);
output(1, 108) <= input(25);
output(1, 109) <= input(26);
output(1, 110) <= input(27);
output(1, 111) <= input(28);
output(1, 112) <= input(37);
output(1, 113) <= input(35);
output(1, 114) <= input(33);
output(1, 115) <= input(16);
output(1, 116) <= input(17);
output(1, 117) <= input(18);
output(1, 118) <= input(19);
output(1, 119) <= input(20);
output(1, 120) <= input(21);
output(1, 121) <= input(22);
output(1, 122) <= input(23);
output(1, 123) <= input(24);
output(1, 124) <= input(25);
output(1, 125) <= input(26);
output(1, 126) <= input(27);
output(1, 127) <= input(28);
output(1, 128) <= input(38);
output(1, 129) <= input(36);
output(1, 130) <= input(34);
output(1, 131) <= input(32);
output(1, 132) <= input(0);
output(1, 133) <= input(1);
output(1, 134) <= input(2);
output(1, 135) <= input(3);
output(1, 136) <= input(4);
output(1, 137) <= input(5);
output(1, 138) <= input(6);
output(1, 139) <= input(7);
output(1, 140) <= input(8);
output(1, 141) <= input(9);
output(1, 142) <= input(10);
output(1, 143) <= input(11);
output(1, 144) <= input(39);
output(1, 145) <= input(37);
output(1, 146) <= input(35);
output(1, 147) <= input(33);
output(1, 148) <= input(16);
output(1, 149) <= input(17);
output(1, 150) <= input(18);
output(1, 151) <= input(19);
output(1, 152) <= input(20);
output(1, 153) <= input(21);
output(1, 154) <= input(22);
output(1, 155) <= input(23);
output(1, 156) <= input(24);
output(1, 157) <= input(25);
output(1, 158) <= input(26);
output(1, 159) <= input(27);
output(1, 160) <= input(40);
output(1, 161) <= input(38);
output(1, 162) <= input(36);
output(1, 163) <= input(34);
output(1, 164) <= input(32);
output(1, 165) <= input(0);
output(1, 166) <= input(1);
output(1, 167) <= input(2);
output(1, 168) <= input(3);
output(1, 169) <= input(4);
output(1, 170) <= input(5);
output(1, 171) <= input(6);
output(1, 172) <= input(7);
output(1, 173) <= input(8);
output(1, 174) <= input(9);
output(1, 175) <= input(10);
output(1, 176) <= input(40);
output(1, 177) <= input(38);
output(1, 178) <= input(36);
output(1, 179) <= input(34);
output(1, 180) <= input(32);
output(1, 181) <= input(0);
output(1, 182) <= input(1);
output(1, 183) <= input(2);
output(1, 184) <= input(3);
output(1, 185) <= input(4);
output(1, 186) <= input(5);
output(1, 187) <= input(6);
output(1, 188) <= input(7);
output(1, 189) <= input(8);
output(1, 190) <= input(9);
output(1, 191) <= input(10);
output(1, 192) <= input(41);
output(1, 193) <= input(39);
output(1, 194) <= input(37);
output(1, 195) <= input(35);
output(1, 196) <= input(33);
output(1, 197) <= input(16);
output(1, 198) <= input(17);
output(1, 199) <= input(18);
output(1, 200) <= input(19);
output(1, 201) <= input(20);
output(1, 202) <= input(21);
output(1, 203) <= input(22);
output(1, 204) <= input(23);
output(1, 205) <= input(24);
output(1, 206) <= input(25);
output(1, 207) <= input(26);
output(1, 208) <= input(42);
output(1, 209) <= input(40);
output(1, 210) <= input(38);
output(1, 211) <= input(36);
output(1, 212) <= input(34);
output(1, 213) <= input(32);
output(1, 214) <= input(0);
output(1, 215) <= input(1);
output(1, 216) <= input(2);
output(1, 217) <= input(3);
output(1, 218) <= input(4);
output(1, 219) <= input(5);
output(1, 220) <= input(6);
output(1, 221) <= input(7);
output(1, 222) <= input(8);
output(1, 223) <= input(9);
output(1, 224) <= input(43);
output(1, 225) <= input(41);
output(1, 226) <= input(39);
output(1, 227) <= input(37);
output(1, 228) <= input(35);
output(1, 229) <= input(33);
output(1, 230) <= input(16);
output(1, 231) <= input(17);
output(1, 232) <= input(18);
output(1, 233) <= input(19);
output(1, 234) <= input(20);
output(1, 235) <= input(21);
output(1, 236) <= input(22);
output(1, 237) <= input(23);
output(1, 238) <= input(24);
output(1, 239) <= input(25);
output(1, 240) <= input(43);
output(1, 241) <= input(41);
output(1, 242) <= input(39);
output(1, 243) <= input(37);
output(1, 244) <= input(35);
output(1, 245) <= input(33);
output(1, 246) <= input(16);
output(1, 247) <= input(17);
output(1, 248) <= input(18);
output(1, 249) <= input(19);
output(1, 250) <= input(20);
output(1, 251) <= input(21);
output(1, 252) <= input(22);
output(1, 253) <= input(23);
output(1, 254) <= input(24);
output(1, 255) <= input(25);
output(2, 0) <= input(34);
output(2, 1) <= input(32);
output(2, 2) <= input(0);
output(2, 3) <= input(1);
output(2, 4) <= input(2);
output(2, 5) <= input(3);
output(2, 6) <= input(4);
output(2, 7) <= input(5);
output(2, 8) <= input(6);
output(2, 9) <= input(7);
output(2, 10) <= input(8);
output(2, 11) <= input(9);
output(2, 12) <= input(10);
output(2, 13) <= input(11);
output(2, 14) <= input(12);
output(2, 15) <= input(13);
output(2, 16) <= input(35);
output(2, 17) <= input(33);
output(2, 18) <= input(16);
output(2, 19) <= input(17);
output(2, 20) <= input(18);
output(2, 21) <= input(19);
output(2, 22) <= input(20);
output(2, 23) <= input(21);
output(2, 24) <= input(22);
output(2, 25) <= input(23);
output(2, 26) <= input(24);
output(2, 27) <= input(25);
output(2, 28) <= input(26);
output(2, 29) <= input(27);
output(2, 30) <= input(28);
output(2, 31) <= input(29);
output(2, 32) <= input(36);
output(2, 33) <= input(34);
output(2, 34) <= input(32);
output(2, 35) <= input(0);
output(2, 36) <= input(1);
output(2, 37) <= input(2);
output(2, 38) <= input(3);
output(2, 39) <= input(4);
output(2, 40) <= input(5);
output(2, 41) <= input(6);
output(2, 42) <= input(7);
output(2, 43) <= input(8);
output(2, 44) <= input(9);
output(2, 45) <= input(10);
output(2, 46) <= input(11);
output(2, 47) <= input(12);
output(2, 48) <= input(37);
output(2, 49) <= input(35);
output(2, 50) <= input(33);
output(2, 51) <= input(16);
output(2, 52) <= input(17);
output(2, 53) <= input(18);
output(2, 54) <= input(19);
output(2, 55) <= input(20);
output(2, 56) <= input(21);
output(2, 57) <= input(22);
output(2, 58) <= input(23);
output(2, 59) <= input(24);
output(2, 60) <= input(25);
output(2, 61) <= input(26);
output(2, 62) <= input(27);
output(2, 63) <= input(28);
output(2, 64) <= input(38);
output(2, 65) <= input(36);
output(2, 66) <= input(34);
output(2, 67) <= input(32);
output(2, 68) <= input(0);
output(2, 69) <= input(1);
output(2, 70) <= input(2);
output(2, 71) <= input(3);
output(2, 72) <= input(4);
output(2, 73) <= input(5);
output(2, 74) <= input(6);
output(2, 75) <= input(7);
output(2, 76) <= input(8);
output(2, 77) <= input(9);
output(2, 78) <= input(10);
output(2, 79) <= input(11);
output(2, 80) <= input(39);
output(2, 81) <= input(37);
output(2, 82) <= input(35);
output(2, 83) <= input(33);
output(2, 84) <= input(16);
output(2, 85) <= input(17);
output(2, 86) <= input(18);
output(2, 87) <= input(19);
output(2, 88) <= input(20);
output(2, 89) <= input(21);
output(2, 90) <= input(22);
output(2, 91) <= input(23);
output(2, 92) <= input(24);
output(2, 93) <= input(25);
output(2, 94) <= input(26);
output(2, 95) <= input(27);
output(2, 96) <= input(40);
output(2, 97) <= input(38);
output(2, 98) <= input(36);
output(2, 99) <= input(34);
output(2, 100) <= input(32);
output(2, 101) <= input(0);
output(2, 102) <= input(1);
output(2, 103) <= input(2);
output(2, 104) <= input(3);
output(2, 105) <= input(4);
output(2, 106) <= input(5);
output(2, 107) <= input(6);
output(2, 108) <= input(7);
output(2, 109) <= input(8);
output(2, 110) <= input(9);
output(2, 111) <= input(10);
output(2, 112) <= input(40);
output(2, 113) <= input(38);
output(2, 114) <= input(36);
output(2, 115) <= input(34);
output(2, 116) <= input(32);
output(2, 117) <= input(0);
output(2, 118) <= input(1);
output(2, 119) <= input(2);
output(2, 120) <= input(3);
output(2, 121) <= input(4);
output(2, 122) <= input(5);
output(2, 123) <= input(6);
output(2, 124) <= input(7);
output(2, 125) <= input(8);
output(2, 126) <= input(9);
output(2, 127) <= input(10);
output(2, 128) <= input(41);
output(2, 129) <= input(39);
output(2, 130) <= input(37);
output(2, 131) <= input(35);
output(2, 132) <= input(33);
output(2, 133) <= input(16);
output(2, 134) <= input(17);
output(2, 135) <= input(18);
output(2, 136) <= input(19);
output(2, 137) <= input(20);
output(2, 138) <= input(21);
output(2, 139) <= input(22);
output(2, 140) <= input(23);
output(2, 141) <= input(24);
output(2, 142) <= input(25);
output(2, 143) <= input(26);
output(2, 144) <= input(42);
output(2, 145) <= input(40);
output(2, 146) <= input(38);
output(2, 147) <= input(36);
output(2, 148) <= input(34);
output(2, 149) <= input(32);
output(2, 150) <= input(0);
output(2, 151) <= input(1);
output(2, 152) <= input(2);
output(2, 153) <= input(3);
output(2, 154) <= input(4);
output(2, 155) <= input(5);
output(2, 156) <= input(6);
output(2, 157) <= input(7);
output(2, 158) <= input(8);
output(2, 159) <= input(9);
output(2, 160) <= input(43);
output(2, 161) <= input(41);
output(2, 162) <= input(39);
output(2, 163) <= input(37);
output(2, 164) <= input(35);
output(2, 165) <= input(33);
output(2, 166) <= input(16);
output(2, 167) <= input(17);
output(2, 168) <= input(18);
output(2, 169) <= input(19);
output(2, 170) <= input(20);
output(2, 171) <= input(21);
output(2, 172) <= input(22);
output(2, 173) <= input(23);
output(2, 174) <= input(24);
output(2, 175) <= input(25);
output(2, 176) <= input(44);
output(2, 177) <= input(42);
output(2, 178) <= input(40);
output(2, 179) <= input(38);
output(2, 180) <= input(36);
output(2, 181) <= input(34);
output(2, 182) <= input(32);
output(2, 183) <= input(0);
output(2, 184) <= input(1);
output(2, 185) <= input(2);
output(2, 186) <= input(3);
output(2, 187) <= input(4);
output(2, 188) <= input(5);
output(2, 189) <= input(6);
output(2, 190) <= input(7);
output(2, 191) <= input(8);
output(2, 192) <= input(45);
output(2, 193) <= input(43);
output(2, 194) <= input(41);
output(2, 195) <= input(39);
output(2, 196) <= input(37);
output(2, 197) <= input(35);
output(2, 198) <= input(33);
output(2, 199) <= input(16);
output(2, 200) <= input(17);
output(2, 201) <= input(18);
output(2, 202) <= input(19);
output(2, 203) <= input(20);
output(2, 204) <= input(21);
output(2, 205) <= input(22);
output(2, 206) <= input(23);
output(2, 207) <= input(24);
output(2, 208) <= input(46);
output(2, 209) <= input(44);
output(2, 210) <= input(42);
output(2, 211) <= input(40);
output(2, 212) <= input(38);
output(2, 213) <= input(36);
output(2, 214) <= input(34);
output(2, 215) <= input(32);
output(2, 216) <= input(0);
output(2, 217) <= input(1);
output(2, 218) <= input(2);
output(2, 219) <= input(3);
output(2, 220) <= input(4);
output(2, 221) <= input(5);
output(2, 222) <= input(6);
output(2, 223) <= input(7);
output(2, 224) <= input(47);
output(2, 225) <= input(45);
output(2, 226) <= input(43);
output(2, 227) <= input(41);
output(2, 228) <= input(39);
output(2, 229) <= input(37);
output(2, 230) <= input(35);
output(2, 231) <= input(33);
output(2, 232) <= input(16);
output(2, 233) <= input(17);
output(2, 234) <= input(18);
output(2, 235) <= input(19);
output(2, 236) <= input(20);
output(2, 237) <= input(21);
output(2, 238) <= input(22);
output(2, 239) <= input(23);
output(2, 240) <= input(47);
output(2, 241) <= input(45);
output(2, 242) <= input(43);
output(2, 243) <= input(41);
output(2, 244) <= input(39);
output(2, 245) <= input(37);
output(2, 246) <= input(35);
output(2, 247) <= input(33);
output(2, 248) <= input(16);
output(2, 249) <= input(17);
output(2, 250) <= input(18);
output(2, 251) <= input(19);
output(2, 252) <= input(20);
output(2, 253) <= input(21);
output(2, 254) <= input(22);
output(2, 255) <= input(23);
when "0101" =>
output(0, 0) <= input(0);
output(0, 1) <= input(1);
output(0, 2) <= input(2);
output(0, 3) <= input(3);
output(0, 4) <= input(4);
output(0, 5) <= input(5);
output(0, 6) <= input(6);
output(0, 7) <= input(7);
output(0, 8) <= input(8);
output(0, 9) <= input(9);
output(0, 10) <= input(10);
output(0, 11) <= input(11);
output(0, 12) <= input(12);
output(0, 13) <= input(13);
output(0, 14) <= input(14);
output(0, 15) <= input(15);
output(0, 16) <= input(16);
output(0, 17) <= input(17);
output(0, 18) <= input(18);
output(0, 19) <= input(19);
output(0, 20) <= input(20);
output(0, 21) <= input(21);
output(0, 22) <= input(22);
output(0, 23) <= input(23);
output(0, 24) <= input(24);
output(0, 25) <= input(25);
output(0, 26) <= input(26);
output(0, 27) <= input(27);
output(0, 28) <= input(28);
output(0, 29) <= input(29);
output(0, 30) <= input(30);
output(0, 31) <= input(31);
output(0, 32) <= input(32);
output(0, 33) <= input(0);
output(0, 34) <= input(1);
output(0, 35) <= input(2);
output(0, 36) <= input(3);
output(0, 37) <= input(4);
output(0, 38) <= input(5);
output(0, 39) <= input(6);
output(0, 40) <= input(7);
output(0, 41) <= input(8);
output(0, 42) <= input(9);
output(0, 43) <= input(10);
output(0, 44) <= input(11);
output(0, 45) <= input(12);
output(0, 46) <= input(13);
output(0, 47) <= input(14);
output(0, 48) <= input(33);
output(0, 49) <= input(16);
output(0, 50) <= input(17);
output(0, 51) <= input(18);
output(0, 52) <= input(19);
output(0, 53) <= input(20);
output(0, 54) <= input(21);
output(0, 55) <= input(22);
output(0, 56) <= input(23);
output(0, 57) <= input(24);
output(0, 58) <= input(25);
output(0, 59) <= input(26);
output(0, 60) <= input(27);
output(0, 61) <= input(28);
output(0, 62) <= input(29);
output(0, 63) <= input(30);
output(0, 64) <= input(34);
output(0, 65) <= input(32);
output(0, 66) <= input(0);
output(0, 67) <= input(1);
output(0, 68) <= input(2);
output(0, 69) <= input(3);
output(0, 70) <= input(4);
output(0, 71) <= input(5);
output(0, 72) <= input(6);
output(0, 73) <= input(7);
output(0, 74) <= input(8);
output(0, 75) <= input(9);
output(0, 76) <= input(10);
output(0, 77) <= input(11);
output(0, 78) <= input(12);
output(0, 79) <= input(13);
output(0, 80) <= input(35);
output(0, 81) <= input(33);
output(0, 82) <= input(16);
output(0, 83) <= input(17);
output(0, 84) <= input(18);
output(0, 85) <= input(19);
output(0, 86) <= input(20);
output(0, 87) <= input(21);
output(0, 88) <= input(22);
output(0, 89) <= input(23);
output(0, 90) <= input(24);
output(0, 91) <= input(25);
output(0, 92) <= input(26);
output(0, 93) <= input(27);
output(0, 94) <= input(28);
output(0, 95) <= input(29);
output(0, 96) <= input(36);
output(0, 97) <= input(34);
output(0, 98) <= input(32);
output(0, 99) <= input(0);
output(0, 100) <= input(1);
output(0, 101) <= input(2);
output(0, 102) <= input(3);
output(0, 103) <= input(4);
output(0, 104) <= input(5);
output(0, 105) <= input(6);
output(0, 106) <= input(7);
output(0, 107) <= input(8);
output(0, 108) <= input(9);
output(0, 109) <= input(10);
output(0, 110) <= input(11);
output(0, 111) <= input(12);
output(0, 112) <= input(37);
output(0, 113) <= input(35);
output(0, 114) <= input(33);
output(0, 115) <= input(16);
output(0, 116) <= input(17);
output(0, 117) <= input(18);
output(0, 118) <= input(19);
output(0, 119) <= input(20);
output(0, 120) <= input(21);
output(0, 121) <= input(22);
output(0, 122) <= input(23);
output(0, 123) <= input(24);
output(0, 124) <= input(25);
output(0, 125) <= input(26);
output(0, 126) <= input(27);
output(0, 127) <= input(28);
output(0, 128) <= input(38);
output(0, 129) <= input(36);
output(0, 130) <= input(34);
output(0, 131) <= input(32);
output(0, 132) <= input(0);
output(0, 133) <= input(1);
output(0, 134) <= input(2);
output(0, 135) <= input(3);
output(0, 136) <= input(4);
output(0, 137) <= input(5);
output(0, 138) <= input(6);
output(0, 139) <= input(7);
output(0, 140) <= input(8);
output(0, 141) <= input(9);
output(0, 142) <= input(10);
output(0, 143) <= input(11);
output(0, 144) <= input(39);
output(0, 145) <= input(37);
output(0, 146) <= input(35);
output(0, 147) <= input(33);
output(0, 148) <= input(16);
output(0, 149) <= input(17);
output(0, 150) <= input(18);
output(0, 151) <= input(19);
output(0, 152) <= input(20);
output(0, 153) <= input(21);
output(0, 154) <= input(22);
output(0, 155) <= input(23);
output(0, 156) <= input(24);
output(0, 157) <= input(25);
output(0, 158) <= input(26);
output(0, 159) <= input(27);
output(0, 160) <= input(40);
output(0, 161) <= input(38);
output(0, 162) <= input(36);
output(0, 163) <= input(34);
output(0, 164) <= input(32);
output(0, 165) <= input(0);
output(0, 166) <= input(1);
output(0, 167) <= input(2);
output(0, 168) <= input(3);
output(0, 169) <= input(4);
output(0, 170) <= input(5);
output(0, 171) <= input(6);
output(0, 172) <= input(7);
output(0, 173) <= input(8);
output(0, 174) <= input(9);
output(0, 175) <= input(10);
output(0, 176) <= input(41);
output(0, 177) <= input(39);
output(0, 178) <= input(37);
output(0, 179) <= input(35);
output(0, 180) <= input(33);
output(0, 181) <= input(16);
output(0, 182) <= input(17);
output(0, 183) <= input(18);
output(0, 184) <= input(19);
output(0, 185) <= input(20);
output(0, 186) <= input(21);
output(0, 187) <= input(22);
output(0, 188) <= input(23);
output(0, 189) <= input(24);
output(0, 190) <= input(25);
output(0, 191) <= input(26);
output(0, 192) <= input(42);
output(0, 193) <= input(40);
output(0, 194) <= input(38);
output(0, 195) <= input(36);
output(0, 196) <= input(34);
output(0, 197) <= input(32);
output(0, 198) <= input(0);
output(0, 199) <= input(1);
output(0, 200) <= input(2);
output(0, 201) <= input(3);
output(0, 202) <= input(4);
output(0, 203) <= input(5);
output(0, 204) <= input(6);
output(0, 205) <= input(7);
output(0, 206) <= input(8);
output(0, 207) <= input(9);
output(0, 208) <= input(43);
output(0, 209) <= input(41);
output(0, 210) <= input(39);
output(0, 211) <= input(37);
output(0, 212) <= input(35);
output(0, 213) <= input(33);
output(0, 214) <= input(16);
output(0, 215) <= input(17);
output(0, 216) <= input(18);
output(0, 217) <= input(19);
output(0, 218) <= input(20);
output(0, 219) <= input(21);
output(0, 220) <= input(22);
output(0, 221) <= input(23);
output(0, 222) <= input(24);
output(0, 223) <= input(25);
output(0, 224) <= input(44);
output(0, 225) <= input(42);
output(0, 226) <= input(40);
output(0, 227) <= input(38);
output(0, 228) <= input(36);
output(0, 229) <= input(34);
output(0, 230) <= input(32);
output(0, 231) <= input(0);
output(0, 232) <= input(1);
output(0, 233) <= input(2);
output(0, 234) <= input(3);
output(0, 235) <= input(4);
output(0, 236) <= input(5);
output(0, 237) <= input(6);
output(0, 238) <= input(7);
output(0, 239) <= input(8);
output(0, 240) <= input(45);
output(0, 241) <= input(43);
output(0, 242) <= input(41);
output(0, 243) <= input(39);
output(0, 244) <= input(37);
output(0, 245) <= input(35);
output(0, 246) <= input(33);
output(0, 247) <= input(16);
output(0, 248) <= input(17);
output(0, 249) <= input(18);
output(0, 250) <= input(19);
output(0, 251) <= input(20);
output(0, 252) <= input(21);
output(0, 253) <= input(22);
output(0, 254) <= input(23);
output(0, 255) <= input(24);
output(1, 0) <= input(33);
output(1, 1) <= input(16);
output(1, 2) <= input(17);
output(1, 3) <= input(18);
output(1, 4) <= input(19);
output(1, 5) <= input(20);
output(1, 6) <= input(21);
output(1, 7) <= input(22);
output(1, 8) <= input(23);
output(1, 9) <= input(24);
output(1, 10) <= input(25);
output(1, 11) <= input(26);
output(1, 12) <= input(27);
output(1, 13) <= input(28);
output(1, 14) <= input(29);
output(1, 15) <= input(30);
output(1, 16) <= input(34);
output(1, 17) <= input(32);
output(1, 18) <= input(0);
output(1, 19) <= input(1);
output(1, 20) <= input(2);
output(1, 21) <= input(3);
output(1, 22) <= input(4);
output(1, 23) <= input(5);
output(1, 24) <= input(6);
output(1, 25) <= input(7);
output(1, 26) <= input(8);
output(1, 27) <= input(9);
output(1, 28) <= input(10);
output(1, 29) <= input(11);
output(1, 30) <= input(12);
output(1, 31) <= input(13);
output(1, 32) <= input(35);
output(1, 33) <= input(33);
output(1, 34) <= input(16);
output(1, 35) <= input(17);
output(1, 36) <= input(18);
output(1, 37) <= input(19);
output(1, 38) <= input(20);
output(1, 39) <= input(21);
output(1, 40) <= input(22);
output(1, 41) <= input(23);
output(1, 42) <= input(24);
output(1, 43) <= input(25);
output(1, 44) <= input(26);
output(1, 45) <= input(27);
output(1, 46) <= input(28);
output(1, 47) <= input(29);
output(1, 48) <= input(36);
output(1, 49) <= input(34);
output(1, 50) <= input(32);
output(1, 51) <= input(0);
output(1, 52) <= input(1);
output(1, 53) <= input(2);
output(1, 54) <= input(3);
output(1, 55) <= input(4);
output(1, 56) <= input(5);
output(1, 57) <= input(6);
output(1, 58) <= input(7);
output(1, 59) <= input(8);
output(1, 60) <= input(9);
output(1, 61) <= input(10);
output(1, 62) <= input(11);
output(1, 63) <= input(12);
output(1, 64) <= input(37);
output(1, 65) <= input(35);
output(1, 66) <= input(33);
output(1, 67) <= input(16);
output(1, 68) <= input(17);
output(1, 69) <= input(18);
output(1, 70) <= input(19);
output(1, 71) <= input(20);
output(1, 72) <= input(21);
output(1, 73) <= input(22);
output(1, 74) <= input(23);
output(1, 75) <= input(24);
output(1, 76) <= input(25);
output(1, 77) <= input(26);
output(1, 78) <= input(27);
output(1, 79) <= input(28);
output(1, 80) <= input(38);
output(1, 81) <= input(36);
output(1, 82) <= input(34);
output(1, 83) <= input(32);
output(1, 84) <= input(0);
output(1, 85) <= input(1);
output(1, 86) <= input(2);
output(1, 87) <= input(3);
output(1, 88) <= input(4);
output(1, 89) <= input(5);
output(1, 90) <= input(6);
output(1, 91) <= input(7);
output(1, 92) <= input(8);
output(1, 93) <= input(9);
output(1, 94) <= input(10);
output(1, 95) <= input(11);
output(1, 96) <= input(39);
output(1, 97) <= input(37);
output(1, 98) <= input(35);
output(1, 99) <= input(33);
output(1, 100) <= input(16);
output(1, 101) <= input(17);
output(1, 102) <= input(18);
output(1, 103) <= input(19);
output(1, 104) <= input(20);
output(1, 105) <= input(21);
output(1, 106) <= input(22);
output(1, 107) <= input(23);
output(1, 108) <= input(24);
output(1, 109) <= input(25);
output(1, 110) <= input(26);
output(1, 111) <= input(27);
output(1, 112) <= input(40);
output(1, 113) <= input(38);
output(1, 114) <= input(36);
output(1, 115) <= input(34);
output(1, 116) <= input(32);
output(1, 117) <= input(0);
output(1, 118) <= input(1);
output(1, 119) <= input(2);
output(1, 120) <= input(3);
output(1, 121) <= input(4);
output(1, 122) <= input(5);
output(1, 123) <= input(6);
output(1, 124) <= input(7);
output(1, 125) <= input(8);
output(1, 126) <= input(9);
output(1, 127) <= input(10);
output(1, 128) <= input(42);
output(1, 129) <= input(40);
output(1, 130) <= input(38);
output(1, 131) <= input(36);
output(1, 132) <= input(34);
output(1, 133) <= input(32);
output(1, 134) <= input(0);
output(1, 135) <= input(1);
output(1, 136) <= input(2);
output(1, 137) <= input(3);
output(1, 138) <= input(4);
output(1, 139) <= input(5);
output(1, 140) <= input(6);
output(1, 141) <= input(7);
output(1, 142) <= input(8);
output(1, 143) <= input(9);
output(1, 144) <= input(43);
output(1, 145) <= input(41);
output(1, 146) <= input(39);
output(1, 147) <= input(37);
output(1, 148) <= input(35);
output(1, 149) <= input(33);
output(1, 150) <= input(16);
output(1, 151) <= input(17);
output(1, 152) <= input(18);
output(1, 153) <= input(19);
output(1, 154) <= input(20);
output(1, 155) <= input(21);
output(1, 156) <= input(22);
output(1, 157) <= input(23);
output(1, 158) <= input(24);
output(1, 159) <= input(25);
output(1, 160) <= input(44);
output(1, 161) <= input(42);
output(1, 162) <= input(40);
output(1, 163) <= input(38);
output(1, 164) <= input(36);
output(1, 165) <= input(34);
output(1, 166) <= input(32);
output(1, 167) <= input(0);
output(1, 168) <= input(1);
output(1, 169) <= input(2);
output(1, 170) <= input(3);
output(1, 171) <= input(4);
output(1, 172) <= input(5);
output(1, 173) <= input(6);
output(1, 174) <= input(7);
output(1, 175) <= input(8);
output(1, 176) <= input(45);
output(1, 177) <= input(43);
output(1, 178) <= input(41);
output(1, 179) <= input(39);
output(1, 180) <= input(37);
output(1, 181) <= input(35);
output(1, 182) <= input(33);
output(1, 183) <= input(16);
output(1, 184) <= input(17);
output(1, 185) <= input(18);
output(1, 186) <= input(19);
output(1, 187) <= input(20);
output(1, 188) <= input(21);
output(1, 189) <= input(22);
output(1, 190) <= input(23);
output(1, 191) <= input(24);
output(1, 192) <= input(46);
output(1, 193) <= input(44);
output(1, 194) <= input(42);
output(1, 195) <= input(40);
output(1, 196) <= input(38);
output(1, 197) <= input(36);
output(1, 198) <= input(34);
output(1, 199) <= input(32);
output(1, 200) <= input(0);
output(1, 201) <= input(1);
output(1, 202) <= input(2);
output(1, 203) <= input(3);
output(1, 204) <= input(4);
output(1, 205) <= input(5);
output(1, 206) <= input(6);
output(1, 207) <= input(7);
output(1, 208) <= input(47);
output(1, 209) <= input(45);
output(1, 210) <= input(43);
output(1, 211) <= input(41);
output(1, 212) <= input(39);
output(1, 213) <= input(37);
output(1, 214) <= input(35);
output(1, 215) <= input(33);
output(1, 216) <= input(16);
output(1, 217) <= input(17);
output(1, 218) <= input(18);
output(1, 219) <= input(19);
output(1, 220) <= input(20);
output(1, 221) <= input(21);
output(1, 222) <= input(22);
output(1, 223) <= input(23);
output(1, 224) <= input(48);
output(1, 225) <= input(46);
output(1, 226) <= input(44);
output(1, 227) <= input(42);
output(1, 228) <= input(40);
output(1, 229) <= input(38);
output(1, 230) <= input(36);
output(1, 231) <= input(34);
output(1, 232) <= input(32);
output(1, 233) <= input(0);
output(1, 234) <= input(1);
output(1, 235) <= input(2);
output(1, 236) <= input(3);
output(1, 237) <= input(4);
output(1, 238) <= input(5);
output(1, 239) <= input(6);
output(1, 240) <= input(49);
output(1, 241) <= input(47);
output(1, 242) <= input(45);
output(1, 243) <= input(43);
output(1, 244) <= input(41);
output(1, 245) <= input(39);
output(1, 246) <= input(37);
output(1, 247) <= input(35);
output(1, 248) <= input(33);
output(1, 249) <= input(16);
output(1, 250) <= input(17);
output(1, 251) <= input(18);
output(1, 252) <= input(19);
output(1, 253) <= input(20);
output(1, 254) <= input(21);
output(1, 255) <= input(22);
when "0110" =>
output(0, 0) <= input(0);
output(0, 1) <= input(1);
output(0, 2) <= input(2);
output(0, 3) <= input(3);
output(0, 4) <= input(4);
output(0, 5) <= input(5);
output(0, 6) <= input(6);
output(0, 7) <= input(7);
output(0, 8) <= input(8);
output(0, 9) <= input(9);
output(0, 10) <= input(10);
output(0, 11) <= input(11);
output(0, 12) <= input(12);
output(0, 13) <= input(13);
output(0, 14) <= input(14);
output(0, 15) <= input(15);
output(0, 16) <= input(16);
output(0, 17) <= input(17);
output(0, 18) <= input(18);
output(0, 19) <= input(19);
output(0, 20) <= input(20);
output(0, 21) <= input(21);
output(0, 22) <= input(22);
output(0, 23) <= input(23);
output(0, 24) <= input(24);
output(0, 25) <= input(25);
output(0, 26) <= input(26);
output(0, 27) <= input(27);
output(0, 28) <= input(28);
output(0, 29) <= input(29);
output(0, 30) <= input(30);
output(0, 31) <= input(31);
output(0, 32) <= input(32);
output(0, 33) <= input(0);
output(0, 34) <= input(1);
output(0, 35) <= input(2);
output(0, 36) <= input(3);
output(0, 37) <= input(4);
output(0, 38) <= input(5);
output(0, 39) <= input(6);
output(0, 40) <= input(7);
output(0, 41) <= input(8);
output(0, 42) <= input(9);
output(0, 43) <= input(10);
output(0, 44) <= input(11);
output(0, 45) <= input(12);
output(0, 46) <= input(13);
output(0, 47) <= input(14);
output(0, 48) <= input(33);
output(0, 49) <= input(16);
output(0, 50) <= input(17);
output(0, 51) <= input(18);
output(0, 52) <= input(19);
output(0, 53) <= input(20);
output(0, 54) <= input(21);
output(0, 55) <= input(22);
output(0, 56) <= input(23);
output(0, 57) <= input(24);
output(0, 58) <= input(25);
output(0, 59) <= input(26);
output(0, 60) <= input(27);
output(0, 61) <= input(28);
output(0, 62) <= input(29);
output(0, 63) <= input(30);
output(0, 64) <= input(34);
output(0, 65) <= input(33);
output(0, 66) <= input(16);
output(0, 67) <= input(17);
output(0, 68) <= input(18);
output(0, 69) <= input(19);
output(0, 70) <= input(20);
output(0, 71) <= input(21);
output(0, 72) <= input(22);
output(0, 73) <= input(23);
output(0, 74) <= input(24);
output(0, 75) <= input(25);
output(0, 76) <= input(26);
output(0, 77) <= input(27);
output(0, 78) <= input(28);
output(0, 79) <= input(29);
output(0, 80) <= input(35);
output(0, 81) <= input(36);
output(0, 82) <= input(32);
output(0, 83) <= input(0);
output(0, 84) <= input(1);
output(0, 85) <= input(2);
output(0, 86) <= input(3);
output(0, 87) <= input(4);
output(0, 88) <= input(5);
output(0, 89) <= input(6);
output(0, 90) <= input(7);
output(0, 91) <= input(8);
output(0, 92) <= input(9);
output(0, 93) <= input(10);
output(0, 94) <= input(11);
output(0, 95) <= input(12);
output(0, 96) <= input(37);
output(0, 97) <= input(34);
output(0, 98) <= input(33);
output(0, 99) <= input(16);
output(0, 100) <= input(17);
output(0, 101) <= input(18);
output(0, 102) <= input(19);
output(0, 103) <= input(20);
output(0, 104) <= input(21);
output(0, 105) <= input(22);
output(0, 106) <= input(23);
output(0, 107) <= input(24);
output(0, 108) <= input(25);
output(0, 109) <= input(26);
output(0, 110) <= input(27);
output(0, 111) <= input(28);
output(0, 112) <= input(38);
output(0, 113) <= input(35);
output(0, 114) <= input(36);
output(0, 115) <= input(32);
output(0, 116) <= input(0);
output(0, 117) <= input(1);
output(0, 118) <= input(2);
output(0, 119) <= input(3);
output(0, 120) <= input(4);
output(0, 121) <= input(5);
output(0, 122) <= input(6);
output(0, 123) <= input(7);
output(0, 124) <= input(8);
output(0, 125) <= input(9);
output(0, 126) <= input(10);
output(0, 127) <= input(11);
output(0, 128) <= input(39);
output(0, 129) <= input(38);
output(0, 130) <= input(35);
output(0, 131) <= input(36);
output(0, 132) <= input(32);
output(0, 133) <= input(0);
output(0, 134) <= input(1);
output(0, 135) <= input(2);
output(0, 136) <= input(3);
output(0, 137) <= input(4);
output(0, 138) <= input(5);
output(0, 139) <= input(6);
output(0, 140) <= input(7);
output(0, 141) <= input(8);
output(0, 142) <= input(9);
output(0, 143) <= input(10);
output(0, 144) <= input(40);
output(0, 145) <= input(41);
output(0, 146) <= input(37);
output(0, 147) <= input(34);
output(0, 148) <= input(33);
output(0, 149) <= input(16);
output(0, 150) <= input(17);
output(0, 151) <= input(18);
output(0, 152) <= input(19);
output(0, 153) <= input(20);
output(0, 154) <= input(21);
output(0, 155) <= input(22);
output(0, 156) <= input(23);
output(0, 157) <= input(24);
output(0, 158) <= input(25);
output(0, 159) <= input(26);
output(0, 160) <= input(42);
output(0, 161) <= input(39);
output(0, 162) <= input(38);
output(0, 163) <= input(35);
output(0, 164) <= input(36);
output(0, 165) <= input(32);
output(0, 166) <= input(0);
output(0, 167) <= input(1);
output(0, 168) <= input(2);
output(0, 169) <= input(3);
output(0, 170) <= input(4);
output(0, 171) <= input(5);
output(0, 172) <= input(6);
output(0, 173) <= input(7);
output(0, 174) <= input(8);
output(0, 175) <= input(9);
output(0, 176) <= input(43);
output(0, 177) <= input(40);
output(0, 178) <= input(41);
output(0, 179) <= input(37);
output(0, 180) <= input(34);
output(0, 181) <= input(33);
output(0, 182) <= input(16);
output(0, 183) <= input(17);
output(0, 184) <= input(18);
output(0, 185) <= input(19);
output(0, 186) <= input(20);
output(0, 187) <= input(21);
output(0, 188) <= input(22);
output(0, 189) <= input(23);
output(0, 190) <= input(24);
output(0, 191) <= input(25);
output(0, 192) <= input(44);
output(0, 193) <= input(43);
output(0, 194) <= input(40);
output(0, 195) <= input(41);
output(0, 196) <= input(37);
output(0, 197) <= input(34);
output(0, 198) <= input(33);
output(0, 199) <= input(16);
output(0, 200) <= input(17);
output(0, 201) <= input(18);
output(0, 202) <= input(19);
output(0, 203) <= input(20);
output(0, 204) <= input(21);
output(0, 205) <= input(22);
output(0, 206) <= input(23);
output(0, 207) <= input(24);
output(0, 208) <= input(45);
output(0, 209) <= input(46);
output(0, 210) <= input(42);
output(0, 211) <= input(39);
output(0, 212) <= input(38);
output(0, 213) <= input(35);
output(0, 214) <= input(36);
output(0, 215) <= input(32);
output(0, 216) <= input(0);
output(0, 217) <= input(1);
output(0, 218) <= input(2);
output(0, 219) <= input(3);
output(0, 220) <= input(4);
output(0, 221) <= input(5);
output(0, 222) <= input(6);
output(0, 223) <= input(7);
output(0, 224) <= input(47);
output(0, 225) <= input(44);
output(0, 226) <= input(43);
output(0, 227) <= input(40);
output(0, 228) <= input(41);
output(0, 229) <= input(37);
output(0, 230) <= input(34);
output(0, 231) <= input(33);
output(0, 232) <= input(16);
output(0, 233) <= input(17);
output(0, 234) <= input(18);
output(0, 235) <= input(19);
output(0, 236) <= input(20);
output(0, 237) <= input(21);
output(0, 238) <= input(22);
output(0, 239) <= input(23);
output(0, 240) <= input(48);
output(0, 241) <= input(45);
output(0, 242) <= input(46);
output(0, 243) <= input(42);
output(0, 244) <= input(39);
output(0, 245) <= input(38);
output(0, 246) <= input(35);
output(0, 247) <= input(36);
output(0, 248) <= input(32);
output(0, 249) <= input(0);
output(0, 250) <= input(1);
output(0, 251) <= input(2);
output(0, 252) <= input(3);
output(0, 253) <= input(4);
output(0, 254) <= input(5);
output(0, 255) <= input(6);
output(1, 0) <= input(33);
output(1, 1) <= input(16);
output(1, 2) <= input(17);
output(1, 3) <= input(18);
output(1, 4) <= input(19);
output(1, 5) <= input(20);
output(1, 6) <= input(21);
output(1, 7) <= input(22);
output(1, 8) <= input(23);
output(1, 9) <= input(24);
output(1, 10) <= input(25);
output(1, 11) <= input(26);
output(1, 12) <= input(27);
output(1, 13) <= input(28);
output(1, 14) <= input(29);
output(1, 15) <= input(30);
output(1, 16) <= input(36);
output(1, 17) <= input(32);
output(1, 18) <= input(0);
output(1, 19) <= input(1);
output(1, 20) <= input(2);
output(1, 21) <= input(3);
output(1, 22) <= input(4);
output(1, 23) <= input(5);
output(1, 24) <= input(6);
output(1, 25) <= input(7);
output(1, 26) <= input(8);
output(1, 27) <= input(9);
output(1, 28) <= input(10);
output(1, 29) <= input(11);
output(1, 30) <= input(12);
output(1, 31) <= input(13);
output(1, 32) <= input(35);
output(1, 33) <= input(36);
output(1, 34) <= input(32);
output(1, 35) <= input(0);
output(1, 36) <= input(1);
output(1, 37) <= input(2);
output(1, 38) <= input(3);
output(1, 39) <= input(4);
output(1, 40) <= input(5);
output(1, 41) <= input(6);
output(1, 42) <= input(7);
output(1, 43) <= input(8);
output(1, 44) <= input(9);
output(1, 45) <= input(10);
output(1, 46) <= input(11);
output(1, 47) <= input(12);
output(1, 48) <= input(37);
output(1, 49) <= input(34);
output(1, 50) <= input(33);
output(1, 51) <= input(16);
output(1, 52) <= input(17);
output(1, 53) <= input(18);
output(1, 54) <= input(19);
output(1, 55) <= input(20);
output(1, 56) <= input(21);
output(1, 57) <= input(22);
output(1, 58) <= input(23);
output(1, 59) <= input(24);
output(1, 60) <= input(25);
output(1, 61) <= input(26);
output(1, 62) <= input(27);
output(1, 63) <= input(28);
output(1, 64) <= input(41);
output(1, 65) <= input(37);
output(1, 66) <= input(34);
output(1, 67) <= input(33);
output(1, 68) <= input(16);
output(1, 69) <= input(17);
output(1, 70) <= input(18);
output(1, 71) <= input(19);
output(1, 72) <= input(20);
output(1, 73) <= input(21);
output(1, 74) <= input(22);
output(1, 75) <= input(23);
output(1, 76) <= input(24);
output(1, 77) <= input(25);
output(1, 78) <= input(26);
output(1, 79) <= input(27);
output(1, 80) <= input(39);
output(1, 81) <= input(38);
output(1, 82) <= input(35);
output(1, 83) <= input(36);
output(1, 84) <= input(32);
output(1, 85) <= input(0);
output(1, 86) <= input(1);
output(1, 87) <= input(2);
output(1, 88) <= input(3);
output(1, 89) <= input(4);
output(1, 90) <= input(5);
output(1, 91) <= input(6);
output(1, 92) <= input(7);
output(1, 93) <= input(8);
output(1, 94) <= input(9);
output(1, 95) <= input(10);
output(1, 96) <= input(42);
output(1, 97) <= input(39);
output(1, 98) <= input(38);
output(1, 99) <= input(35);
output(1, 100) <= input(36);
output(1, 101) <= input(32);
output(1, 102) <= input(0);
output(1, 103) <= input(1);
output(1, 104) <= input(2);
output(1, 105) <= input(3);
output(1, 106) <= input(4);
output(1, 107) <= input(5);
output(1, 108) <= input(6);
output(1, 109) <= input(7);
output(1, 110) <= input(8);
output(1, 111) <= input(9);
output(1, 112) <= input(43);
output(1, 113) <= input(40);
output(1, 114) <= input(41);
output(1, 115) <= input(37);
output(1, 116) <= input(34);
output(1, 117) <= input(33);
output(1, 118) <= input(16);
output(1, 119) <= input(17);
output(1, 120) <= input(18);
output(1, 121) <= input(19);
output(1, 122) <= input(20);
output(1, 123) <= input(21);
output(1, 124) <= input(22);
output(1, 125) <= input(23);
output(1, 126) <= input(24);
output(1, 127) <= input(25);
output(1, 128) <= input(46);
output(1, 129) <= input(42);
output(1, 130) <= input(39);
output(1, 131) <= input(38);
output(1, 132) <= input(35);
output(1, 133) <= input(36);
output(1, 134) <= input(32);
output(1, 135) <= input(0);
output(1, 136) <= input(1);
output(1, 137) <= input(2);
output(1, 138) <= input(3);
output(1, 139) <= input(4);
output(1, 140) <= input(5);
output(1, 141) <= input(6);
output(1, 142) <= input(7);
output(1, 143) <= input(8);
output(1, 144) <= input(45);
output(1, 145) <= input(46);
output(1, 146) <= input(42);
output(1, 147) <= input(39);
output(1, 148) <= input(38);
output(1, 149) <= input(35);
output(1, 150) <= input(36);
output(1, 151) <= input(32);
output(1, 152) <= input(0);
output(1, 153) <= input(1);
output(1, 154) <= input(2);
output(1, 155) <= input(3);
output(1, 156) <= input(4);
output(1, 157) <= input(5);
output(1, 158) <= input(6);
output(1, 159) <= input(7);
output(1, 160) <= input(47);
output(1, 161) <= input(44);
output(1, 162) <= input(43);
output(1, 163) <= input(40);
output(1, 164) <= input(41);
output(1, 165) <= input(37);
output(1, 166) <= input(34);
output(1, 167) <= input(33);
output(1, 168) <= input(16);
output(1, 169) <= input(17);
output(1, 170) <= input(18);
output(1, 171) <= input(19);
output(1, 172) <= input(20);
output(1, 173) <= input(21);
output(1, 174) <= input(22);
output(1, 175) <= input(23);
output(1, 176) <= input(49);
output(1, 177) <= input(47);
output(1, 178) <= input(44);
output(1, 179) <= input(43);
output(1, 180) <= input(40);
output(1, 181) <= input(41);
output(1, 182) <= input(37);
output(1, 183) <= input(34);
output(1, 184) <= input(33);
output(1, 185) <= input(16);
output(1, 186) <= input(17);
output(1, 187) <= input(18);
output(1, 188) <= input(19);
output(1, 189) <= input(20);
output(1, 190) <= input(21);
output(1, 191) <= input(22);
output(1, 192) <= input(50);
output(1, 193) <= input(48);
output(1, 194) <= input(45);
output(1, 195) <= input(46);
output(1, 196) <= input(42);
output(1, 197) <= input(39);
output(1, 198) <= input(38);
output(1, 199) <= input(35);
output(1, 200) <= input(36);
output(1, 201) <= input(32);
output(1, 202) <= input(0);
output(1, 203) <= input(1);
output(1, 204) <= input(2);
output(1, 205) <= input(3);
output(1, 206) <= input(4);
output(1, 207) <= input(5);
output(1, 208) <= input(51);
output(1, 209) <= input(50);
output(1, 210) <= input(48);
output(1, 211) <= input(45);
output(1, 212) <= input(46);
output(1, 213) <= input(42);
output(1, 214) <= input(39);
output(1, 215) <= input(38);
output(1, 216) <= input(35);
output(1, 217) <= input(36);
output(1, 218) <= input(32);
output(1, 219) <= input(0);
output(1, 220) <= input(1);
output(1, 221) <= input(2);
output(1, 222) <= input(3);
output(1, 223) <= input(4);
output(1, 224) <= input(52);
output(1, 225) <= input(53);
output(1, 226) <= input(49);
output(1, 227) <= input(47);
output(1, 228) <= input(44);
output(1, 229) <= input(43);
output(1, 230) <= input(40);
output(1, 231) <= input(41);
output(1, 232) <= input(37);
output(1, 233) <= input(34);
output(1, 234) <= input(33);
output(1, 235) <= input(16);
output(1, 236) <= input(17);
output(1, 237) <= input(18);
output(1, 238) <= input(19);
output(1, 239) <= input(20);
output(1, 240) <= input(54);
output(1, 241) <= input(51);
output(1, 242) <= input(50);
output(1, 243) <= input(48);
output(1, 244) <= input(45);
output(1, 245) <= input(46);
output(1, 246) <= input(42);
output(1, 247) <= input(39);
output(1, 248) <= input(38);
output(1, 249) <= input(35);
output(1, 250) <= input(36);
output(1, 251) <= input(32);
output(1, 252) <= input(0);
output(1, 253) <= input(1);
output(1, 254) <= input(2);
output(1, 255) <= input(3);
output(2, 0) <= input(35);
output(2, 1) <= input(36);
output(2, 2) <= input(32);
output(2, 3) <= input(0);
output(2, 4) <= input(1);
output(2, 5) <= input(2);
output(2, 6) <= input(3);
output(2, 7) <= input(4);
output(2, 8) <= input(5);
output(2, 9) <= input(6);
output(2, 10) <= input(7);
output(2, 11) <= input(8);
output(2, 12) <= input(9);
output(2, 13) <= input(10);
output(2, 14) <= input(11);
output(2, 15) <= input(12);
output(2, 16) <= input(38);
output(2, 17) <= input(35);
output(2, 18) <= input(36);
output(2, 19) <= input(32);
output(2, 20) <= input(0);
output(2, 21) <= input(1);
output(2, 22) <= input(2);
output(2, 23) <= input(3);
output(2, 24) <= input(4);
output(2, 25) <= input(5);
output(2, 26) <= input(6);
output(2, 27) <= input(7);
output(2, 28) <= input(8);
output(2, 29) <= input(9);
output(2, 30) <= input(10);
output(2, 31) <= input(11);
output(2, 32) <= input(41);
output(2, 33) <= input(37);
output(2, 34) <= input(34);
output(2, 35) <= input(33);
output(2, 36) <= input(16);
output(2, 37) <= input(17);
output(2, 38) <= input(18);
output(2, 39) <= input(19);
output(2, 40) <= input(20);
output(2, 41) <= input(21);
output(2, 42) <= input(22);
output(2, 43) <= input(23);
output(2, 44) <= input(24);
output(2, 45) <= input(25);
output(2, 46) <= input(26);
output(2, 47) <= input(27);
output(2, 48) <= input(40);
output(2, 49) <= input(41);
output(2, 50) <= input(37);
output(2, 51) <= input(34);
output(2, 52) <= input(33);
output(2, 53) <= input(16);
output(2, 54) <= input(17);
output(2, 55) <= input(18);
output(2, 56) <= input(19);
output(2, 57) <= input(20);
output(2, 58) <= input(21);
output(2, 59) <= input(22);
output(2, 60) <= input(23);
output(2, 61) <= input(24);
output(2, 62) <= input(25);
output(2, 63) <= input(26);
output(2, 64) <= input(43);
output(2, 65) <= input(40);
output(2, 66) <= input(41);
output(2, 67) <= input(37);
output(2, 68) <= input(34);
output(2, 69) <= input(33);
output(2, 70) <= input(16);
output(2, 71) <= input(17);
output(2, 72) <= input(18);
output(2, 73) <= input(19);
output(2, 74) <= input(20);
output(2, 75) <= input(21);
output(2, 76) <= input(22);
output(2, 77) <= input(23);
output(2, 78) <= input(24);
output(2, 79) <= input(25);
output(2, 80) <= input(46);
output(2, 81) <= input(42);
output(2, 82) <= input(39);
output(2, 83) <= input(38);
output(2, 84) <= input(35);
output(2, 85) <= input(36);
output(2, 86) <= input(32);
output(2, 87) <= input(0);
output(2, 88) <= input(1);
output(2, 89) <= input(2);
output(2, 90) <= input(3);
output(2, 91) <= input(4);
output(2, 92) <= input(5);
output(2, 93) <= input(6);
output(2, 94) <= input(7);
output(2, 95) <= input(8);
output(2, 96) <= input(45);
output(2, 97) <= input(46);
output(2, 98) <= input(42);
output(2, 99) <= input(39);
output(2, 100) <= input(38);
output(2, 101) <= input(35);
output(2, 102) <= input(36);
output(2, 103) <= input(32);
output(2, 104) <= input(0);
output(2, 105) <= input(1);
output(2, 106) <= input(2);
output(2, 107) <= input(3);
output(2, 108) <= input(4);
output(2, 109) <= input(5);
output(2, 110) <= input(6);
output(2, 111) <= input(7);
output(2, 112) <= input(47);
output(2, 113) <= input(44);
output(2, 114) <= input(43);
output(2, 115) <= input(40);
output(2, 116) <= input(41);
output(2, 117) <= input(37);
output(2, 118) <= input(34);
output(2, 119) <= input(33);
output(2, 120) <= input(16);
output(2, 121) <= input(17);
output(2, 122) <= input(18);
output(2, 123) <= input(19);
output(2, 124) <= input(20);
output(2, 125) <= input(21);
output(2, 126) <= input(22);
output(2, 127) <= input(23);
output(2, 128) <= input(49);
output(2, 129) <= input(47);
output(2, 130) <= input(44);
output(2, 131) <= input(43);
output(2, 132) <= input(40);
output(2, 133) <= input(41);
output(2, 134) <= input(37);
output(2, 135) <= input(34);
output(2, 136) <= input(33);
output(2, 137) <= input(16);
output(2, 138) <= input(17);
output(2, 139) <= input(18);
output(2, 140) <= input(19);
output(2, 141) <= input(20);
output(2, 142) <= input(21);
output(2, 143) <= input(22);
output(2, 144) <= input(53);
output(2, 145) <= input(49);
output(2, 146) <= input(47);
output(2, 147) <= input(44);
output(2, 148) <= input(43);
output(2, 149) <= input(40);
output(2, 150) <= input(41);
output(2, 151) <= input(37);
output(2, 152) <= input(34);
output(2, 153) <= input(33);
output(2, 154) <= input(16);
output(2, 155) <= input(17);
output(2, 156) <= input(18);
output(2, 157) <= input(19);
output(2, 158) <= input(20);
output(2, 159) <= input(21);
output(2, 160) <= input(51);
output(2, 161) <= input(50);
output(2, 162) <= input(48);
output(2, 163) <= input(45);
output(2, 164) <= input(46);
output(2, 165) <= input(42);
output(2, 166) <= input(39);
output(2, 167) <= input(38);
output(2, 168) <= input(35);
output(2, 169) <= input(36);
output(2, 170) <= input(32);
output(2, 171) <= input(0);
output(2, 172) <= input(1);
output(2, 173) <= input(2);
output(2, 174) <= input(3);
output(2, 175) <= input(4);
output(2, 176) <= input(54);
output(2, 177) <= input(51);
output(2, 178) <= input(50);
output(2, 179) <= input(48);
output(2, 180) <= input(45);
output(2, 181) <= input(46);
output(2, 182) <= input(42);
output(2, 183) <= input(39);
output(2, 184) <= input(38);
output(2, 185) <= input(35);
output(2, 186) <= input(36);
output(2, 187) <= input(32);
output(2, 188) <= input(0);
output(2, 189) <= input(1);
output(2, 190) <= input(2);
output(2, 191) <= input(3);
output(2, 192) <= input(55);
output(2, 193) <= input(54);
output(2, 194) <= input(51);
output(2, 195) <= input(50);
output(2, 196) <= input(48);
output(2, 197) <= input(45);
output(2, 198) <= input(46);
output(2, 199) <= input(42);
output(2, 200) <= input(39);
output(2, 201) <= input(38);
output(2, 202) <= input(35);
output(2, 203) <= input(36);
output(2, 204) <= input(32);
output(2, 205) <= input(0);
output(2, 206) <= input(1);
output(2, 207) <= input(2);
output(2, 208) <= input(56);
output(2, 209) <= input(57);
output(2, 210) <= input(52);
output(2, 211) <= input(53);
output(2, 212) <= input(49);
output(2, 213) <= input(47);
output(2, 214) <= input(44);
output(2, 215) <= input(43);
output(2, 216) <= input(40);
output(2, 217) <= input(41);
output(2, 218) <= input(37);
output(2, 219) <= input(34);
output(2, 220) <= input(33);
output(2, 221) <= input(16);
output(2, 222) <= input(17);
output(2, 223) <= input(18);
output(2, 224) <= input(58);
output(2, 225) <= input(56);
output(2, 226) <= input(57);
output(2, 227) <= input(52);
output(2, 228) <= input(53);
output(2, 229) <= input(49);
output(2, 230) <= input(47);
output(2, 231) <= input(44);
output(2, 232) <= input(43);
output(2, 233) <= input(40);
output(2, 234) <= input(41);
output(2, 235) <= input(37);
output(2, 236) <= input(34);
output(2, 237) <= input(33);
output(2, 238) <= input(16);
output(2, 239) <= input(17);
output(2, 240) <= input(59);
output(2, 241) <= input(60);
output(2, 242) <= input(55);
output(2, 243) <= input(54);
output(2, 244) <= input(51);
output(2, 245) <= input(50);
output(2, 246) <= input(48);
output(2, 247) <= input(45);
output(2, 248) <= input(46);
output(2, 249) <= input(42);
output(2, 250) <= input(39);
output(2, 251) <= input(38);
output(2, 252) <= input(35);
output(2, 253) <= input(36);
output(2, 254) <= input(32);
output(2, 255) <= input(0);
when "0111" =>
output(0, 0) <= input(0);
output(0, 1) <= input(1);
output(0, 2) <= input(2);
output(0, 3) <= input(3);
output(0, 4) <= input(4);
output(0, 5) <= input(5);
output(0, 6) <= input(6);
output(0, 7) <= input(7);
output(0, 8) <= input(8);
output(0, 9) <= input(9);
output(0, 10) <= input(10);
output(0, 11) <= input(11);
output(0, 12) <= input(12);
output(0, 13) <= input(13);
output(0, 14) <= input(14);
output(0, 15) <= input(15);
output(0, 16) <= input(16);
output(0, 17) <= input(0);
output(0, 18) <= input(1);
output(0, 19) <= input(2);
output(0, 20) <= input(3);
output(0, 21) <= input(4);
output(0, 22) <= input(5);
output(0, 23) <= input(6);
output(0, 24) <= input(7);
output(0, 25) <= input(8);
output(0, 26) <= input(9);
output(0, 27) <= input(10);
output(0, 28) <= input(11);
output(0, 29) <= input(12);
output(0, 30) <= input(13);
output(0, 31) <= input(14);
output(0, 32) <= input(17);
output(0, 33) <= input(16);
output(0, 34) <= input(0);
output(0, 35) <= input(1);
output(0, 36) <= input(2);
output(0, 37) <= input(3);
output(0, 38) <= input(4);
output(0, 39) <= input(5);
output(0, 40) <= input(6);
output(0, 41) <= input(7);
output(0, 42) <= input(8);
output(0, 43) <= input(9);
output(0, 44) <= input(10);
output(0, 45) <= input(11);
output(0, 46) <= input(12);
output(0, 47) <= input(13);
output(0, 48) <= input(18);
output(0, 49) <= input(17);
output(0, 50) <= input(16);
output(0, 51) <= input(0);
output(0, 52) <= input(1);
output(0, 53) <= input(2);
output(0, 54) <= input(3);
output(0, 55) <= input(4);
output(0, 56) <= input(5);
output(0, 57) <= input(6);
output(0, 58) <= input(7);
output(0, 59) <= input(8);
output(0, 60) <= input(9);
output(0, 61) <= input(10);
output(0, 62) <= input(11);
output(0, 63) <= input(12);
output(0, 64) <= input(19);
output(0, 65) <= input(18);
output(0, 66) <= input(17);
output(0, 67) <= input(16);
output(0, 68) <= input(0);
output(0, 69) <= input(1);
output(0, 70) <= input(2);
output(0, 71) <= input(3);
output(0, 72) <= input(4);
output(0, 73) <= input(5);
output(0, 74) <= input(6);
output(0, 75) <= input(7);
output(0, 76) <= input(8);
output(0, 77) <= input(9);
output(0, 78) <= input(10);
output(0, 79) <= input(11);
output(0, 80) <= input(20);
output(0, 81) <= input(21);
output(0, 82) <= input(22);
output(0, 83) <= input(23);
output(0, 84) <= input(24);
output(0, 85) <= input(25);
output(0, 86) <= input(26);
output(0, 87) <= input(27);
output(0, 88) <= input(28);
output(0, 89) <= input(29);
output(0, 90) <= input(30);
output(0, 91) <= input(31);
output(0, 92) <= input(32);
output(0, 93) <= input(33);
output(0, 94) <= input(34);
output(0, 95) <= input(35);
output(0, 96) <= input(36);
output(0, 97) <= input(20);
output(0, 98) <= input(21);
output(0, 99) <= input(22);
output(0, 100) <= input(23);
output(0, 101) <= input(24);
output(0, 102) <= input(25);
output(0, 103) <= input(26);
output(0, 104) <= input(27);
output(0, 105) <= input(28);
output(0, 106) <= input(29);
output(0, 107) <= input(30);
output(0, 108) <= input(31);
output(0, 109) <= input(32);
output(0, 110) <= input(33);
output(0, 111) <= input(34);
output(0, 112) <= input(37);
output(0, 113) <= input(36);
output(0, 114) <= input(20);
output(0, 115) <= input(21);
output(0, 116) <= input(22);
output(0, 117) <= input(23);
output(0, 118) <= input(24);
output(0, 119) <= input(25);
output(0, 120) <= input(26);
output(0, 121) <= input(27);
output(0, 122) <= input(28);
output(0, 123) <= input(29);
output(0, 124) <= input(30);
output(0, 125) <= input(31);
output(0, 126) <= input(32);
output(0, 127) <= input(33);
output(0, 128) <= input(38);
output(0, 129) <= input(37);
output(0, 130) <= input(36);
output(0, 131) <= input(20);
output(0, 132) <= input(21);
output(0, 133) <= input(22);
output(0, 134) <= input(23);
output(0, 135) <= input(24);
output(0, 136) <= input(25);
output(0, 137) <= input(26);
output(0, 138) <= input(27);
output(0, 139) <= input(28);
output(0, 140) <= input(29);
output(0, 141) <= input(30);
output(0, 142) <= input(31);
output(0, 143) <= input(32);
output(0, 144) <= input(39);
output(0, 145) <= input(38);
output(0, 146) <= input(37);
output(0, 147) <= input(36);
output(0, 148) <= input(20);
output(0, 149) <= input(21);
output(0, 150) <= input(22);
output(0, 151) <= input(23);
output(0, 152) <= input(24);
output(0, 153) <= input(25);
output(0, 154) <= input(26);
output(0, 155) <= input(27);
output(0, 156) <= input(28);
output(0, 157) <= input(29);
output(0, 158) <= input(30);
output(0, 159) <= input(31);
output(0, 160) <= input(40);
output(0, 161) <= input(41);
output(0, 162) <= input(42);
output(0, 163) <= input(43);
output(0, 164) <= input(44);
output(0, 165) <= input(19);
output(0, 166) <= input(18);
output(0, 167) <= input(17);
output(0, 168) <= input(16);
output(0, 169) <= input(0);
output(0, 170) <= input(1);
output(0, 171) <= input(2);
output(0, 172) <= input(3);
output(0, 173) <= input(4);
output(0, 174) <= input(5);
output(0, 175) <= input(6);
output(0, 176) <= input(45);
output(0, 177) <= input(40);
output(0, 178) <= input(41);
output(0, 179) <= input(42);
output(0, 180) <= input(43);
output(0, 181) <= input(44);
output(0, 182) <= input(19);
output(0, 183) <= input(18);
output(0, 184) <= input(17);
output(0, 185) <= input(16);
output(0, 186) <= input(0);
output(0, 187) <= input(1);
output(0, 188) <= input(2);
output(0, 189) <= input(3);
output(0, 190) <= input(4);
output(0, 191) <= input(5);
output(0, 192) <= input(46);
output(0, 193) <= input(45);
output(0, 194) <= input(40);
output(0, 195) <= input(41);
output(0, 196) <= input(42);
output(0, 197) <= input(43);
output(0, 198) <= input(44);
output(0, 199) <= input(19);
output(0, 200) <= input(18);
output(0, 201) <= input(17);
output(0, 202) <= input(16);
output(0, 203) <= input(0);
output(0, 204) <= input(1);
output(0, 205) <= input(2);
output(0, 206) <= input(3);
output(0, 207) <= input(4);
output(0, 208) <= input(47);
output(0, 209) <= input(46);
output(0, 210) <= input(45);
output(0, 211) <= input(40);
output(0, 212) <= input(41);
output(0, 213) <= input(42);
output(0, 214) <= input(43);
output(0, 215) <= input(44);
output(0, 216) <= input(19);
output(0, 217) <= input(18);
output(0, 218) <= input(17);
output(0, 219) <= input(16);
output(0, 220) <= input(0);
output(0, 221) <= input(1);
output(0, 222) <= input(2);
output(0, 223) <= input(3);
output(0, 224) <= input(48);
output(0, 225) <= input(47);
output(0, 226) <= input(46);
output(0, 227) <= input(45);
output(0, 228) <= input(40);
output(0, 229) <= input(41);
output(0, 230) <= input(42);
output(0, 231) <= input(43);
output(0, 232) <= input(44);
output(0, 233) <= input(19);
output(0, 234) <= input(18);
output(0, 235) <= input(17);
output(0, 236) <= input(16);
output(0, 237) <= input(0);
output(0, 238) <= input(1);
output(0, 239) <= input(2);
output(0, 240) <= input(49);
output(0, 241) <= input(50);
output(0, 242) <= input(51);
output(0, 243) <= input(52);
output(0, 244) <= input(53);
output(0, 245) <= input(39);
output(0, 246) <= input(38);
output(0, 247) <= input(37);
output(0, 248) <= input(36);
output(0, 249) <= input(20);
output(0, 250) <= input(21);
output(0, 251) <= input(22);
output(0, 252) <= input(23);
output(0, 253) <= input(24);
output(0, 254) <= input(25);
output(0, 255) <= input(26);
output(1, 0) <= input(54);
output(1, 1) <= input(55);
output(1, 2) <= input(56);
output(1, 3) <= input(57);
output(1, 4) <= input(58);
output(1, 5) <= input(59);
output(1, 6) <= input(60);
output(1, 7) <= input(61);
output(1, 8) <= input(62);
output(1, 9) <= input(63);
output(1, 10) <= input(64);
output(1, 11) <= input(65);
output(1, 12) <= input(66);
output(1, 13) <= input(67);
output(1, 14) <= input(68);
output(1, 15) <= input(69);
output(1, 16) <= input(70);
output(1, 17) <= input(54);
output(1, 18) <= input(55);
output(1, 19) <= input(56);
output(1, 20) <= input(57);
output(1, 21) <= input(58);
output(1, 22) <= input(59);
output(1, 23) <= input(60);
output(1, 24) <= input(61);
output(1, 25) <= input(62);
output(1, 26) <= input(63);
output(1, 27) <= input(64);
output(1, 28) <= input(65);
output(1, 29) <= input(66);
output(1, 30) <= input(67);
output(1, 31) <= input(68);
output(1, 32) <= input(71);
output(1, 33) <= input(70);
output(1, 34) <= input(54);
output(1, 35) <= input(55);
output(1, 36) <= input(56);
output(1, 37) <= input(57);
output(1, 38) <= input(58);
output(1, 39) <= input(59);
output(1, 40) <= input(60);
output(1, 41) <= input(61);
output(1, 42) <= input(62);
output(1, 43) <= input(63);
output(1, 44) <= input(64);
output(1, 45) <= input(65);
output(1, 46) <= input(66);
output(1, 47) <= input(67);
output(1, 48) <= input(72);
output(1, 49) <= input(71);
output(1, 50) <= input(70);
output(1, 51) <= input(54);
output(1, 52) <= input(55);
output(1, 53) <= input(56);
output(1, 54) <= input(57);
output(1, 55) <= input(58);
output(1, 56) <= input(59);
output(1, 57) <= input(60);
output(1, 58) <= input(61);
output(1, 59) <= input(62);
output(1, 60) <= input(63);
output(1, 61) <= input(64);
output(1, 62) <= input(65);
output(1, 63) <= input(66);
output(1, 64) <= input(73);
output(1, 65) <= input(72);
output(1, 66) <= input(71);
output(1, 67) <= input(70);
output(1, 68) <= input(54);
output(1, 69) <= input(55);
output(1, 70) <= input(56);
output(1, 71) <= input(57);
output(1, 72) <= input(58);
output(1, 73) <= input(59);
output(1, 74) <= input(60);
output(1, 75) <= input(61);
output(1, 76) <= input(62);
output(1, 77) <= input(63);
output(1, 78) <= input(64);
output(1, 79) <= input(65);
output(1, 80) <= input(74);
output(1, 81) <= input(73);
output(1, 82) <= input(72);
output(1, 83) <= input(71);
output(1, 84) <= input(70);
output(1, 85) <= input(54);
output(1, 86) <= input(55);
output(1, 87) <= input(56);
output(1, 88) <= input(57);
output(1, 89) <= input(58);
output(1, 90) <= input(59);
output(1, 91) <= input(60);
output(1, 92) <= input(61);
output(1, 93) <= input(62);
output(1, 94) <= input(63);
output(1, 95) <= input(64);
output(1, 96) <= input(75);
output(1, 97) <= input(74);
output(1, 98) <= input(73);
output(1, 99) <= input(72);
output(1, 100) <= input(71);
output(1, 101) <= input(70);
output(1, 102) <= input(54);
output(1, 103) <= input(55);
output(1, 104) <= input(56);
output(1, 105) <= input(57);
output(1, 106) <= input(58);
output(1, 107) <= input(59);
output(1, 108) <= input(60);
output(1, 109) <= input(61);
output(1, 110) <= input(62);
output(1, 111) <= input(63);
output(1, 112) <= input(76);
output(1, 113) <= input(75);
output(1, 114) <= input(74);
output(1, 115) <= input(73);
output(1, 116) <= input(72);
output(1, 117) <= input(71);
output(1, 118) <= input(70);
output(1, 119) <= input(54);
output(1, 120) <= input(55);
output(1, 121) <= input(56);
output(1, 122) <= input(57);
output(1, 123) <= input(58);
output(1, 124) <= input(59);
output(1, 125) <= input(60);
output(1, 126) <= input(61);
output(1, 127) <= input(62);
output(1, 128) <= input(77);
output(1, 129) <= input(76);
output(1, 130) <= input(75);
output(1, 131) <= input(74);
output(1, 132) <= input(73);
output(1, 133) <= input(72);
output(1, 134) <= input(71);
output(1, 135) <= input(70);
output(1, 136) <= input(54);
output(1, 137) <= input(55);
output(1, 138) <= input(56);
output(1, 139) <= input(57);
output(1, 140) <= input(58);
output(1, 141) <= input(59);
output(1, 142) <= input(60);
output(1, 143) <= input(61);
output(1, 144) <= input(78);
output(1, 145) <= input(77);
output(1, 146) <= input(76);
output(1, 147) <= input(75);
output(1, 148) <= input(74);
output(1, 149) <= input(73);
output(1, 150) <= input(72);
output(1, 151) <= input(71);
output(1, 152) <= input(70);
output(1, 153) <= input(54);
output(1, 154) <= input(55);
output(1, 155) <= input(56);
output(1, 156) <= input(57);
output(1, 157) <= input(58);
output(1, 158) <= input(59);
output(1, 159) <= input(60);
output(1, 160) <= input(79);
output(1, 161) <= input(78);
output(1, 162) <= input(77);
output(1, 163) <= input(76);
output(1, 164) <= input(75);
output(1, 165) <= input(74);
output(1, 166) <= input(73);
output(1, 167) <= input(72);
output(1, 168) <= input(71);
output(1, 169) <= input(70);
output(1, 170) <= input(54);
output(1, 171) <= input(55);
output(1, 172) <= input(56);
output(1, 173) <= input(57);
output(1, 174) <= input(58);
output(1, 175) <= input(59);
output(1, 176) <= input(80);
output(1, 177) <= input(79);
output(1, 178) <= input(78);
output(1, 179) <= input(77);
output(1, 180) <= input(76);
output(1, 181) <= input(75);
output(1, 182) <= input(74);
output(1, 183) <= input(73);
output(1, 184) <= input(72);
output(1, 185) <= input(71);
output(1, 186) <= input(70);
output(1, 187) <= input(54);
output(1, 188) <= input(55);
output(1, 189) <= input(56);
output(1, 190) <= input(57);
output(1, 191) <= input(58);
output(1, 192) <= input(81);
output(1, 193) <= input(80);
output(1, 194) <= input(79);
output(1, 195) <= input(78);
output(1, 196) <= input(77);
output(1, 197) <= input(76);
output(1, 198) <= input(75);
output(1, 199) <= input(74);
output(1, 200) <= input(73);
output(1, 201) <= input(72);
output(1, 202) <= input(71);
output(1, 203) <= input(70);
output(1, 204) <= input(54);
output(1, 205) <= input(55);
output(1, 206) <= input(56);
output(1, 207) <= input(57);
output(1, 208) <= input(82);
output(1, 209) <= input(81);
output(1, 210) <= input(80);
output(1, 211) <= input(79);
output(1, 212) <= input(78);
output(1, 213) <= input(77);
output(1, 214) <= input(76);
output(1, 215) <= input(75);
output(1, 216) <= input(74);
output(1, 217) <= input(73);
output(1, 218) <= input(72);
output(1, 219) <= input(71);
output(1, 220) <= input(70);
output(1, 221) <= input(54);
output(1, 222) <= input(55);
output(1, 223) <= input(56);
output(1, 224) <= input(83);
output(1, 225) <= input(82);
output(1, 226) <= input(81);
output(1, 227) <= input(80);
output(1, 228) <= input(79);
output(1, 229) <= input(78);
output(1, 230) <= input(77);
output(1, 231) <= input(76);
output(1, 232) <= input(75);
output(1, 233) <= input(74);
output(1, 234) <= input(73);
output(1, 235) <= input(72);
output(1, 236) <= input(71);
output(1, 237) <= input(70);
output(1, 238) <= input(54);
output(1, 239) <= input(55);
output(1, 240) <= input(84);
output(1, 241) <= input(83);
output(1, 242) <= input(82);
output(1, 243) <= input(81);
output(1, 244) <= input(80);
output(1, 245) <= input(79);
output(1, 246) <= input(78);
output(1, 247) <= input(77);
output(1, 248) <= input(76);
output(1, 249) <= input(75);
output(1, 250) <= input(74);
output(1, 251) <= input(73);
output(1, 252) <= input(72);
output(1, 253) <= input(71);
output(1, 254) <= input(70);
output(1, 255) <= input(54);
when "1000" =>
output(0, 0) <= input(0);
output(0, 1) <= input(1);
output(0, 2) <= input(2);
output(0, 3) <= input(3);
output(0, 4) <= input(4);
output(0, 5) <= input(5);
output(0, 6) <= input(6);
output(0, 7) <= input(7);
output(0, 8) <= input(8);
output(0, 9) <= input(9);
output(0, 10) <= input(10);
output(0, 11) <= input(11);
output(0, 12) <= input(12);
output(0, 13) <= input(13);
output(0, 14) <= input(14);
output(0, 15) <= input(15);
output(0, 16) <= input(16);
output(0, 17) <= input(0);
output(0, 18) <= input(1);
output(0, 19) <= input(2);
output(0, 20) <= input(3);
output(0, 21) <= input(4);
output(0, 22) <= input(5);
output(0, 23) <= input(6);
output(0, 24) <= input(7);
output(0, 25) <= input(8);
output(0, 26) <= input(9);
output(0, 27) <= input(10);
output(0, 28) <= input(11);
output(0, 29) <= input(12);
output(0, 30) <= input(13);
output(0, 31) <= input(14);
output(0, 32) <= input(17);
output(0, 33) <= input(16);
output(0, 34) <= input(0);
output(0, 35) <= input(1);
output(0, 36) <= input(2);
output(0, 37) <= input(3);
output(0, 38) <= input(4);
output(0, 39) <= input(5);
output(0, 40) <= input(6);
output(0, 41) <= input(7);
output(0, 42) <= input(8);
output(0, 43) <= input(9);
output(0, 44) <= input(10);
output(0, 45) <= input(11);
output(0, 46) <= input(12);
output(0, 47) <= input(13);
output(0, 48) <= input(18);
output(0, 49) <= input(17);
output(0, 50) <= input(16);
output(0, 51) <= input(0);
output(0, 52) <= input(1);
output(0, 53) <= input(2);
output(0, 54) <= input(3);
output(0, 55) <= input(4);
output(0, 56) <= input(5);
output(0, 57) <= input(6);
output(0, 58) <= input(7);
output(0, 59) <= input(8);
output(0, 60) <= input(9);
output(0, 61) <= input(10);
output(0, 62) <= input(11);
output(0, 63) <= input(12);
output(0, 64) <= input(19);
output(0, 65) <= input(18);
output(0, 66) <= input(17);
output(0, 67) <= input(16);
output(0, 68) <= input(0);
output(0, 69) <= input(1);
output(0, 70) <= input(2);
output(0, 71) <= input(3);
output(0, 72) <= input(4);
output(0, 73) <= input(5);
output(0, 74) <= input(6);
output(0, 75) <= input(7);
output(0, 76) <= input(8);
output(0, 77) <= input(9);
output(0, 78) <= input(10);
output(0, 79) <= input(11);
output(0, 80) <= input(20);
output(0, 81) <= input(21);
output(0, 82) <= input(22);
output(0, 83) <= input(23);
output(0, 84) <= input(24);
output(0, 85) <= input(25);
output(0, 86) <= input(26);
output(0, 87) <= input(27);
output(0, 88) <= input(28);
output(0, 89) <= input(29);
output(0, 90) <= input(30);
output(0, 91) <= input(31);
output(0, 92) <= input(32);
output(0, 93) <= input(33);
output(0, 94) <= input(34);
output(0, 95) <= input(35);
output(0, 96) <= input(36);
output(0, 97) <= input(20);
output(0, 98) <= input(21);
output(0, 99) <= input(22);
output(0, 100) <= input(23);
output(0, 101) <= input(24);
output(0, 102) <= input(25);
output(0, 103) <= input(26);
output(0, 104) <= input(27);
output(0, 105) <= input(28);
output(0, 106) <= input(29);
output(0, 107) <= input(30);
output(0, 108) <= input(31);
output(0, 109) <= input(32);
output(0, 110) <= input(33);
output(0, 111) <= input(34);
output(0, 112) <= input(37);
output(0, 113) <= input(36);
output(0, 114) <= input(20);
output(0, 115) <= input(21);
output(0, 116) <= input(22);
output(0, 117) <= input(23);
output(0, 118) <= input(24);
output(0, 119) <= input(25);
output(0, 120) <= input(26);
output(0, 121) <= input(27);
output(0, 122) <= input(28);
output(0, 123) <= input(29);
output(0, 124) <= input(30);
output(0, 125) <= input(31);
output(0, 126) <= input(32);
output(0, 127) <= input(33);
output(0, 128) <= input(38);
output(0, 129) <= input(37);
output(0, 130) <= input(36);
output(0, 131) <= input(20);
output(0, 132) <= input(21);
output(0, 133) <= input(22);
output(0, 134) <= input(23);
output(0, 135) <= input(24);
output(0, 136) <= input(25);
output(0, 137) <= input(26);
output(0, 138) <= input(27);
output(0, 139) <= input(28);
output(0, 140) <= input(29);
output(0, 141) <= input(30);
output(0, 142) <= input(31);
output(0, 143) <= input(32);
output(0, 144) <= input(39);
output(0, 145) <= input(38);
output(0, 146) <= input(37);
output(0, 147) <= input(36);
output(0, 148) <= input(20);
output(0, 149) <= input(21);
output(0, 150) <= input(22);
output(0, 151) <= input(23);
output(0, 152) <= input(24);
output(0, 153) <= input(25);
output(0, 154) <= input(26);
output(0, 155) <= input(27);
output(0, 156) <= input(28);
output(0, 157) <= input(29);
output(0, 158) <= input(30);
output(0, 159) <= input(31);
output(0, 160) <= input(40);
output(0, 161) <= input(41);
output(0, 162) <= input(42);
output(0, 163) <= input(43);
output(0, 164) <= input(44);
output(0, 165) <= input(19);
output(0, 166) <= input(18);
output(0, 167) <= input(17);
output(0, 168) <= input(16);
output(0, 169) <= input(0);
output(0, 170) <= input(1);
output(0, 171) <= input(2);
output(0, 172) <= input(3);
output(0, 173) <= input(4);
output(0, 174) <= input(5);
output(0, 175) <= input(6);
output(0, 176) <= input(45);
output(0, 177) <= input(40);
output(0, 178) <= input(41);
output(0, 179) <= input(42);
output(0, 180) <= input(43);
output(0, 181) <= input(44);
output(0, 182) <= input(19);
output(0, 183) <= input(18);
output(0, 184) <= input(17);
output(0, 185) <= input(16);
output(0, 186) <= input(0);
output(0, 187) <= input(1);
output(0, 188) <= input(2);
output(0, 189) <= input(3);
output(0, 190) <= input(4);
output(0, 191) <= input(5);
output(0, 192) <= input(46);
output(0, 193) <= input(45);
output(0, 194) <= input(40);
output(0, 195) <= input(41);
output(0, 196) <= input(42);
output(0, 197) <= input(43);
output(0, 198) <= input(44);
output(0, 199) <= input(19);
output(0, 200) <= input(18);
output(0, 201) <= input(17);
output(0, 202) <= input(16);
output(0, 203) <= input(0);
output(0, 204) <= input(1);
output(0, 205) <= input(2);
output(0, 206) <= input(3);
output(0, 207) <= input(4);
output(0, 208) <= input(47);
output(0, 209) <= input(46);
output(0, 210) <= input(45);
output(0, 211) <= input(40);
output(0, 212) <= input(41);
output(0, 213) <= input(42);
output(0, 214) <= input(43);
output(0, 215) <= input(44);
output(0, 216) <= input(19);
output(0, 217) <= input(18);
output(0, 218) <= input(17);
output(0, 219) <= input(16);
output(0, 220) <= input(0);
output(0, 221) <= input(1);
output(0, 222) <= input(2);
output(0, 223) <= input(3);
output(0, 224) <= input(48);
output(0, 225) <= input(47);
output(0, 226) <= input(46);
output(0, 227) <= input(45);
output(0, 228) <= input(40);
output(0, 229) <= input(41);
output(0, 230) <= input(42);
output(0, 231) <= input(43);
output(0, 232) <= input(44);
output(0, 233) <= input(19);
output(0, 234) <= input(18);
output(0, 235) <= input(17);
output(0, 236) <= input(16);
output(0, 237) <= input(0);
output(0, 238) <= input(1);
output(0, 239) <= input(2);
output(0, 240) <= input(49);
output(0, 241) <= input(50);
output(0, 242) <= input(51);
output(0, 243) <= input(52);
output(0, 244) <= input(53);
output(0, 245) <= input(39);
output(0, 246) <= input(38);
output(0, 247) <= input(37);
output(0, 248) <= input(36);
output(0, 249) <= input(20);
output(0, 250) <= input(21);
output(0, 251) <= input(22);
output(0, 252) <= input(23);
output(0, 253) <= input(24);
output(0, 254) <= input(25);
output(0, 255) <= input(26);
when "1001" =>
output(0, 0) <= input(0);
output(0, 1) <= input(1);
output(0, 2) <= input(2);
output(0, 3) <= input(3);
output(0, 4) <= input(4);
output(0, 5) <= input(5);
output(0, 6) <= input(6);
output(0, 7) <= input(7);
output(0, 8) <= input(8);
output(0, 9) <= input(9);
output(0, 10) <= input(10);
output(0, 11) <= input(11);
output(0, 12) <= input(12);
output(0, 13) <= input(13);
output(0, 14) <= input(14);
output(0, 15) <= input(15);
output(0, 16) <= input(16);
output(0, 17) <= input(0);
output(0, 18) <= input(1);
output(0, 19) <= input(2);
output(0, 20) <= input(3);
output(0, 21) <= input(4);
output(0, 22) <= input(5);
output(0, 23) <= input(6);
output(0, 24) <= input(7);
output(0, 25) <= input(8);
output(0, 26) <= input(9);
output(0, 27) <= input(10);
output(0, 28) <= input(11);
output(0, 29) <= input(12);
output(0, 30) <= input(13);
output(0, 31) <= input(14);
output(0, 32) <= input(17);
output(0, 33) <= input(18);
output(0, 34) <= input(19);
output(0, 35) <= input(20);
output(0, 36) <= input(21);
output(0, 37) <= input(22);
output(0, 38) <= input(23);
output(0, 39) <= input(24);
output(0, 40) <= input(25);
output(0, 41) <= input(26);
output(0, 42) <= input(27);
output(0, 43) <= input(28);
output(0, 44) <= input(29);
output(0, 45) <= input(30);
output(0, 46) <= input(31);
output(0, 47) <= input(32);
output(0, 48) <= input(33);
output(0, 49) <= input(17);
output(0, 50) <= input(18);
output(0, 51) <= input(19);
output(0, 52) <= input(20);
output(0, 53) <= input(21);
output(0, 54) <= input(22);
output(0, 55) <= input(23);
output(0, 56) <= input(24);
output(0, 57) <= input(25);
output(0, 58) <= input(26);
output(0, 59) <= input(27);
output(0, 60) <= input(28);
output(0, 61) <= input(29);
output(0, 62) <= input(30);
output(0, 63) <= input(31);
output(0, 64) <= input(34);
output(0, 65) <= input(33);
output(0, 66) <= input(17);
output(0, 67) <= input(18);
output(0, 68) <= input(19);
output(0, 69) <= input(20);
output(0, 70) <= input(21);
output(0, 71) <= input(22);
output(0, 72) <= input(23);
output(0, 73) <= input(24);
output(0, 74) <= input(25);
output(0, 75) <= input(26);
output(0, 76) <= input(27);
output(0, 77) <= input(28);
output(0, 78) <= input(29);
output(0, 79) <= input(30);
output(0, 80) <= input(35);
output(0, 81) <= input(36);
output(0, 82) <= input(37);
output(0, 83) <= input(16);
output(0, 84) <= input(0);
output(0, 85) <= input(1);
output(0, 86) <= input(2);
output(0, 87) <= input(3);
output(0, 88) <= input(4);
output(0, 89) <= input(5);
output(0, 90) <= input(6);
output(0, 91) <= input(7);
output(0, 92) <= input(8);
output(0, 93) <= input(9);
output(0, 94) <= input(10);
output(0, 95) <= input(11);
output(0, 96) <= input(38);
output(0, 97) <= input(35);
output(0, 98) <= input(36);
output(0, 99) <= input(37);
output(0, 100) <= input(16);
output(0, 101) <= input(0);
output(0, 102) <= input(1);
output(0, 103) <= input(2);
output(0, 104) <= input(3);
output(0, 105) <= input(4);
output(0, 106) <= input(5);
output(0, 107) <= input(6);
output(0, 108) <= input(7);
output(0, 109) <= input(8);
output(0, 110) <= input(9);
output(0, 111) <= input(10);
output(0, 112) <= input(39);
output(0, 113) <= input(40);
output(0, 114) <= input(34);
output(0, 115) <= input(33);
output(0, 116) <= input(17);
output(0, 117) <= input(18);
output(0, 118) <= input(19);
output(0, 119) <= input(20);
output(0, 120) <= input(21);
output(0, 121) <= input(22);
output(0, 122) <= input(23);
output(0, 123) <= input(24);
output(0, 124) <= input(25);
output(0, 125) <= input(26);
output(0, 126) <= input(27);
output(0, 127) <= input(28);
output(0, 128) <= input(41);
output(0, 129) <= input(39);
output(0, 130) <= input(40);
output(0, 131) <= input(34);
output(0, 132) <= input(33);
output(0, 133) <= input(17);
output(0, 134) <= input(18);
output(0, 135) <= input(19);
output(0, 136) <= input(20);
output(0, 137) <= input(21);
output(0, 138) <= input(22);
output(0, 139) <= input(23);
output(0, 140) <= input(24);
output(0, 141) <= input(25);
output(0, 142) <= input(26);
output(0, 143) <= input(27);
output(0, 144) <= input(42);
output(0, 145) <= input(41);
output(0, 146) <= input(39);
output(0, 147) <= input(40);
output(0, 148) <= input(34);
output(0, 149) <= input(33);
output(0, 150) <= input(17);
output(0, 151) <= input(18);
output(0, 152) <= input(19);
output(0, 153) <= input(20);
output(0, 154) <= input(21);
output(0, 155) <= input(22);
output(0, 156) <= input(23);
output(0, 157) <= input(24);
output(0, 158) <= input(25);
output(0, 159) <= input(26);
output(0, 160) <= input(43);
output(0, 161) <= input(44);
output(0, 162) <= input(45);
output(0, 163) <= input(38);
output(0, 164) <= input(35);
output(0, 165) <= input(36);
output(0, 166) <= input(37);
output(0, 167) <= input(16);
output(0, 168) <= input(0);
output(0, 169) <= input(1);
output(0, 170) <= input(2);
output(0, 171) <= input(3);
output(0, 172) <= input(4);
output(0, 173) <= input(5);
output(0, 174) <= input(6);
output(0, 175) <= input(7);
output(0, 176) <= input(46);
output(0, 177) <= input(43);
output(0, 178) <= input(44);
output(0, 179) <= input(45);
output(0, 180) <= input(38);
output(0, 181) <= input(35);
output(0, 182) <= input(36);
output(0, 183) <= input(37);
output(0, 184) <= input(16);
output(0, 185) <= input(0);
output(0, 186) <= input(1);
output(0, 187) <= input(2);
output(0, 188) <= input(3);
output(0, 189) <= input(4);
output(0, 190) <= input(5);
output(0, 191) <= input(6);
output(0, 192) <= input(47);
output(0, 193) <= input(46);
output(0, 194) <= input(43);
output(0, 195) <= input(44);
output(0, 196) <= input(45);
output(0, 197) <= input(38);
output(0, 198) <= input(35);
output(0, 199) <= input(36);
output(0, 200) <= input(37);
output(0, 201) <= input(16);
output(0, 202) <= input(0);
output(0, 203) <= input(1);
output(0, 204) <= input(2);
output(0, 205) <= input(3);
output(0, 206) <= input(4);
output(0, 207) <= input(5);
output(0, 208) <= input(48);
output(0, 209) <= input(49);
output(0, 210) <= input(50);
output(0, 211) <= input(42);
output(0, 212) <= input(41);
output(0, 213) <= input(39);
output(0, 214) <= input(40);
output(0, 215) <= input(34);
output(0, 216) <= input(33);
output(0, 217) <= input(17);
output(0, 218) <= input(18);
output(0, 219) <= input(19);
output(0, 220) <= input(20);
output(0, 221) <= input(21);
output(0, 222) <= input(22);
output(0, 223) <= input(23);
output(0, 224) <= input(51);
output(0, 225) <= input(48);
output(0, 226) <= input(49);
output(0, 227) <= input(50);
output(0, 228) <= input(42);
output(0, 229) <= input(41);
output(0, 230) <= input(39);
output(0, 231) <= input(40);
output(0, 232) <= input(34);
output(0, 233) <= input(33);
output(0, 234) <= input(17);
output(0, 235) <= input(18);
output(0, 236) <= input(19);
output(0, 237) <= input(20);
output(0, 238) <= input(21);
output(0, 239) <= input(22);
output(0, 240) <= input(52);
output(0, 241) <= input(53);
output(0, 242) <= input(47);
output(0, 243) <= input(46);
output(0, 244) <= input(43);
output(0, 245) <= input(44);
output(0, 246) <= input(45);
output(0, 247) <= input(38);
output(0, 248) <= input(35);
output(0, 249) <= input(36);
output(0, 250) <= input(37);
output(0, 251) <= input(16);
output(0, 252) <= input(0);
output(0, 253) <= input(1);
output(0, 254) <= input(2);
output(0, 255) <= input(3);
output(1, 0) <= input(20);
output(1, 1) <= input(21);
output(1, 2) <= input(22);
output(1, 3) <= input(23);
output(1, 4) <= input(24);
output(1, 5) <= input(25);
output(1, 6) <= input(26);
output(1, 7) <= input(27);
output(1, 8) <= input(28);
output(1, 9) <= input(29);
output(1, 10) <= input(30);
output(1, 11) <= input(31);
output(1, 12) <= input(32);
output(1, 13) <= input(54);
output(1, 14) <= input(55);
output(1, 15) <= input(56);
output(1, 16) <= input(1);
output(1, 17) <= input(2);
output(1, 18) <= input(3);
output(1, 19) <= input(4);
output(1, 20) <= input(5);
output(1, 21) <= input(6);
output(1, 22) <= input(7);
output(1, 23) <= input(8);
output(1, 24) <= input(9);
output(1, 25) <= input(10);
output(1, 26) <= input(11);
output(1, 27) <= input(12);
output(1, 28) <= input(13);
output(1, 29) <= input(14);
output(1, 30) <= input(15);
output(1, 31) <= input(57);
output(1, 32) <= input(0);
output(1, 33) <= input(1);
output(1, 34) <= input(2);
output(1, 35) <= input(3);
output(1, 36) <= input(4);
output(1, 37) <= input(5);
output(1, 38) <= input(6);
output(1, 39) <= input(7);
output(1, 40) <= input(8);
output(1, 41) <= input(9);
output(1, 42) <= input(10);
output(1, 43) <= input(11);
output(1, 44) <= input(12);
output(1, 45) <= input(13);
output(1, 46) <= input(14);
output(1, 47) <= input(15);
output(1, 48) <= input(18);
output(1, 49) <= input(19);
output(1, 50) <= input(20);
output(1, 51) <= input(21);
output(1, 52) <= input(22);
output(1, 53) <= input(23);
output(1, 54) <= input(24);
output(1, 55) <= input(25);
output(1, 56) <= input(26);
output(1, 57) <= input(27);
output(1, 58) <= input(28);
output(1, 59) <= input(29);
output(1, 60) <= input(30);
output(1, 61) <= input(31);
output(1, 62) <= input(32);
output(1, 63) <= input(54);
output(1, 64) <= input(17);
output(1, 65) <= input(18);
output(1, 66) <= input(19);
output(1, 67) <= input(20);
output(1, 68) <= input(21);
output(1, 69) <= input(22);
output(1, 70) <= input(23);
output(1, 71) <= input(24);
output(1, 72) <= input(25);
output(1, 73) <= input(26);
output(1, 74) <= input(27);
output(1, 75) <= input(28);
output(1, 76) <= input(29);
output(1, 77) <= input(30);
output(1, 78) <= input(31);
output(1, 79) <= input(32);
output(1, 80) <= input(37);
output(1, 81) <= input(16);
output(1, 82) <= input(0);
output(1, 83) <= input(1);
output(1, 84) <= input(2);
output(1, 85) <= input(3);
output(1, 86) <= input(4);
output(1, 87) <= input(5);
output(1, 88) <= input(6);
output(1, 89) <= input(7);
output(1, 90) <= input(8);
output(1, 91) <= input(9);
output(1, 92) <= input(10);
output(1, 93) <= input(11);
output(1, 94) <= input(12);
output(1, 95) <= input(13);
output(1, 96) <= input(36);
output(1, 97) <= input(37);
output(1, 98) <= input(16);
output(1, 99) <= input(0);
output(1, 100) <= input(1);
output(1, 101) <= input(2);
output(1, 102) <= input(3);
output(1, 103) <= input(4);
output(1, 104) <= input(5);
output(1, 105) <= input(6);
output(1, 106) <= input(7);
output(1, 107) <= input(8);
output(1, 108) <= input(9);
output(1, 109) <= input(10);
output(1, 110) <= input(11);
output(1, 111) <= input(12);
output(1, 112) <= input(34);
output(1, 113) <= input(33);
output(1, 114) <= input(17);
output(1, 115) <= input(18);
output(1, 116) <= input(19);
output(1, 117) <= input(20);
output(1, 118) <= input(21);
output(1, 119) <= input(22);
output(1, 120) <= input(23);
output(1, 121) <= input(24);
output(1, 122) <= input(25);
output(1, 123) <= input(26);
output(1, 124) <= input(27);
output(1, 125) <= input(28);
output(1, 126) <= input(29);
output(1, 127) <= input(30);
output(1, 128) <= input(35);
output(1, 129) <= input(36);
output(1, 130) <= input(37);
output(1, 131) <= input(16);
output(1, 132) <= input(0);
output(1, 133) <= input(1);
output(1, 134) <= input(2);
output(1, 135) <= input(3);
output(1, 136) <= input(4);
output(1, 137) <= input(5);
output(1, 138) <= input(6);
output(1, 139) <= input(7);
output(1, 140) <= input(8);
output(1, 141) <= input(9);
output(1, 142) <= input(10);
output(1, 143) <= input(11);
output(1, 144) <= input(38);
output(1, 145) <= input(35);
output(1, 146) <= input(36);
output(1, 147) <= input(37);
output(1, 148) <= input(16);
output(1, 149) <= input(0);
output(1, 150) <= input(1);
output(1, 151) <= input(2);
output(1, 152) <= input(3);
output(1, 153) <= input(4);
output(1, 154) <= input(5);
output(1, 155) <= input(6);
output(1, 156) <= input(7);
output(1, 157) <= input(8);
output(1, 158) <= input(9);
output(1, 159) <= input(10);
output(1, 160) <= input(39);
output(1, 161) <= input(40);
output(1, 162) <= input(34);
output(1, 163) <= input(33);
output(1, 164) <= input(17);
output(1, 165) <= input(18);
output(1, 166) <= input(19);
output(1, 167) <= input(20);
output(1, 168) <= input(21);
output(1, 169) <= input(22);
output(1, 170) <= input(23);
output(1, 171) <= input(24);
output(1, 172) <= input(25);
output(1, 173) <= input(26);
output(1, 174) <= input(27);
output(1, 175) <= input(28);
output(1, 176) <= input(41);
output(1, 177) <= input(39);
output(1, 178) <= input(40);
output(1, 179) <= input(34);
output(1, 180) <= input(33);
output(1, 181) <= input(17);
output(1, 182) <= input(18);
output(1, 183) <= input(19);
output(1, 184) <= input(20);
output(1, 185) <= input(21);
output(1, 186) <= input(22);
output(1, 187) <= input(23);
output(1, 188) <= input(24);
output(1, 189) <= input(25);
output(1, 190) <= input(26);
output(1, 191) <= input(27);
output(1, 192) <= input(44);
output(1, 193) <= input(45);
output(1, 194) <= input(38);
output(1, 195) <= input(35);
output(1, 196) <= input(36);
output(1, 197) <= input(37);
output(1, 198) <= input(16);
output(1, 199) <= input(0);
output(1, 200) <= input(1);
output(1, 201) <= input(2);
output(1, 202) <= input(3);
output(1, 203) <= input(4);
output(1, 204) <= input(5);
output(1, 205) <= input(6);
output(1, 206) <= input(7);
output(1, 207) <= input(8);
output(1, 208) <= input(43);
output(1, 209) <= input(44);
output(1, 210) <= input(45);
output(1, 211) <= input(38);
output(1, 212) <= input(35);
output(1, 213) <= input(36);
output(1, 214) <= input(37);
output(1, 215) <= input(16);
output(1, 216) <= input(0);
output(1, 217) <= input(1);
output(1, 218) <= input(2);
output(1, 219) <= input(3);
output(1, 220) <= input(4);
output(1, 221) <= input(5);
output(1, 222) <= input(6);
output(1, 223) <= input(7);
output(1, 224) <= input(50);
output(1, 225) <= input(42);
output(1, 226) <= input(41);
output(1, 227) <= input(39);
output(1, 228) <= input(40);
output(1, 229) <= input(34);
output(1, 230) <= input(33);
output(1, 231) <= input(17);
output(1, 232) <= input(18);
output(1, 233) <= input(19);
output(1, 234) <= input(20);
output(1, 235) <= input(21);
output(1, 236) <= input(22);
output(1, 237) <= input(23);
output(1, 238) <= input(24);
output(1, 239) <= input(25);
output(1, 240) <= input(46);
output(1, 241) <= input(43);
output(1, 242) <= input(44);
output(1, 243) <= input(45);
output(1, 244) <= input(38);
output(1, 245) <= input(35);
output(1, 246) <= input(36);
output(1, 247) <= input(37);
output(1, 248) <= input(16);
output(1, 249) <= input(0);
output(1, 250) <= input(1);
output(1, 251) <= input(2);
output(1, 252) <= input(3);
output(1, 253) <= input(4);
output(1, 254) <= input(5);
output(1, 255) <= input(6);
output(2, 0) <= input(3);
output(2, 1) <= input(4);
output(2, 2) <= input(5);
output(2, 3) <= input(6);
output(2, 4) <= input(7);
output(2, 5) <= input(8);
output(2, 6) <= input(9);
output(2, 7) <= input(10);
output(2, 8) <= input(11);
output(2, 9) <= input(12);
output(2, 10) <= input(13);
output(2, 11) <= input(14);
output(2, 12) <= input(15);
output(2, 13) <= input(57);
output(2, 14) <= input(58);
output(2, 15) <= input(59);
output(2, 16) <= input(21);
output(2, 17) <= input(22);
output(2, 18) <= input(23);
output(2, 19) <= input(24);
output(2, 20) <= input(25);
output(2, 21) <= input(26);
output(2, 22) <= input(27);
output(2, 23) <= input(28);
output(2, 24) <= input(29);
output(2, 25) <= input(30);
output(2, 26) <= input(31);
output(2, 27) <= input(32);
output(2, 28) <= input(54);
output(2, 29) <= input(55);
output(2, 30) <= input(56);
output(2, 31) <= input(60);
output(2, 32) <= input(2);
output(2, 33) <= input(3);
output(2, 34) <= input(4);
output(2, 35) <= input(5);
output(2, 36) <= input(6);
output(2, 37) <= input(7);
output(2, 38) <= input(8);
output(2, 39) <= input(9);
output(2, 40) <= input(10);
output(2, 41) <= input(11);
output(2, 42) <= input(12);
output(2, 43) <= input(13);
output(2, 44) <= input(14);
output(2, 45) <= input(15);
output(2, 46) <= input(57);
output(2, 47) <= input(58);
output(2, 48) <= input(20);
output(2, 49) <= input(21);
output(2, 50) <= input(22);
output(2, 51) <= input(23);
output(2, 52) <= input(24);
output(2, 53) <= input(25);
output(2, 54) <= input(26);
output(2, 55) <= input(27);
output(2, 56) <= input(28);
output(2, 57) <= input(29);
output(2, 58) <= input(30);
output(2, 59) <= input(31);
output(2, 60) <= input(32);
output(2, 61) <= input(54);
output(2, 62) <= input(55);
output(2, 63) <= input(56);
output(2, 64) <= input(19);
output(2, 65) <= input(20);
output(2, 66) <= input(21);
output(2, 67) <= input(22);
output(2, 68) <= input(23);
output(2, 69) <= input(24);
output(2, 70) <= input(25);
output(2, 71) <= input(26);
output(2, 72) <= input(27);
output(2, 73) <= input(28);
output(2, 74) <= input(29);
output(2, 75) <= input(30);
output(2, 76) <= input(31);
output(2, 77) <= input(32);
output(2, 78) <= input(54);
output(2, 79) <= input(55);
output(2, 80) <= input(0);
output(2, 81) <= input(1);
output(2, 82) <= input(2);
output(2, 83) <= input(3);
output(2, 84) <= input(4);
output(2, 85) <= input(5);
output(2, 86) <= input(6);
output(2, 87) <= input(7);
output(2, 88) <= input(8);
output(2, 89) <= input(9);
output(2, 90) <= input(10);
output(2, 91) <= input(11);
output(2, 92) <= input(12);
output(2, 93) <= input(13);
output(2, 94) <= input(14);
output(2, 95) <= input(15);
output(2, 96) <= input(18);
output(2, 97) <= input(19);
output(2, 98) <= input(20);
output(2, 99) <= input(21);
output(2, 100) <= input(22);
output(2, 101) <= input(23);
output(2, 102) <= input(24);
output(2, 103) <= input(25);
output(2, 104) <= input(26);
output(2, 105) <= input(27);
output(2, 106) <= input(28);
output(2, 107) <= input(29);
output(2, 108) <= input(30);
output(2, 109) <= input(31);
output(2, 110) <= input(32);
output(2, 111) <= input(54);
output(2, 112) <= input(16);
output(2, 113) <= input(0);
output(2, 114) <= input(1);
output(2, 115) <= input(2);
output(2, 116) <= input(3);
output(2, 117) <= input(4);
output(2, 118) <= input(5);
output(2, 119) <= input(6);
output(2, 120) <= input(7);
output(2, 121) <= input(8);
output(2, 122) <= input(9);
output(2, 123) <= input(10);
output(2, 124) <= input(11);
output(2, 125) <= input(12);
output(2, 126) <= input(13);
output(2, 127) <= input(14);
output(2, 128) <= input(37);
output(2, 129) <= input(16);
output(2, 130) <= input(0);
output(2, 131) <= input(1);
output(2, 132) <= input(2);
output(2, 133) <= input(3);
output(2, 134) <= input(4);
output(2, 135) <= input(5);
output(2, 136) <= input(6);
output(2, 137) <= input(7);
output(2, 138) <= input(8);
output(2, 139) <= input(9);
output(2, 140) <= input(10);
output(2, 141) <= input(11);
output(2, 142) <= input(12);
output(2, 143) <= input(13);
output(2, 144) <= input(33);
output(2, 145) <= input(17);
output(2, 146) <= input(18);
output(2, 147) <= input(19);
output(2, 148) <= input(20);
output(2, 149) <= input(21);
output(2, 150) <= input(22);
output(2, 151) <= input(23);
output(2, 152) <= input(24);
output(2, 153) <= input(25);
output(2, 154) <= input(26);
output(2, 155) <= input(27);
output(2, 156) <= input(28);
output(2, 157) <= input(29);
output(2, 158) <= input(30);
output(2, 159) <= input(31);
output(2, 160) <= input(36);
output(2, 161) <= input(37);
output(2, 162) <= input(16);
output(2, 163) <= input(0);
output(2, 164) <= input(1);
output(2, 165) <= input(2);
output(2, 166) <= input(3);
output(2, 167) <= input(4);
output(2, 168) <= input(5);
output(2, 169) <= input(6);
output(2, 170) <= input(7);
output(2, 171) <= input(8);
output(2, 172) <= input(9);
output(2, 173) <= input(10);
output(2, 174) <= input(11);
output(2, 175) <= input(12);
output(2, 176) <= input(34);
output(2, 177) <= input(33);
output(2, 178) <= input(17);
output(2, 179) <= input(18);
output(2, 180) <= input(19);
output(2, 181) <= input(20);
output(2, 182) <= input(21);
output(2, 183) <= input(22);
output(2, 184) <= input(23);
output(2, 185) <= input(24);
output(2, 186) <= input(25);
output(2, 187) <= input(26);
output(2, 188) <= input(27);
output(2, 189) <= input(28);
output(2, 190) <= input(29);
output(2, 191) <= input(30);
output(2, 192) <= input(40);
output(2, 193) <= input(34);
output(2, 194) <= input(33);
output(2, 195) <= input(17);
output(2, 196) <= input(18);
output(2, 197) <= input(19);
output(2, 198) <= input(20);
output(2, 199) <= input(21);
output(2, 200) <= input(22);
output(2, 201) <= input(23);
output(2, 202) <= input(24);
output(2, 203) <= input(25);
output(2, 204) <= input(26);
output(2, 205) <= input(27);
output(2, 206) <= input(28);
output(2, 207) <= input(29);
output(2, 208) <= input(38);
output(2, 209) <= input(35);
output(2, 210) <= input(36);
output(2, 211) <= input(37);
output(2, 212) <= input(16);
output(2, 213) <= input(0);
output(2, 214) <= input(1);
output(2, 215) <= input(2);
output(2, 216) <= input(3);
output(2, 217) <= input(4);
output(2, 218) <= input(5);
output(2, 219) <= input(6);
output(2, 220) <= input(7);
output(2, 221) <= input(8);
output(2, 222) <= input(9);
output(2, 223) <= input(10);
output(2, 224) <= input(39);
output(2, 225) <= input(40);
output(2, 226) <= input(34);
output(2, 227) <= input(33);
output(2, 228) <= input(17);
output(2, 229) <= input(18);
output(2, 230) <= input(19);
output(2, 231) <= input(20);
output(2, 232) <= input(21);
output(2, 233) <= input(22);
output(2, 234) <= input(23);
output(2, 235) <= input(24);
output(2, 236) <= input(25);
output(2, 237) <= input(26);
output(2, 238) <= input(27);
output(2, 239) <= input(28);
output(2, 240) <= input(45);
output(2, 241) <= input(38);
output(2, 242) <= input(35);
output(2, 243) <= input(36);
output(2, 244) <= input(37);
output(2, 245) <= input(16);
output(2, 246) <= input(0);
output(2, 247) <= input(1);
output(2, 248) <= input(2);
output(2, 249) <= input(3);
output(2, 250) <= input(4);
output(2, 251) <= input(5);
output(2, 252) <= input(6);
output(2, 253) <= input(7);
output(2, 254) <= input(8);
output(2, 255) <= input(9);
when "1010" =>
output(0, 0) <= input(0);
output(0, 1) <= input(1);
output(0, 2) <= input(2);
output(0, 3) <= input(3);
output(0, 4) <= input(4);
output(0, 5) <= input(5);
output(0, 6) <= input(6);
output(0, 7) <= input(7);
output(0, 8) <= input(8);
output(0, 9) <= input(9);
output(0, 10) <= input(10);
output(0, 11) <= input(11);
output(0, 12) <= input(12);
output(0, 13) <= input(13);
output(0, 14) <= input(14);
output(0, 15) <= input(15);
output(0, 16) <= input(16);
output(0, 17) <= input(17);
output(0, 18) <= input(18);
output(0, 19) <= input(19);
output(0, 20) <= input(20);
output(0, 21) <= input(21);
output(0, 22) <= input(22);
output(0, 23) <= input(23);
output(0, 24) <= input(24);
output(0, 25) <= input(25);
output(0, 26) <= input(26);
output(0, 27) <= input(27);
output(0, 28) <= input(28);
output(0, 29) <= input(29);
output(0, 30) <= input(30);
output(0, 31) <= input(31);
output(0, 32) <= input(32);
output(0, 33) <= input(0);
output(0, 34) <= input(1);
output(0, 35) <= input(2);
output(0, 36) <= input(3);
output(0, 37) <= input(4);
output(0, 38) <= input(5);
output(0, 39) <= input(6);
output(0, 40) <= input(7);
output(0, 41) <= input(8);
output(0, 42) <= input(9);
output(0, 43) <= input(10);
output(0, 44) <= input(11);
output(0, 45) <= input(12);
output(0, 46) <= input(13);
output(0, 47) <= input(14);
output(0, 48) <= input(33);
output(0, 49) <= input(16);
output(0, 50) <= input(17);
output(0, 51) <= input(18);
output(0, 52) <= input(19);
output(0, 53) <= input(20);
output(0, 54) <= input(21);
output(0, 55) <= input(22);
output(0, 56) <= input(23);
output(0, 57) <= input(24);
output(0, 58) <= input(25);
output(0, 59) <= input(26);
output(0, 60) <= input(27);
output(0, 61) <= input(28);
output(0, 62) <= input(29);
output(0, 63) <= input(30);
output(0, 64) <= input(34);
output(0, 65) <= input(32);
output(0, 66) <= input(0);
output(0, 67) <= input(1);
output(0, 68) <= input(2);
output(0, 69) <= input(3);
output(0, 70) <= input(4);
output(0, 71) <= input(5);
output(0, 72) <= input(6);
output(0, 73) <= input(7);
output(0, 74) <= input(8);
output(0, 75) <= input(9);
output(0, 76) <= input(10);
output(0, 77) <= input(11);
output(0, 78) <= input(12);
output(0, 79) <= input(13);
output(0, 80) <= input(35);
output(0, 81) <= input(33);
output(0, 82) <= input(16);
output(0, 83) <= input(17);
output(0, 84) <= input(18);
output(0, 85) <= input(19);
output(0, 86) <= input(20);
output(0, 87) <= input(21);
output(0, 88) <= input(22);
output(0, 89) <= input(23);
output(0, 90) <= input(24);
output(0, 91) <= input(25);
output(0, 92) <= input(26);
output(0, 93) <= input(27);
output(0, 94) <= input(28);
output(0, 95) <= input(29);
output(0, 96) <= input(36);
output(0, 97) <= input(34);
output(0, 98) <= input(32);
output(0, 99) <= input(0);
output(0, 100) <= input(1);
output(0, 101) <= input(2);
output(0, 102) <= input(3);
output(0, 103) <= input(4);
output(0, 104) <= input(5);
output(0, 105) <= input(6);
output(0, 106) <= input(7);
output(0, 107) <= input(8);
output(0, 108) <= input(9);
output(0, 109) <= input(10);
output(0, 110) <= input(11);
output(0, 111) <= input(12);
output(0, 112) <= input(37);
output(0, 113) <= input(35);
output(0, 114) <= input(33);
output(0, 115) <= input(16);
output(0, 116) <= input(17);
output(0, 117) <= input(18);
output(0, 118) <= input(19);
output(0, 119) <= input(20);
output(0, 120) <= input(21);
output(0, 121) <= input(22);
output(0, 122) <= input(23);
output(0, 123) <= input(24);
output(0, 124) <= input(25);
output(0, 125) <= input(26);
output(0, 126) <= input(27);
output(0, 127) <= input(28);
output(0, 128) <= input(38);
output(0, 129) <= input(37);
output(0, 130) <= input(35);
output(0, 131) <= input(33);
output(0, 132) <= input(16);
output(0, 133) <= input(17);
output(0, 134) <= input(18);
output(0, 135) <= input(19);
output(0, 136) <= input(20);
output(0, 137) <= input(21);
output(0, 138) <= input(22);
output(0, 139) <= input(23);
output(0, 140) <= input(24);
output(0, 141) <= input(25);
output(0, 142) <= input(26);
output(0, 143) <= input(27);
output(0, 144) <= input(39);
output(0, 145) <= input(40);
output(0, 146) <= input(36);
output(0, 147) <= input(34);
output(0, 148) <= input(32);
output(0, 149) <= input(0);
output(0, 150) <= input(1);
output(0, 151) <= input(2);
output(0, 152) <= input(3);
output(0, 153) <= input(4);
output(0, 154) <= input(5);
output(0, 155) <= input(6);
output(0, 156) <= input(7);
output(0, 157) <= input(8);
output(0, 158) <= input(9);
output(0, 159) <= input(10);
output(0, 160) <= input(41);
output(0, 161) <= input(38);
output(0, 162) <= input(37);
output(0, 163) <= input(35);
output(0, 164) <= input(33);
output(0, 165) <= input(16);
output(0, 166) <= input(17);
output(0, 167) <= input(18);
output(0, 168) <= input(19);
output(0, 169) <= input(20);
output(0, 170) <= input(21);
output(0, 171) <= input(22);
output(0, 172) <= input(23);
output(0, 173) <= input(24);
output(0, 174) <= input(25);
output(0, 175) <= input(26);
output(0, 176) <= input(42);
output(0, 177) <= input(39);
output(0, 178) <= input(40);
output(0, 179) <= input(36);
output(0, 180) <= input(34);
output(0, 181) <= input(32);
output(0, 182) <= input(0);
output(0, 183) <= input(1);
output(0, 184) <= input(2);
output(0, 185) <= input(3);
output(0, 186) <= input(4);
output(0, 187) <= input(5);
output(0, 188) <= input(6);
output(0, 189) <= input(7);
output(0, 190) <= input(8);
output(0, 191) <= input(9);
output(0, 192) <= input(43);
output(0, 193) <= input(41);
output(0, 194) <= input(38);
output(0, 195) <= input(37);
output(0, 196) <= input(35);
output(0, 197) <= input(33);
output(0, 198) <= input(16);
output(0, 199) <= input(17);
output(0, 200) <= input(18);
output(0, 201) <= input(19);
output(0, 202) <= input(20);
output(0, 203) <= input(21);
output(0, 204) <= input(22);
output(0, 205) <= input(23);
output(0, 206) <= input(24);
output(0, 207) <= input(25);
output(0, 208) <= input(44);
output(0, 209) <= input(42);
output(0, 210) <= input(39);
output(0, 211) <= input(40);
output(0, 212) <= input(36);
output(0, 213) <= input(34);
output(0, 214) <= input(32);
output(0, 215) <= input(0);
output(0, 216) <= input(1);
output(0, 217) <= input(2);
output(0, 218) <= input(3);
output(0, 219) <= input(4);
output(0, 220) <= input(5);
output(0, 221) <= input(6);
output(0, 222) <= input(7);
output(0, 223) <= input(8);
output(0, 224) <= input(45);
output(0, 225) <= input(43);
output(0, 226) <= input(41);
output(0, 227) <= input(38);
output(0, 228) <= input(37);
output(0, 229) <= input(35);
output(0, 230) <= input(33);
output(0, 231) <= input(16);
output(0, 232) <= input(17);
output(0, 233) <= input(18);
output(0, 234) <= input(19);
output(0, 235) <= input(20);
output(0, 236) <= input(21);
output(0, 237) <= input(22);
output(0, 238) <= input(23);
output(0, 239) <= input(24);
output(0, 240) <= input(46);
output(0, 241) <= input(44);
output(0, 242) <= input(42);
output(0, 243) <= input(39);
output(0, 244) <= input(40);
output(0, 245) <= input(36);
output(0, 246) <= input(34);
output(0, 247) <= input(32);
output(0, 248) <= input(0);
output(0, 249) <= input(1);
output(0, 250) <= input(2);
output(0, 251) <= input(3);
output(0, 252) <= input(4);
output(0, 253) <= input(5);
output(0, 254) <= input(6);
output(0, 255) <= input(7);
output(1, 0) <= input(18);
output(1, 1) <= input(19);
output(1, 2) <= input(20);
output(1, 3) <= input(21);
output(1, 4) <= input(22);
output(1, 5) <= input(23);
output(1, 6) <= input(24);
output(1, 7) <= input(25);
output(1, 8) <= input(26);
output(1, 9) <= input(27);
output(1, 10) <= input(28);
output(1, 11) <= input(29);
output(1, 12) <= input(30);
output(1, 13) <= input(31);
output(1, 14) <= input(47);
output(1, 15) <= input(48);
output(1, 16) <= input(1);
output(1, 17) <= input(2);
output(1, 18) <= input(3);
output(1, 19) <= input(4);
output(1, 20) <= input(5);
output(1, 21) <= input(6);
output(1, 22) <= input(7);
output(1, 23) <= input(8);
output(1, 24) <= input(9);
output(1, 25) <= input(10);
output(1, 26) <= input(11);
output(1, 27) <= input(12);
output(1, 28) <= input(13);
output(1, 29) <= input(14);
output(1, 30) <= input(15);
output(1, 31) <= input(49);
output(1, 32) <= input(17);
output(1, 33) <= input(18);
output(1, 34) <= input(19);
output(1, 35) <= input(20);
output(1, 36) <= input(21);
output(1, 37) <= input(22);
output(1, 38) <= input(23);
output(1, 39) <= input(24);
output(1, 40) <= input(25);
output(1, 41) <= input(26);
output(1, 42) <= input(27);
output(1, 43) <= input(28);
output(1, 44) <= input(29);
output(1, 45) <= input(30);
output(1, 46) <= input(31);
output(1, 47) <= input(47);
output(1, 48) <= input(0);
output(1, 49) <= input(1);
output(1, 50) <= input(2);
output(1, 51) <= input(3);
output(1, 52) <= input(4);
output(1, 53) <= input(5);
output(1, 54) <= input(6);
output(1, 55) <= input(7);
output(1, 56) <= input(8);
output(1, 57) <= input(9);
output(1, 58) <= input(10);
output(1, 59) <= input(11);
output(1, 60) <= input(12);
output(1, 61) <= input(13);
output(1, 62) <= input(14);
output(1, 63) <= input(15);
output(1, 64) <= input(16);
output(1, 65) <= input(17);
output(1, 66) <= input(18);
output(1, 67) <= input(19);
output(1, 68) <= input(20);
output(1, 69) <= input(21);
output(1, 70) <= input(22);
output(1, 71) <= input(23);
output(1, 72) <= input(24);
output(1, 73) <= input(25);
output(1, 74) <= input(26);
output(1, 75) <= input(27);
output(1, 76) <= input(28);
output(1, 77) <= input(29);
output(1, 78) <= input(30);
output(1, 79) <= input(31);
output(1, 80) <= input(32);
output(1, 81) <= input(0);
output(1, 82) <= input(1);
output(1, 83) <= input(2);
output(1, 84) <= input(3);
output(1, 85) <= input(4);
output(1, 86) <= input(5);
output(1, 87) <= input(6);
output(1, 88) <= input(7);
output(1, 89) <= input(8);
output(1, 90) <= input(9);
output(1, 91) <= input(10);
output(1, 92) <= input(11);
output(1, 93) <= input(12);
output(1, 94) <= input(13);
output(1, 95) <= input(14);
output(1, 96) <= input(33);
output(1, 97) <= input(16);
output(1, 98) <= input(17);
output(1, 99) <= input(18);
output(1, 100) <= input(19);
output(1, 101) <= input(20);
output(1, 102) <= input(21);
output(1, 103) <= input(22);
output(1, 104) <= input(23);
output(1, 105) <= input(24);
output(1, 106) <= input(25);
output(1, 107) <= input(26);
output(1, 108) <= input(27);
output(1, 109) <= input(28);
output(1, 110) <= input(29);
output(1, 111) <= input(30);
output(1, 112) <= input(34);
output(1, 113) <= input(32);
output(1, 114) <= input(0);
output(1, 115) <= input(1);
output(1, 116) <= input(2);
output(1, 117) <= input(3);
output(1, 118) <= input(4);
output(1, 119) <= input(5);
output(1, 120) <= input(6);
output(1, 121) <= input(7);
output(1, 122) <= input(8);
output(1, 123) <= input(9);
output(1, 124) <= input(10);
output(1, 125) <= input(11);
output(1, 126) <= input(12);
output(1, 127) <= input(13);
output(1, 128) <= input(35);
output(1, 129) <= input(33);
output(1, 130) <= input(16);
output(1, 131) <= input(17);
output(1, 132) <= input(18);
output(1, 133) <= input(19);
output(1, 134) <= input(20);
output(1, 135) <= input(21);
output(1, 136) <= input(22);
output(1, 137) <= input(23);
output(1, 138) <= input(24);
output(1, 139) <= input(25);
output(1, 140) <= input(26);
output(1, 141) <= input(27);
output(1, 142) <= input(28);
output(1, 143) <= input(29);
output(1, 144) <= input(36);
output(1, 145) <= input(34);
output(1, 146) <= input(32);
output(1, 147) <= input(0);
output(1, 148) <= input(1);
output(1, 149) <= input(2);
output(1, 150) <= input(3);
output(1, 151) <= input(4);
output(1, 152) <= input(5);
output(1, 153) <= input(6);
output(1, 154) <= input(7);
output(1, 155) <= input(8);
output(1, 156) <= input(9);
output(1, 157) <= input(10);
output(1, 158) <= input(11);
output(1, 159) <= input(12);
output(1, 160) <= input(37);
output(1, 161) <= input(35);
output(1, 162) <= input(33);
output(1, 163) <= input(16);
output(1, 164) <= input(17);
output(1, 165) <= input(18);
output(1, 166) <= input(19);
output(1, 167) <= input(20);
output(1, 168) <= input(21);
output(1, 169) <= input(22);
output(1, 170) <= input(23);
output(1, 171) <= input(24);
output(1, 172) <= input(25);
output(1, 173) <= input(26);
output(1, 174) <= input(27);
output(1, 175) <= input(28);
output(1, 176) <= input(40);
output(1, 177) <= input(36);
output(1, 178) <= input(34);
output(1, 179) <= input(32);
output(1, 180) <= input(0);
output(1, 181) <= input(1);
output(1, 182) <= input(2);
output(1, 183) <= input(3);
output(1, 184) <= input(4);
output(1, 185) <= input(5);
output(1, 186) <= input(6);
output(1, 187) <= input(7);
output(1, 188) <= input(8);
output(1, 189) <= input(9);
output(1, 190) <= input(10);
output(1, 191) <= input(11);
output(1, 192) <= input(38);
output(1, 193) <= input(37);
output(1, 194) <= input(35);
output(1, 195) <= input(33);
output(1, 196) <= input(16);
output(1, 197) <= input(17);
output(1, 198) <= input(18);
output(1, 199) <= input(19);
output(1, 200) <= input(20);
output(1, 201) <= input(21);
output(1, 202) <= input(22);
output(1, 203) <= input(23);
output(1, 204) <= input(24);
output(1, 205) <= input(25);
output(1, 206) <= input(26);
output(1, 207) <= input(27);
output(1, 208) <= input(39);
output(1, 209) <= input(40);
output(1, 210) <= input(36);
output(1, 211) <= input(34);
output(1, 212) <= input(32);
output(1, 213) <= input(0);
output(1, 214) <= input(1);
output(1, 215) <= input(2);
output(1, 216) <= input(3);
output(1, 217) <= input(4);
output(1, 218) <= input(5);
output(1, 219) <= input(6);
output(1, 220) <= input(7);
output(1, 221) <= input(8);
output(1, 222) <= input(9);
output(1, 223) <= input(10);
output(1, 224) <= input(41);
output(1, 225) <= input(38);
output(1, 226) <= input(37);
output(1, 227) <= input(35);
output(1, 228) <= input(33);
output(1, 229) <= input(16);
output(1, 230) <= input(17);
output(1, 231) <= input(18);
output(1, 232) <= input(19);
output(1, 233) <= input(20);
output(1, 234) <= input(21);
output(1, 235) <= input(22);
output(1, 236) <= input(23);
output(1, 237) <= input(24);
output(1, 238) <= input(25);
output(1, 239) <= input(26);
output(1, 240) <= input(42);
output(1, 241) <= input(39);
output(1, 242) <= input(40);
output(1, 243) <= input(36);
output(1, 244) <= input(34);
output(1, 245) <= input(32);
output(1, 246) <= input(0);
output(1, 247) <= input(1);
output(1, 248) <= input(2);
output(1, 249) <= input(3);
output(1, 250) <= input(4);
output(1, 251) <= input(5);
output(1, 252) <= input(6);
output(1, 253) <= input(7);
output(1, 254) <= input(8);
output(1, 255) <= input(9);
when "1011" =>
output(0, 0) <= input(0);
output(0, 1) <= input(1);
output(0, 2) <= input(2);
output(0, 3) <= input(3);
output(0, 4) <= input(4);
output(0, 5) <= input(5);
output(0, 6) <= input(6);
output(0, 7) <= input(7);
output(0, 8) <= input(8);
output(0, 9) <= input(9);
output(0, 10) <= input(10);
output(0, 11) <= input(11);
output(0, 12) <= input(12);
output(0, 13) <= input(13);
output(0, 14) <= input(14);
output(0, 15) <= input(15);
output(0, 16) <= input(16);
output(0, 17) <= input(17);
output(0, 18) <= input(18);
output(0, 19) <= input(19);
output(0, 20) <= input(20);
output(0, 21) <= input(21);
output(0, 22) <= input(22);
output(0, 23) <= input(23);
output(0, 24) <= input(24);
output(0, 25) <= input(25);
output(0, 26) <= input(26);
output(0, 27) <= input(27);
output(0, 28) <= input(28);
output(0, 29) <= input(29);
output(0, 30) <= input(30);
output(0, 31) <= input(31);
output(0, 32) <= input(32);
output(0, 33) <= input(0);
output(0, 34) <= input(1);
output(0, 35) <= input(2);
output(0, 36) <= input(3);
output(0, 37) <= input(4);
output(0, 38) <= input(5);
output(0, 39) <= input(6);
output(0, 40) <= input(7);
output(0, 41) <= input(8);
output(0, 42) <= input(9);
output(0, 43) <= input(10);
output(0, 44) <= input(11);
output(0, 45) <= input(12);
output(0, 46) <= input(13);
output(0, 47) <= input(14);
output(0, 48) <= input(33);
output(0, 49) <= input(16);
output(0, 50) <= input(17);
output(0, 51) <= input(18);
output(0, 52) <= input(19);
output(0, 53) <= input(20);
output(0, 54) <= input(21);
output(0, 55) <= input(22);
output(0, 56) <= input(23);
output(0, 57) <= input(24);
output(0, 58) <= input(25);
output(0, 59) <= input(26);
output(0, 60) <= input(27);
output(0, 61) <= input(28);
output(0, 62) <= input(29);
output(0, 63) <= input(30);
output(0, 64) <= input(34);
output(0, 65) <= input(32);
output(0, 66) <= input(0);
output(0, 67) <= input(1);
output(0, 68) <= input(2);
output(0, 69) <= input(3);
output(0, 70) <= input(4);
output(0, 71) <= input(5);
output(0, 72) <= input(6);
output(0, 73) <= input(7);
output(0, 74) <= input(8);
output(0, 75) <= input(9);
output(0, 76) <= input(10);
output(0, 77) <= input(11);
output(0, 78) <= input(12);
output(0, 79) <= input(13);
output(0, 80) <= input(35);
output(0, 81) <= input(33);
output(0, 82) <= input(16);
output(0, 83) <= input(17);
output(0, 84) <= input(18);
output(0, 85) <= input(19);
output(0, 86) <= input(20);
output(0, 87) <= input(21);
output(0, 88) <= input(22);
output(0, 89) <= input(23);
output(0, 90) <= input(24);
output(0, 91) <= input(25);
output(0, 92) <= input(26);
output(0, 93) <= input(27);
output(0, 94) <= input(28);
output(0, 95) <= input(29);
output(0, 96) <= input(36);
output(0, 97) <= input(34);
output(0, 98) <= input(32);
output(0, 99) <= input(0);
output(0, 100) <= input(1);
output(0, 101) <= input(2);
output(0, 102) <= input(3);
output(0, 103) <= input(4);
output(0, 104) <= input(5);
output(0, 105) <= input(6);
output(0, 106) <= input(7);
output(0, 107) <= input(8);
output(0, 108) <= input(9);
output(0, 109) <= input(10);
output(0, 110) <= input(11);
output(0, 111) <= input(12);
output(0, 112) <= input(36);
output(0, 113) <= input(34);
output(0, 114) <= input(32);
output(0, 115) <= input(0);
output(0, 116) <= input(1);
output(0, 117) <= input(2);
output(0, 118) <= input(3);
output(0, 119) <= input(4);
output(0, 120) <= input(5);
output(0, 121) <= input(6);
output(0, 122) <= input(7);
output(0, 123) <= input(8);
output(0, 124) <= input(9);
output(0, 125) <= input(10);
output(0, 126) <= input(11);
output(0, 127) <= input(12);
output(0, 128) <= input(37);
output(0, 129) <= input(35);
output(0, 130) <= input(33);
output(0, 131) <= input(16);
output(0, 132) <= input(17);
output(0, 133) <= input(18);
output(0, 134) <= input(19);
output(0, 135) <= input(20);
output(0, 136) <= input(21);
output(0, 137) <= input(22);
output(0, 138) <= input(23);
output(0, 139) <= input(24);
output(0, 140) <= input(25);
output(0, 141) <= input(26);
output(0, 142) <= input(27);
output(0, 143) <= input(28);
output(0, 144) <= input(38);
output(0, 145) <= input(36);
output(0, 146) <= input(34);
output(0, 147) <= input(32);
output(0, 148) <= input(0);
output(0, 149) <= input(1);
output(0, 150) <= input(2);
output(0, 151) <= input(3);
output(0, 152) <= input(4);
output(0, 153) <= input(5);
output(0, 154) <= input(6);
output(0, 155) <= input(7);
output(0, 156) <= input(8);
output(0, 157) <= input(9);
output(0, 158) <= input(10);
output(0, 159) <= input(11);
output(0, 160) <= input(39);
output(0, 161) <= input(37);
output(0, 162) <= input(35);
output(0, 163) <= input(33);
output(0, 164) <= input(16);
output(0, 165) <= input(17);
output(0, 166) <= input(18);
output(0, 167) <= input(19);
output(0, 168) <= input(20);
output(0, 169) <= input(21);
output(0, 170) <= input(22);
output(0, 171) <= input(23);
output(0, 172) <= input(24);
output(0, 173) <= input(25);
output(0, 174) <= input(26);
output(0, 175) <= input(27);
output(0, 176) <= input(40);
output(0, 177) <= input(38);
output(0, 178) <= input(36);
output(0, 179) <= input(34);
output(0, 180) <= input(32);
output(0, 181) <= input(0);
output(0, 182) <= input(1);
output(0, 183) <= input(2);
output(0, 184) <= input(3);
output(0, 185) <= input(4);
output(0, 186) <= input(5);
output(0, 187) <= input(6);
output(0, 188) <= input(7);
output(0, 189) <= input(8);
output(0, 190) <= input(9);
output(0, 191) <= input(10);
output(0, 192) <= input(41);
output(0, 193) <= input(39);
output(0, 194) <= input(37);
output(0, 195) <= input(35);
output(0, 196) <= input(33);
output(0, 197) <= input(16);
output(0, 198) <= input(17);
output(0, 199) <= input(18);
output(0, 200) <= input(19);
output(0, 201) <= input(20);
output(0, 202) <= input(21);
output(0, 203) <= input(22);
output(0, 204) <= input(23);
output(0, 205) <= input(24);
output(0, 206) <= input(25);
output(0, 207) <= input(26);
output(0, 208) <= input(42);
output(0, 209) <= input(40);
output(0, 210) <= input(38);
output(0, 211) <= input(36);
output(0, 212) <= input(34);
output(0, 213) <= input(32);
output(0, 214) <= input(0);
output(0, 215) <= input(1);
output(0, 216) <= input(2);
output(0, 217) <= input(3);
output(0, 218) <= input(4);
output(0, 219) <= input(5);
output(0, 220) <= input(6);
output(0, 221) <= input(7);
output(0, 222) <= input(8);
output(0, 223) <= input(9);
output(0, 224) <= input(43);
output(0, 225) <= input(41);
output(0, 226) <= input(39);
output(0, 227) <= input(37);
output(0, 228) <= input(35);
output(0, 229) <= input(33);
output(0, 230) <= input(16);
output(0, 231) <= input(17);
output(0, 232) <= input(18);
output(0, 233) <= input(19);
output(0, 234) <= input(20);
output(0, 235) <= input(21);
output(0, 236) <= input(22);
output(0, 237) <= input(23);
output(0, 238) <= input(24);
output(0, 239) <= input(25);
output(0, 240) <= input(43);
output(0, 241) <= input(41);
output(0, 242) <= input(39);
output(0, 243) <= input(37);
output(0, 244) <= input(35);
output(0, 245) <= input(33);
output(0, 246) <= input(16);
output(0, 247) <= input(17);
output(0, 248) <= input(18);
output(0, 249) <= input(19);
output(0, 250) <= input(20);
output(0, 251) <= input(21);
output(0, 252) <= input(22);
output(0, 253) <= input(23);
output(0, 254) <= input(24);
output(0, 255) <= input(25);
output(1, 0) <= input(1);
output(1, 1) <= input(2);
output(1, 2) <= input(3);
output(1, 3) <= input(4);
output(1, 4) <= input(5);
output(1, 5) <= input(6);
output(1, 6) <= input(7);
output(1, 7) <= input(8);
output(1, 8) <= input(9);
output(1, 9) <= input(10);
output(1, 10) <= input(11);
output(1, 11) <= input(12);
output(1, 12) <= input(13);
output(1, 13) <= input(14);
output(1, 14) <= input(15);
output(1, 15) <= input(44);
output(1, 16) <= input(17);
output(1, 17) <= input(18);
output(1, 18) <= input(19);
output(1, 19) <= input(20);
output(1, 20) <= input(21);
output(1, 21) <= input(22);
output(1, 22) <= input(23);
output(1, 23) <= input(24);
output(1, 24) <= input(25);
output(1, 25) <= input(26);
output(1, 26) <= input(27);
output(1, 27) <= input(28);
output(1, 28) <= input(29);
output(1, 29) <= input(30);
output(1, 30) <= input(31);
output(1, 31) <= input(45);
output(1, 32) <= input(0);
output(1, 33) <= input(1);
output(1, 34) <= input(2);
output(1, 35) <= input(3);
output(1, 36) <= input(4);
output(1, 37) <= input(5);
output(1, 38) <= input(6);
output(1, 39) <= input(7);
output(1, 40) <= input(8);
output(1, 41) <= input(9);
output(1, 42) <= input(10);
output(1, 43) <= input(11);
output(1, 44) <= input(12);
output(1, 45) <= input(13);
output(1, 46) <= input(14);
output(1, 47) <= input(15);
output(1, 48) <= input(0);
output(1, 49) <= input(1);
output(1, 50) <= input(2);
output(1, 51) <= input(3);
output(1, 52) <= input(4);
output(1, 53) <= input(5);
output(1, 54) <= input(6);
output(1, 55) <= input(7);
output(1, 56) <= input(8);
output(1, 57) <= input(9);
output(1, 58) <= input(10);
output(1, 59) <= input(11);
output(1, 60) <= input(12);
output(1, 61) <= input(13);
output(1, 62) <= input(14);
output(1, 63) <= input(15);
output(1, 64) <= input(16);
output(1, 65) <= input(17);
output(1, 66) <= input(18);
output(1, 67) <= input(19);
output(1, 68) <= input(20);
output(1, 69) <= input(21);
output(1, 70) <= input(22);
output(1, 71) <= input(23);
output(1, 72) <= input(24);
output(1, 73) <= input(25);
output(1, 74) <= input(26);
output(1, 75) <= input(27);
output(1, 76) <= input(28);
output(1, 77) <= input(29);
output(1, 78) <= input(30);
output(1, 79) <= input(31);
output(1, 80) <= input(32);
output(1, 81) <= input(0);
output(1, 82) <= input(1);
output(1, 83) <= input(2);
output(1, 84) <= input(3);
output(1, 85) <= input(4);
output(1, 86) <= input(5);
output(1, 87) <= input(6);
output(1, 88) <= input(7);
output(1, 89) <= input(8);
output(1, 90) <= input(9);
output(1, 91) <= input(10);
output(1, 92) <= input(11);
output(1, 93) <= input(12);
output(1, 94) <= input(13);
output(1, 95) <= input(14);
output(1, 96) <= input(33);
output(1, 97) <= input(16);
output(1, 98) <= input(17);
output(1, 99) <= input(18);
output(1, 100) <= input(19);
output(1, 101) <= input(20);
output(1, 102) <= input(21);
output(1, 103) <= input(22);
output(1, 104) <= input(23);
output(1, 105) <= input(24);
output(1, 106) <= input(25);
output(1, 107) <= input(26);
output(1, 108) <= input(27);
output(1, 109) <= input(28);
output(1, 110) <= input(29);
output(1, 111) <= input(30);
output(1, 112) <= input(33);
output(1, 113) <= input(16);
output(1, 114) <= input(17);
output(1, 115) <= input(18);
output(1, 116) <= input(19);
output(1, 117) <= input(20);
output(1, 118) <= input(21);
output(1, 119) <= input(22);
output(1, 120) <= input(23);
output(1, 121) <= input(24);
output(1, 122) <= input(25);
output(1, 123) <= input(26);
output(1, 124) <= input(27);
output(1, 125) <= input(28);
output(1, 126) <= input(29);
output(1, 127) <= input(30);
output(1, 128) <= input(34);
output(1, 129) <= input(32);
output(1, 130) <= input(0);
output(1, 131) <= input(1);
output(1, 132) <= input(2);
output(1, 133) <= input(3);
output(1, 134) <= input(4);
output(1, 135) <= input(5);
output(1, 136) <= input(6);
output(1, 137) <= input(7);
output(1, 138) <= input(8);
output(1, 139) <= input(9);
output(1, 140) <= input(10);
output(1, 141) <= input(11);
output(1, 142) <= input(12);
output(1, 143) <= input(13);
output(1, 144) <= input(35);
output(1, 145) <= input(33);
output(1, 146) <= input(16);
output(1, 147) <= input(17);
output(1, 148) <= input(18);
output(1, 149) <= input(19);
output(1, 150) <= input(20);
output(1, 151) <= input(21);
output(1, 152) <= input(22);
output(1, 153) <= input(23);
output(1, 154) <= input(24);
output(1, 155) <= input(25);
output(1, 156) <= input(26);
output(1, 157) <= input(27);
output(1, 158) <= input(28);
output(1, 159) <= input(29);
output(1, 160) <= input(36);
output(1, 161) <= input(34);
output(1, 162) <= input(32);
output(1, 163) <= input(0);
output(1, 164) <= input(1);
output(1, 165) <= input(2);
output(1, 166) <= input(3);
output(1, 167) <= input(4);
output(1, 168) <= input(5);
output(1, 169) <= input(6);
output(1, 170) <= input(7);
output(1, 171) <= input(8);
output(1, 172) <= input(9);
output(1, 173) <= input(10);
output(1, 174) <= input(11);
output(1, 175) <= input(12);
output(1, 176) <= input(36);
output(1, 177) <= input(34);
output(1, 178) <= input(32);
output(1, 179) <= input(0);
output(1, 180) <= input(1);
output(1, 181) <= input(2);
output(1, 182) <= input(3);
output(1, 183) <= input(4);
output(1, 184) <= input(5);
output(1, 185) <= input(6);
output(1, 186) <= input(7);
output(1, 187) <= input(8);
output(1, 188) <= input(9);
output(1, 189) <= input(10);
output(1, 190) <= input(11);
output(1, 191) <= input(12);
output(1, 192) <= input(37);
output(1, 193) <= input(35);
output(1, 194) <= input(33);
output(1, 195) <= input(16);
output(1, 196) <= input(17);
output(1, 197) <= input(18);
output(1, 198) <= input(19);
output(1, 199) <= input(20);
output(1, 200) <= input(21);
output(1, 201) <= input(22);
output(1, 202) <= input(23);
output(1, 203) <= input(24);
output(1, 204) <= input(25);
output(1, 205) <= input(26);
output(1, 206) <= input(27);
output(1, 207) <= input(28);
output(1, 208) <= input(38);
output(1, 209) <= input(36);
output(1, 210) <= input(34);
output(1, 211) <= input(32);
output(1, 212) <= input(0);
output(1, 213) <= input(1);
output(1, 214) <= input(2);
output(1, 215) <= input(3);
output(1, 216) <= input(4);
output(1, 217) <= input(5);
output(1, 218) <= input(6);
output(1, 219) <= input(7);
output(1, 220) <= input(8);
output(1, 221) <= input(9);
output(1, 222) <= input(10);
output(1, 223) <= input(11);
output(1, 224) <= input(39);
output(1, 225) <= input(37);
output(1, 226) <= input(35);
output(1, 227) <= input(33);
output(1, 228) <= input(16);
output(1, 229) <= input(17);
output(1, 230) <= input(18);
output(1, 231) <= input(19);
output(1, 232) <= input(20);
output(1, 233) <= input(21);
output(1, 234) <= input(22);
output(1, 235) <= input(23);
output(1, 236) <= input(24);
output(1, 237) <= input(25);
output(1, 238) <= input(26);
output(1, 239) <= input(27);
output(1, 240) <= input(39);
output(1, 241) <= input(37);
output(1, 242) <= input(35);
output(1, 243) <= input(33);
output(1, 244) <= input(16);
output(1, 245) <= input(17);
output(1, 246) <= input(18);
output(1, 247) <= input(19);
output(1, 248) <= input(20);
output(1, 249) <= input(21);
output(1, 250) <= input(22);
output(1, 251) <= input(23);
output(1, 252) <= input(24);
output(1, 253) <= input(25);
output(1, 254) <= input(26);
output(1, 255) <= input(27);
output(2, 0) <= input(2);
output(2, 1) <= input(3);
output(2, 2) <= input(4);
output(2, 3) <= input(5);
output(2, 4) <= input(6);
output(2, 5) <= input(7);
output(2, 6) <= input(8);
output(2, 7) <= input(9);
output(2, 8) <= input(10);
output(2, 9) <= input(11);
output(2, 10) <= input(12);
output(2, 11) <= input(13);
output(2, 12) <= input(14);
output(2, 13) <= input(15);
output(2, 14) <= input(44);
output(2, 15) <= input(46);
output(2, 16) <= input(18);
output(2, 17) <= input(19);
output(2, 18) <= input(20);
output(2, 19) <= input(21);
output(2, 20) <= input(22);
output(2, 21) <= input(23);
output(2, 22) <= input(24);
output(2, 23) <= input(25);
output(2, 24) <= input(26);
output(2, 25) <= input(27);
output(2, 26) <= input(28);
output(2, 27) <= input(29);
output(2, 28) <= input(30);
output(2, 29) <= input(31);
output(2, 30) <= input(45);
output(2, 31) <= input(47);
output(2, 32) <= input(18);
output(2, 33) <= input(19);
output(2, 34) <= input(20);
output(2, 35) <= input(21);
output(2, 36) <= input(22);
output(2, 37) <= input(23);
output(2, 38) <= input(24);
output(2, 39) <= input(25);
output(2, 40) <= input(26);
output(2, 41) <= input(27);
output(2, 42) <= input(28);
output(2, 43) <= input(29);
output(2, 44) <= input(30);
output(2, 45) <= input(31);
output(2, 46) <= input(45);
output(2, 47) <= input(47);
output(2, 48) <= input(1);
output(2, 49) <= input(2);
output(2, 50) <= input(3);
output(2, 51) <= input(4);
output(2, 52) <= input(5);
output(2, 53) <= input(6);
output(2, 54) <= input(7);
output(2, 55) <= input(8);
output(2, 56) <= input(9);
output(2, 57) <= input(10);
output(2, 58) <= input(11);
output(2, 59) <= input(12);
output(2, 60) <= input(13);
output(2, 61) <= input(14);
output(2, 62) <= input(15);
output(2, 63) <= input(44);
output(2, 64) <= input(17);
output(2, 65) <= input(18);
output(2, 66) <= input(19);
output(2, 67) <= input(20);
output(2, 68) <= input(21);
output(2, 69) <= input(22);
output(2, 70) <= input(23);
output(2, 71) <= input(24);
output(2, 72) <= input(25);
output(2, 73) <= input(26);
output(2, 74) <= input(27);
output(2, 75) <= input(28);
output(2, 76) <= input(29);
output(2, 77) <= input(30);
output(2, 78) <= input(31);
output(2, 79) <= input(45);
output(2, 80) <= input(17);
output(2, 81) <= input(18);
output(2, 82) <= input(19);
output(2, 83) <= input(20);
output(2, 84) <= input(21);
output(2, 85) <= input(22);
output(2, 86) <= input(23);
output(2, 87) <= input(24);
output(2, 88) <= input(25);
output(2, 89) <= input(26);
output(2, 90) <= input(27);
output(2, 91) <= input(28);
output(2, 92) <= input(29);
output(2, 93) <= input(30);
output(2, 94) <= input(31);
output(2, 95) <= input(45);
output(2, 96) <= input(0);
output(2, 97) <= input(1);
output(2, 98) <= input(2);
output(2, 99) <= input(3);
output(2, 100) <= input(4);
output(2, 101) <= input(5);
output(2, 102) <= input(6);
output(2, 103) <= input(7);
output(2, 104) <= input(8);
output(2, 105) <= input(9);
output(2, 106) <= input(10);
output(2, 107) <= input(11);
output(2, 108) <= input(12);
output(2, 109) <= input(13);
output(2, 110) <= input(14);
output(2, 111) <= input(15);
output(2, 112) <= input(0);
output(2, 113) <= input(1);
output(2, 114) <= input(2);
output(2, 115) <= input(3);
output(2, 116) <= input(4);
output(2, 117) <= input(5);
output(2, 118) <= input(6);
output(2, 119) <= input(7);
output(2, 120) <= input(8);
output(2, 121) <= input(9);
output(2, 122) <= input(10);
output(2, 123) <= input(11);
output(2, 124) <= input(12);
output(2, 125) <= input(13);
output(2, 126) <= input(14);
output(2, 127) <= input(15);
output(2, 128) <= input(16);
output(2, 129) <= input(17);
output(2, 130) <= input(18);
output(2, 131) <= input(19);
output(2, 132) <= input(20);
output(2, 133) <= input(21);
output(2, 134) <= input(22);
output(2, 135) <= input(23);
output(2, 136) <= input(24);
output(2, 137) <= input(25);
output(2, 138) <= input(26);
output(2, 139) <= input(27);
output(2, 140) <= input(28);
output(2, 141) <= input(29);
output(2, 142) <= input(30);
output(2, 143) <= input(31);
output(2, 144) <= input(32);
output(2, 145) <= input(0);
output(2, 146) <= input(1);
output(2, 147) <= input(2);
output(2, 148) <= input(3);
output(2, 149) <= input(4);
output(2, 150) <= input(5);
output(2, 151) <= input(6);
output(2, 152) <= input(7);
output(2, 153) <= input(8);
output(2, 154) <= input(9);
output(2, 155) <= input(10);
output(2, 156) <= input(11);
output(2, 157) <= input(12);
output(2, 158) <= input(13);
output(2, 159) <= input(14);
output(2, 160) <= input(32);
output(2, 161) <= input(0);
output(2, 162) <= input(1);
output(2, 163) <= input(2);
output(2, 164) <= input(3);
output(2, 165) <= input(4);
output(2, 166) <= input(5);
output(2, 167) <= input(6);
output(2, 168) <= input(7);
output(2, 169) <= input(8);
output(2, 170) <= input(9);
output(2, 171) <= input(10);
output(2, 172) <= input(11);
output(2, 173) <= input(12);
output(2, 174) <= input(13);
output(2, 175) <= input(14);
output(2, 176) <= input(33);
output(2, 177) <= input(16);
output(2, 178) <= input(17);
output(2, 179) <= input(18);
output(2, 180) <= input(19);
output(2, 181) <= input(20);
output(2, 182) <= input(21);
output(2, 183) <= input(22);
output(2, 184) <= input(23);
output(2, 185) <= input(24);
output(2, 186) <= input(25);
output(2, 187) <= input(26);
output(2, 188) <= input(27);
output(2, 189) <= input(28);
output(2, 190) <= input(29);
output(2, 191) <= input(30);
output(2, 192) <= input(34);
output(2, 193) <= input(32);
output(2, 194) <= input(0);
output(2, 195) <= input(1);
output(2, 196) <= input(2);
output(2, 197) <= input(3);
output(2, 198) <= input(4);
output(2, 199) <= input(5);
output(2, 200) <= input(6);
output(2, 201) <= input(7);
output(2, 202) <= input(8);
output(2, 203) <= input(9);
output(2, 204) <= input(10);
output(2, 205) <= input(11);
output(2, 206) <= input(12);
output(2, 207) <= input(13);
output(2, 208) <= input(34);
output(2, 209) <= input(32);
output(2, 210) <= input(0);
output(2, 211) <= input(1);
output(2, 212) <= input(2);
output(2, 213) <= input(3);
output(2, 214) <= input(4);
output(2, 215) <= input(5);
output(2, 216) <= input(6);
output(2, 217) <= input(7);
output(2, 218) <= input(8);
output(2, 219) <= input(9);
output(2, 220) <= input(10);
output(2, 221) <= input(11);
output(2, 222) <= input(12);
output(2, 223) <= input(13);
output(2, 224) <= input(35);
output(2, 225) <= input(33);
output(2, 226) <= input(16);
output(2, 227) <= input(17);
output(2, 228) <= input(18);
output(2, 229) <= input(19);
output(2, 230) <= input(20);
output(2, 231) <= input(21);
output(2, 232) <= input(22);
output(2, 233) <= input(23);
output(2, 234) <= input(24);
output(2, 235) <= input(25);
output(2, 236) <= input(26);
output(2, 237) <= input(27);
output(2, 238) <= input(28);
output(2, 239) <= input(29);
output(2, 240) <= input(35);
output(2, 241) <= input(33);
output(2, 242) <= input(16);
output(2, 243) <= input(17);
output(2, 244) <= input(18);
output(2, 245) <= input(19);
output(2, 246) <= input(20);
output(2, 247) <= input(21);
output(2, 248) <= input(22);
output(2, 249) <= input(23);
output(2, 250) <= input(24);
output(2, 251) <= input(25);
output(2, 252) <= input(26);
output(2, 253) <= input(27);
output(2, 254) <= input(28);
output(2, 255) <= input(29);
when "1100" =>
output(0, 0) <= input(0);
output(0, 1) <= input(1);
output(0, 2) <= input(2);
output(0, 3) <= input(3);
output(0, 4) <= input(4);
output(0, 5) <= input(5);
output(0, 6) <= input(6);
output(0, 7) <= input(7);
output(0, 8) <= input(8);
output(0, 9) <= input(9);
output(0, 10) <= input(10);
output(0, 11) <= input(11);
output(0, 12) <= input(12);
output(0, 13) <= input(13);
output(0, 14) <= input(14);
output(0, 15) <= input(15);
output(0, 16) <= input(0);
output(0, 17) <= input(1);
output(0, 18) <= input(2);
output(0, 19) <= input(3);
output(0, 20) <= input(4);
output(0, 21) <= input(5);
output(0, 22) <= input(6);
output(0, 23) <= input(7);
output(0, 24) <= input(8);
output(0, 25) <= input(9);
output(0, 26) <= input(10);
output(0, 27) <= input(11);
output(0, 28) <= input(12);
output(0, 29) <= input(13);
output(0, 30) <= input(14);
output(0, 31) <= input(15);
output(0, 32) <= input(16);
output(0, 33) <= input(17);
output(0, 34) <= input(18);
output(0, 35) <= input(19);
output(0, 36) <= input(20);
output(0, 37) <= input(21);
output(0, 38) <= input(22);
output(0, 39) <= input(23);
output(0, 40) <= input(24);
output(0, 41) <= input(25);
output(0, 42) <= input(26);
output(0, 43) <= input(27);
output(0, 44) <= input(28);
output(0, 45) <= input(29);
output(0, 46) <= input(30);
output(0, 47) <= input(31);
output(0, 48) <= input(16);
output(0, 49) <= input(17);
output(0, 50) <= input(18);
output(0, 51) <= input(19);
output(0, 52) <= input(20);
output(0, 53) <= input(21);
output(0, 54) <= input(22);
output(0, 55) <= input(23);
output(0, 56) <= input(24);
output(0, 57) <= input(25);
output(0, 58) <= input(26);
output(0, 59) <= input(27);
output(0, 60) <= input(28);
output(0, 61) <= input(29);
output(0, 62) <= input(30);
output(0, 63) <= input(31);
output(0, 64) <= input(32);
output(0, 65) <= input(0);
output(0, 66) <= input(1);
output(0, 67) <= input(2);
output(0, 68) <= input(3);
output(0, 69) <= input(4);
output(0, 70) <= input(5);
output(0, 71) <= input(6);
output(0, 72) <= input(7);
output(0, 73) <= input(8);
output(0, 74) <= input(9);
output(0, 75) <= input(10);
output(0, 76) <= input(11);
output(0, 77) <= input(12);
output(0, 78) <= input(13);
output(0, 79) <= input(14);
output(0, 80) <= input(32);
output(0, 81) <= input(0);
output(0, 82) <= input(1);
output(0, 83) <= input(2);
output(0, 84) <= input(3);
output(0, 85) <= input(4);
output(0, 86) <= input(5);
output(0, 87) <= input(6);
output(0, 88) <= input(7);
output(0, 89) <= input(8);
output(0, 90) <= input(9);
output(0, 91) <= input(10);
output(0, 92) <= input(11);
output(0, 93) <= input(12);
output(0, 94) <= input(13);
output(0, 95) <= input(14);
output(0, 96) <= input(33);
output(0, 97) <= input(16);
output(0, 98) <= input(17);
output(0, 99) <= input(18);
output(0, 100) <= input(19);
output(0, 101) <= input(20);
output(0, 102) <= input(21);
output(0, 103) <= input(22);
output(0, 104) <= input(23);
output(0, 105) <= input(24);
output(0, 106) <= input(25);
output(0, 107) <= input(26);
output(0, 108) <= input(27);
output(0, 109) <= input(28);
output(0, 110) <= input(29);
output(0, 111) <= input(30);
output(0, 112) <= input(33);
output(0, 113) <= input(16);
output(0, 114) <= input(17);
output(0, 115) <= input(18);
output(0, 116) <= input(19);
output(0, 117) <= input(20);
output(0, 118) <= input(21);
output(0, 119) <= input(22);
output(0, 120) <= input(23);
output(0, 121) <= input(24);
output(0, 122) <= input(25);
output(0, 123) <= input(26);
output(0, 124) <= input(27);
output(0, 125) <= input(28);
output(0, 126) <= input(29);
output(0, 127) <= input(30);
output(0, 128) <= input(34);
output(0, 129) <= input(32);
output(0, 130) <= input(0);
output(0, 131) <= input(1);
output(0, 132) <= input(2);
output(0, 133) <= input(3);
output(0, 134) <= input(4);
output(0, 135) <= input(5);
output(0, 136) <= input(6);
output(0, 137) <= input(7);
output(0, 138) <= input(8);
output(0, 139) <= input(9);
output(0, 140) <= input(10);
output(0, 141) <= input(11);
output(0, 142) <= input(12);
output(0, 143) <= input(13);
output(0, 144) <= input(34);
output(0, 145) <= input(32);
output(0, 146) <= input(0);
output(0, 147) <= input(1);
output(0, 148) <= input(2);
output(0, 149) <= input(3);
output(0, 150) <= input(4);
output(0, 151) <= input(5);
output(0, 152) <= input(6);
output(0, 153) <= input(7);
output(0, 154) <= input(8);
output(0, 155) <= input(9);
output(0, 156) <= input(10);
output(0, 157) <= input(11);
output(0, 158) <= input(12);
output(0, 159) <= input(13);
output(0, 160) <= input(35);
output(0, 161) <= input(33);
output(0, 162) <= input(16);
output(0, 163) <= input(17);
output(0, 164) <= input(18);
output(0, 165) <= input(19);
output(0, 166) <= input(20);
output(0, 167) <= input(21);
output(0, 168) <= input(22);
output(0, 169) <= input(23);
output(0, 170) <= input(24);
output(0, 171) <= input(25);
output(0, 172) <= input(26);
output(0, 173) <= input(27);
output(0, 174) <= input(28);
output(0, 175) <= input(29);
output(0, 176) <= input(35);
output(0, 177) <= input(33);
output(0, 178) <= input(16);
output(0, 179) <= input(17);
output(0, 180) <= input(18);
output(0, 181) <= input(19);
output(0, 182) <= input(20);
output(0, 183) <= input(21);
output(0, 184) <= input(22);
output(0, 185) <= input(23);
output(0, 186) <= input(24);
output(0, 187) <= input(25);
output(0, 188) <= input(26);
output(0, 189) <= input(27);
output(0, 190) <= input(28);
output(0, 191) <= input(29);
output(0, 192) <= input(36);
output(0, 193) <= input(34);
output(0, 194) <= input(32);
output(0, 195) <= input(0);
output(0, 196) <= input(1);
output(0, 197) <= input(2);
output(0, 198) <= input(3);
output(0, 199) <= input(4);
output(0, 200) <= input(5);
output(0, 201) <= input(6);
output(0, 202) <= input(7);
output(0, 203) <= input(8);
output(0, 204) <= input(9);
output(0, 205) <= input(10);
output(0, 206) <= input(11);
output(0, 207) <= input(12);
output(0, 208) <= input(36);
output(0, 209) <= input(34);
output(0, 210) <= input(32);
output(0, 211) <= input(0);
output(0, 212) <= input(1);
output(0, 213) <= input(2);
output(0, 214) <= input(3);
output(0, 215) <= input(4);
output(0, 216) <= input(5);
output(0, 217) <= input(6);
output(0, 218) <= input(7);
output(0, 219) <= input(8);
output(0, 220) <= input(9);
output(0, 221) <= input(10);
output(0, 222) <= input(11);
output(0, 223) <= input(12);
output(0, 224) <= input(37);
output(0, 225) <= input(35);
output(0, 226) <= input(33);
output(0, 227) <= input(16);
output(0, 228) <= input(17);
output(0, 229) <= input(18);
output(0, 230) <= input(19);
output(0, 231) <= input(20);
output(0, 232) <= input(21);
output(0, 233) <= input(22);
output(0, 234) <= input(23);
output(0, 235) <= input(24);
output(0, 236) <= input(25);
output(0, 237) <= input(26);
output(0, 238) <= input(27);
output(0, 239) <= input(28);
output(0, 240) <= input(37);
output(0, 241) <= input(35);
output(0, 242) <= input(33);
output(0, 243) <= input(16);
output(0, 244) <= input(17);
output(0, 245) <= input(18);
output(0, 246) <= input(19);
output(0, 247) <= input(20);
output(0, 248) <= input(21);
output(0, 249) <= input(22);
output(0, 250) <= input(23);
output(0, 251) <= input(24);
output(0, 252) <= input(25);
output(0, 253) <= input(26);
output(0, 254) <= input(27);
output(0, 255) <= input(28);
output(1, 0) <= input(1);
output(1, 1) <= input(2);
output(1, 2) <= input(3);
output(1, 3) <= input(4);
output(1, 4) <= input(5);
output(1, 5) <= input(6);
output(1, 6) <= input(7);
output(1, 7) <= input(8);
output(1, 8) <= input(9);
output(1, 9) <= input(10);
output(1, 10) <= input(11);
output(1, 11) <= input(12);
output(1, 12) <= input(13);
output(1, 13) <= input(14);
output(1, 14) <= input(15);
output(1, 15) <= input(38);
output(1, 16) <= input(1);
output(1, 17) <= input(2);
output(1, 18) <= input(3);
output(1, 19) <= input(4);
output(1, 20) <= input(5);
output(1, 21) <= input(6);
output(1, 22) <= input(7);
output(1, 23) <= input(8);
output(1, 24) <= input(9);
output(1, 25) <= input(10);
output(1, 26) <= input(11);
output(1, 27) <= input(12);
output(1, 28) <= input(13);
output(1, 29) <= input(14);
output(1, 30) <= input(15);
output(1, 31) <= input(38);
output(1, 32) <= input(17);
output(1, 33) <= input(18);
output(1, 34) <= input(19);
output(1, 35) <= input(20);
output(1, 36) <= input(21);
output(1, 37) <= input(22);
output(1, 38) <= input(23);
output(1, 39) <= input(24);
output(1, 40) <= input(25);
output(1, 41) <= input(26);
output(1, 42) <= input(27);
output(1, 43) <= input(28);
output(1, 44) <= input(29);
output(1, 45) <= input(30);
output(1, 46) <= input(31);
output(1, 47) <= input(39);
output(1, 48) <= input(17);
output(1, 49) <= input(18);
output(1, 50) <= input(19);
output(1, 51) <= input(20);
output(1, 52) <= input(21);
output(1, 53) <= input(22);
output(1, 54) <= input(23);
output(1, 55) <= input(24);
output(1, 56) <= input(25);
output(1, 57) <= input(26);
output(1, 58) <= input(27);
output(1, 59) <= input(28);
output(1, 60) <= input(29);
output(1, 61) <= input(30);
output(1, 62) <= input(31);
output(1, 63) <= input(39);
output(1, 64) <= input(17);
output(1, 65) <= input(18);
output(1, 66) <= input(19);
output(1, 67) <= input(20);
output(1, 68) <= input(21);
output(1, 69) <= input(22);
output(1, 70) <= input(23);
output(1, 71) <= input(24);
output(1, 72) <= input(25);
output(1, 73) <= input(26);
output(1, 74) <= input(27);
output(1, 75) <= input(28);
output(1, 76) <= input(29);
output(1, 77) <= input(30);
output(1, 78) <= input(31);
output(1, 79) <= input(39);
output(1, 80) <= input(0);
output(1, 81) <= input(1);
output(1, 82) <= input(2);
output(1, 83) <= input(3);
output(1, 84) <= input(4);
output(1, 85) <= input(5);
output(1, 86) <= input(6);
output(1, 87) <= input(7);
output(1, 88) <= input(8);
output(1, 89) <= input(9);
output(1, 90) <= input(10);
output(1, 91) <= input(11);
output(1, 92) <= input(12);
output(1, 93) <= input(13);
output(1, 94) <= input(14);
output(1, 95) <= input(15);
output(1, 96) <= input(0);
output(1, 97) <= input(1);
output(1, 98) <= input(2);
output(1, 99) <= input(3);
output(1, 100) <= input(4);
output(1, 101) <= input(5);
output(1, 102) <= input(6);
output(1, 103) <= input(7);
output(1, 104) <= input(8);
output(1, 105) <= input(9);
output(1, 106) <= input(10);
output(1, 107) <= input(11);
output(1, 108) <= input(12);
output(1, 109) <= input(13);
output(1, 110) <= input(14);
output(1, 111) <= input(15);
output(1, 112) <= input(0);
output(1, 113) <= input(1);
output(1, 114) <= input(2);
output(1, 115) <= input(3);
output(1, 116) <= input(4);
output(1, 117) <= input(5);
output(1, 118) <= input(6);
output(1, 119) <= input(7);
output(1, 120) <= input(8);
output(1, 121) <= input(9);
output(1, 122) <= input(10);
output(1, 123) <= input(11);
output(1, 124) <= input(12);
output(1, 125) <= input(13);
output(1, 126) <= input(14);
output(1, 127) <= input(15);
output(1, 128) <= input(16);
output(1, 129) <= input(17);
output(1, 130) <= input(18);
output(1, 131) <= input(19);
output(1, 132) <= input(20);
output(1, 133) <= input(21);
output(1, 134) <= input(22);
output(1, 135) <= input(23);
output(1, 136) <= input(24);
output(1, 137) <= input(25);
output(1, 138) <= input(26);
output(1, 139) <= input(27);
output(1, 140) <= input(28);
output(1, 141) <= input(29);
output(1, 142) <= input(30);
output(1, 143) <= input(31);
output(1, 144) <= input(16);
output(1, 145) <= input(17);
output(1, 146) <= input(18);
output(1, 147) <= input(19);
output(1, 148) <= input(20);
output(1, 149) <= input(21);
output(1, 150) <= input(22);
output(1, 151) <= input(23);
output(1, 152) <= input(24);
output(1, 153) <= input(25);
output(1, 154) <= input(26);
output(1, 155) <= input(27);
output(1, 156) <= input(28);
output(1, 157) <= input(29);
output(1, 158) <= input(30);
output(1, 159) <= input(31);
output(1, 160) <= input(32);
output(1, 161) <= input(0);
output(1, 162) <= input(1);
output(1, 163) <= input(2);
output(1, 164) <= input(3);
output(1, 165) <= input(4);
output(1, 166) <= input(5);
output(1, 167) <= input(6);
output(1, 168) <= input(7);
output(1, 169) <= input(8);
output(1, 170) <= input(9);
output(1, 171) <= input(10);
output(1, 172) <= input(11);
output(1, 173) <= input(12);
output(1, 174) <= input(13);
output(1, 175) <= input(14);
output(1, 176) <= input(32);
output(1, 177) <= input(0);
output(1, 178) <= input(1);
output(1, 179) <= input(2);
output(1, 180) <= input(3);
output(1, 181) <= input(4);
output(1, 182) <= input(5);
output(1, 183) <= input(6);
output(1, 184) <= input(7);
output(1, 185) <= input(8);
output(1, 186) <= input(9);
output(1, 187) <= input(10);
output(1, 188) <= input(11);
output(1, 189) <= input(12);
output(1, 190) <= input(13);
output(1, 191) <= input(14);
output(1, 192) <= input(32);
output(1, 193) <= input(0);
output(1, 194) <= input(1);
output(1, 195) <= input(2);
output(1, 196) <= input(3);
output(1, 197) <= input(4);
output(1, 198) <= input(5);
output(1, 199) <= input(6);
output(1, 200) <= input(7);
output(1, 201) <= input(8);
output(1, 202) <= input(9);
output(1, 203) <= input(10);
output(1, 204) <= input(11);
output(1, 205) <= input(12);
output(1, 206) <= input(13);
output(1, 207) <= input(14);
output(1, 208) <= input(33);
output(1, 209) <= input(16);
output(1, 210) <= input(17);
output(1, 211) <= input(18);
output(1, 212) <= input(19);
output(1, 213) <= input(20);
output(1, 214) <= input(21);
output(1, 215) <= input(22);
output(1, 216) <= input(23);
output(1, 217) <= input(24);
output(1, 218) <= input(25);
output(1, 219) <= input(26);
output(1, 220) <= input(27);
output(1, 221) <= input(28);
output(1, 222) <= input(29);
output(1, 223) <= input(30);
output(1, 224) <= input(33);
output(1, 225) <= input(16);
output(1, 226) <= input(17);
output(1, 227) <= input(18);
output(1, 228) <= input(19);
output(1, 229) <= input(20);
output(1, 230) <= input(21);
output(1, 231) <= input(22);
output(1, 232) <= input(23);
output(1, 233) <= input(24);
output(1, 234) <= input(25);
output(1, 235) <= input(26);
output(1, 236) <= input(27);
output(1, 237) <= input(28);
output(1, 238) <= input(29);
output(1, 239) <= input(30);
output(1, 240) <= input(33);
output(1, 241) <= input(16);
output(1, 242) <= input(17);
output(1, 243) <= input(18);
output(1, 244) <= input(19);
output(1, 245) <= input(20);
output(1, 246) <= input(21);
output(1, 247) <= input(22);
output(1, 248) <= input(23);
output(1, 249) <= input(24);
output(1, 250) <= input(25);
output(1, 251) <= input(26);
output(1, 252) <= input(27);
output(1, 253) <= input(28);
output(1, 254) <= input(29);
output(1, 255) <= input(30);
output(2, 0) <= input(2);
output(2, 1) <= input(3);
output(2, 2) <= input(4);
output(2, 3) <= input(5);
output(2, 4) <= input(6);
output(2, 5) <= input(7);
output(2, 6) <= input(8);
output(2, 7) <= input(9);
output(2, 8) <= input(10);
output(2, 9) <= input(11);
output(2, 10) <= input(12);
output(2, 11) <= input(13);
output(2, 12) <= input(14);
output(2, 13) <= input(15);
output(2, 14) <= input(38);
output(2, 15) <= input(40);
output(2, 16) <= input(2);
output(2, 17) <= input(3);
output(2, 18) <= input(4);
output(2, 19) <= input(5);
output(2, 20) <= input(6);
output(2, 21) <= input(7);
output(2, 22) <= input(8);
output(2, 23) <= input(9);
output(2, 24) <= input(10);
output(2, 25) <= input(11);
output(2, 26) <= input(12);
output(2, 27) <= input(13);
output(2, 28) <= input(14);
output(2, 29) <= input(15);
output(2, 30) <= input(38);
output(2, 31) <= input(40);
output(2, 32) <= input(2);
output(2, 33) <= input(3);
output(2, 34) <= input(4);
output(2, 35) <= input(5);
output(2, 36) <= input(6);
output(2, 37) <= input(7);
output(2, 38) <= input(8);
output(2, 39) <= input(9);
output(2, 40) <= input(10);
output(2, 41) <= input(11);
output(2, 42) <= input(12);
output(2, 43) <= input(13);
output(2, 44) <= input(14);
output(2, 45) <= input(15);
output(2, 46) <= input(38);
output(2, 47) <= input(40);
output(2, 48) <= input(2);
output(2, 49) <= input(3);
output(2, 50) <= input(4);
output(2, 51) <= input(5);
output(2, 52) <= input(6);
output(2, 53) <= input(7);
output(2, 54) <= input(8);
output(2, 55) <= input(9);
output(2, 56) <= input(10);
output(2, 57) <= input(11);
output(2, 58) <= input(12);
output(2, 59) <= input(13);
output(2, 60) <= input(14);
output(2, 61) <= input(15);
output(2, 62) <= input(38);
output(2, 63) <= input(40);
output(2, 64) <= input(18);
output(2, 65) <= input(19);
output(2, 66) <= input(20);
output(2, 67) <= input(21);
output(2, 68) <= input(22);
output(2, 69) <= input(23);
output(2, 70) <= input(24);
output(2, 71) <= input(25);
output(2, 72) <= input(26);
output(2, 73) <= input(27);
output(2, 74) <= input(28);
output(2, 75) <= input(29);
output(2, 76) <= input(30);
output(2, 77) <= input(31);
output(2, 78) <= input(39);
output(2, 79) <= input(41);
output(2, 80) <= input(18);
output(2, 81) <= input(19);
output(2, 82) <= input(20);
output(2, 83) <= input(21);
output(2, 84) <= input(22);
output(2, 85) <= input(23);
output(2, 86) <= input(24);
output(2, 87) <= input(25);
output(2, 88) <= input(26);
output(2, 89) <= input(27);
output(2, 90) <= input(28);
output(2, 91) <= input(29);
output(2, 92) <= input(30);
output(2, 93) <= input(31);
output(2, 94) <= input(39);
output(2, 95) <= input(41);
output(2, 96) <= input(18);
output(2, 97) <= input(19);
output(2, 98) <= input(20);
output(2, 99) <= input(21);
output(2, 100) <= input(22);
output(2, 101) <= input(23);
output(2, 102) <= input(24);
output(2, 103) <= input(25);
output(2, 104) <= input(26);
output(2, 105) <= input(27);
output(2, 106) <= input(28);
output(2, 107) <= input(29);
output(2, 108) <= input(30);
output(2, 109) <= input(31);
output(2, 110) <= input(39);
output(2, 111) <= input(41);
output(2, 112) <= input(18);
output(2, 113) <= input(19);
output(2, 114) <= input(20);
output(2, 115) <= input(21);
output(2, 116) <= input(22);
output(2, 117) <= input(23);
output(2, 118) <= input(24);
output(2, 119) <= input(25);
output(2, 120) <= input(26);
output(2, 121) <= input(27);
output(2, 122) <= input(28);
output(2, 123) <= input(29);
output(2, 124) <= input(30);
output(2, 125) <= input(31);
output(2, 126) <= input(39);
output(2, 127) <= input(41);
output(2, 128) <= input(1);
output(2, 129) <= input(2);
output(2, 130) <= input(3);
output(2, 131) <= input(4);
output(2, 132) <= input(5);
output(2, 133) <= input(6);
output(2, 134) <= input(7);
output(2, 135) <= input(8);
output(2, 136) <= input(9);
output(2, 137) <= input(10);
output(2, 138) <= input(11);
output(2, 139) <= input(12);
output(2, 140) <= input(13);
output(2, 141) <= input(14);
output(2, 142) <= input(15);
output(2, 143) <= input(38);
output(2, 144) <= input(1);
output(2, 145) <= input(2);
output(2, 146) <= input(3);
output(2, 147) <= input(4);
output(2, 148) <= input(5);
output(2, 149) <= input(6);
output(2, 150) <= input(7);
output(2, 151) <= input(8);
output(2, 152) <= input(9);
output(2, 153) <= input(10);
output(2, 154) <= input(11);
output(2, 155) <= input(12);
output(2, 156) <= input(13);
output(2, 157) <= input(14);
output(2, 158) <= input(15);
output(2, 159) <= input(38);
output(2, 160) <= input(1);
output(2, 161) <= input(2);
output(2, 162) <= input(3);
output(2, 163) <= input(4);
output(2, 164) <= input(5);
output(2, 165) <= input(6);
output(2, 166) <= input(7);
output(2, 167) <= input(8);
output(2, 168) <= input(9);
output(2, 169) <= input(10);
output(2, 170) <= input(11);
output(2, 171) <= input(12);
output(2, 172) <= input(13);
output(2, 173) <= input(14);
output(2, 174) <= input(15);
output(2, 175) <= input(38);
output(2, 176) <= input(1);
output(2, 177) <= input(2);
output(2, 178) <= input(3);
output(2, 179) <= input(4);
output(2, 180) <= input(5);
output(2, 181) <= input(6);
output(2, 182) <= input(7);
output(2, 183) <= input(8);
output(2, 184) <= input(9);
output(2, 185) <= input(10);
output(2, 186) <= input(11);
output(2, 187) <= input(12);
output(2, 188) <= input(13);
output(2, 189) <= input(14);
output(2, 190) <= input(15);
output(2, 191) <= input(38);
output(2, 192) <= input(17);
output(2, 193) <= input(18);
output(2, 194) <= input(19);
output(2, 195) <= input(20);
output(2, 196) <= input(21);
output(2, 197) <= input(22);
output(2, 198) <= input(23);
output(2, 199) <= input(24);
output(2, 200) <= input(25);
output(2, 201) <= input(26);
output(2, 202) <= input(27);
output(2, 203) <= input(28);
output(2, 204) <= input(29);
output(2, 205) <= input(30);
output(2, 206) <= input(31);
output(2, 207) <= input(39);
output(2, 208) <= input(17);
output(2, 209) <= input(18);
output(2, 210) <= input(19);
output(2, 211) <= input(20);
output(2, 212) <= input(21);
output(2, 213) <= input(22);
output(2, 214) <= input(23);
output(2, 215) <= input(24);
output(2, 216) <= input(25);
output(2, 217) <= input(26);
output(2, 218) <= input(27);
output(2, 219) <= input(28);
output(2, 220) <= input(29);
output(2, 221) <= input(30);
output(2, 222) <= input(31);
output(2, 223) <= input(39);
output(2, 224) <= input(17);
output(2, 225) <= input(18);
output(2, 226) <= input(19);
output(2, 227) <= input(20);
output(2, 228) <= input(21);
output(2, 229) <= input(22);
output(2, 230) <= input(23);
output(2, 231) <= input(24);
output(2, 232) <= input(25);
output(2, 233) <= input(26);
output(2, 234) <= input(27);
output(2, 235) <= input(28);
output(2, 236) <= input(29);
output(2, 237) <= input(30);
output(2, 238) <= input(31);
output(2, 239) <= input(39);
output(2, 240) <= input(17);
output(2, 241) <= input(18);
output(2, 242) <= input(19);
output(2, 243) <= input(20);
output(2, 244) <= input(21);
output(2, 245) <= input(22);
output(2, 246) <= input(23);
output(2, 247) <= input(24);
output(2, 248) <= input(25);
output(2, 249) <= input(26);
output(2, 250) <= input(27);
output(2, 251) <= input(28);
output(2, 252) <= input(29);
output(2, 253) <= input(30);
output(2, 254) <= input(31);
output(2, 255) <= input(39);
when "1101" =>
output(0, 0) <= input(0);
output(0, 1) <= input(1);
output(0, 2) <= input(2);
output(0, 3) <= input(3);
output(0, 4) <= input(4);
output(0, 5) <= input(5);
output(0, 6) <= input(6);
output(0, 7) <= input(7);
output(0, 8) <= input(8);
output(0, 9) <= input(9);
output(0, 10) <= input(10);
output(0, 11) <= input(11);
output(0, 12) <= input(12);
output(0, 13) <= input(13);
output(0, 14) <= input(14);
output(0, 15) <= input(15);
output(0, 16) <= input(0);
output(0, 17) <= input(1);
output(0, 18) <= input(2);
output(0, 19) <= input(3);
output(0, 20) <= input(4);
output(0, 21) <= input(5);
output(0, 22) <= input(6);
output(0, 23) <= input(7);
output(0, 24) <= input(8);
output(0, 25) <= input(9);
output(0, 26) <= input(10);
output(0, 27) <= input(11);
output(0, 28) <= input(12);
output(0, 29) <= input(13);
output(0, 30) <= input(14);
output(0, 31) <= input(15);
output(0, 32) <= input(0);
output(0, 33) <= input(1);
output(0, 34) <= input(2);
output(0, 35) <= input(3);
output(0, 36) <= input(4);
output(0, 37) <= input(5);
output(0, 38) <= input(6);
output(0, 39) <= input(7);
output(0, 40) <= input(8);
output(0, 41) <= input(9);
output(0, 42) <= input(10);
output(0, 43) <= input(11);
output(0, 44) <= input(12);
output(0, 45) <= input(13);
output(0, 46) <= input(14);
output(0, 47) <= input(15);
output(0, 48) <= input(0);
output(0, 49) <= input(1);
output(0, 50) <= input(2);
output(0, 51) <= input(3);
output(0, 52) <= input(4);
output(0, 53) <= input(5);
output(0, 54) <= input(6);
output(0, 55) <= input(7);
output(0, 56) <= input(8);
output(0, 57) <= input(9);
output(0, 58) <= input(10);
output(0, 59) <= input(11);
output(0, 60) <= input(12);
output(0, 61) <= input(13);
output(0, 62) <= input(14);
output(0, 63) <= input(15);
output(0, 64) <= input(0);
output(0, 65) <= input(1);
output(0, 66) <= input(2);
output(0, 67) <= input(3);
output(0, 68) <= input(4);
output(0, 69) <= input(5);
output(0, 70) <= input(6);
output(0, 71) <= input(7);
output(0, 72) <= input(8);
output(0, 73) <= input(9);
output(0, 74) <= input(10);
output(0, 75) <= input(11);
output(0, 76) <= input(12);
output(0, 77) <= input(13);
output(0, 78) <= input(14);
output(0, 79) <= input(15);
output(0, 80) <= input(16);
output(0, 81) <= input(17);
output(0, 82) <= input(18);
output(0, 83) <= input(19);
output(0, 84) <= input(20);
output(0, 85) <= input(21);
output(0, 86) <= input(22);
output(0, 87) <= input(23);
output(0, 88) <= input(24);
output(0, 89) <= input(25);
output(0, 90) <= input(26);
output(0, 91) <= input(27);
output(0, 92) <= input(28);
output(0, 93) <= input(29);
output(0, 94) <= input(30);
output(0, 95) <= input(31);
output(0, 96) <= input(16);
output(0, 97) <= input(17);
output(0, 98) <= input(18);
output(0, 99) <= input(19);
output(0, 100) <= input(20);
output(0, 101) <= input(21);
output(0, 102) <= input(22);
output(0, 103) <= input(23);
output(0, 104) <= input(24);
output(0, 105) <= input(25);
output(0, 106) <= input(26);
output(0, 107) <= input(27);
output(0, 108) <= input(28);
output(0, 109) <= input(29);
output(0, 110) <= input(30);
output(0, 111) <= input(31);
output(0, 112) <= input(16);
output(0, 113) <= input(17);
output(0, 114) <= input(18);
output(0, 115) <= input(19);
output(0, 116) <= input(20);
output(0, 117) <= input(21);
output(0, 118) <= input(22);
output(0, 119) <= input(23);
output(0, 120) <= input(24);
output(0, 121) <= input(25);
output(0, 122) <= input(26);
output(0, 123) <= input(27);
output(0, 124) <= input(28);
output(0, 125) <= input(29);
output(0, 126) <= input(30);
output(0, 127) <= input(31);
output(0, 128) <= input(16);
output(0, 129) <= input(17);
output(0, 130) <= input(18);
output(0, 131) <= input(19);
output(0, 132) <= input(20);
output(0, 133) <= input(21);
output(0, 134) <= input(22);
output(0, 135) <= input(23);
output(0, 136) <= input(24);
output(0, 137) <= input(25);
output(0, 138) <= input(26);
output(0, 139) <= input(27);
output(0, 140) <= input(28);
output(0, 141) <= input(29);
output(0, 142) <= input(30);
output(0, 143) <= input(31);
output(0, 144) <= input(16);
output(0, 145) <= input(17);
output(0, 146) <= input(18);
output(0, 147) <= input(19);
output(0, 148) <= input(20);
output(0, 149) <= input(21);
output(0, 150) <= input(22);
output(0, 151) <= input(23);
output(0, 152) <= input(24);
output(0, 153) <= input(25);
output(0, 154) <= input(26);
output(0, 155) <= input(27);
output(0, 156) <= input(28);
output(0, 157) <= input(29);
output(0, 158) <= input(30);
output(0, 159) <= input(31);
output(0, 160) <= input(32);
output(0, 161) <= input(0);
output(0, 162) <= input(1);
output(0, 163) <= input(2);
output(0, 164) <= input(3);
output(0, 165) <= input(4);
output(0, 166) <= input(5);
output(0, 167) <= input(6);
output(0, 168) <= input(7);
output(0, 169) <= input(8);
output(0, 170) <= input(9);
output(0, 171) <= input(10);
output(0, 172) <= input(11);
output(0, 173) <= input(12);
output(0, 174) <= input(13);
output(0, 175) <= input(14);
output(0, 176) <= input(32);
output(0, 177) <= input(0);
output(0, 178) <= input(1);
output(0, 179) <= input(2);
output(0, 180) <= input(3);
output(0, 181) <= input(4);
output(0, 182) <= input(5);
output(0, 183) <= input(6);
output(0, 184) <= input(7);
output(0, 185) <= input(8);
output(0, 186) <= input(9);
output(0, 187) <= input(10);
output(0, 188) <= input(11);
output(0, 189) <= input(12);
output(0, 190) <= input(13);
output(0, 191) <= input(14);
output(0, 192) <= input(32);
output(0, 193) <= input(0);
output(0, 194) <= input(1);
output(0, 195) <= input(2);
output(0, 196) <= input(3);
output(0, 197) <= input(4);
output(0, 198) <= input(5);
output(0, 199) <= input(6);
output(0, 200) <= input(7);
output(0, 201) <= input(8);
output(0, 202) <= input(9);
output(0, 203) <= input(10);
output(0, 204) <= input(11);
output(0, 205) <= input(12);
output(0, 206) <= input(13);
output(0, 207) <= input(14);
output(0, 208) <= input(32);
output(0, 209) <= input(0);
output(0, 210) <= input(1);
output(0, 211) <= input(2);
output(0, 212) <= input(3);
output(0, 213) <= input(4);
output(0, 214) <= input(5);
output(0, 215) <= input(6);
output(0, 216) <= input(7);
output(0, 217) <= input(8);
output(0, 218) <= input(9);
output(0, 219) <= input(10);
output(0, 220) <= input(11);
output(0, 221) <= input(12);
output(0, 222) <= input(13);
output(0, 223) <= input(14);
output(0, 224) <= input(32);
output(0, 225) <= input(0);
output(0, 226) <= input(1);
output(0, 227) <= input(2);
output(0, 228) <= input(3);
output(0, 229) <= input(4);
output(0, 230) <= input(5);
output(0, 231) <= input(6);
output(0, 232) <= input(7);
output(0, 233) <= input(8);
output(0, 234) <= input(9);
output(0, 235) <= input(10);
output(0, 236) <= input(11);
output(0, 237) <= input(12);
output(0, 238) <= input(13);
output(0, 239) <= input(14);
output(0, 240) <= input(32);
output(0, 241) <= input(0);
output(0, 242) <= input(1);
output(0, 243) <= input(2);
output(0, 244) <= input(3);
output(0, 245) <= input(4);
output(0, 246) <= input(5);
output(0, 247) <= input(6);
output(0, 248) <= input(7);
output(0, 249) <= input(8);
output(0, 250) <= input(9);
output(0, 251) <= input(10);
output(0, 252) <= input(11);
output(0, 253) <= input(12);
output(0, 254) <= input(13);
output(0, 255) <= input(14);
output(1, 0) <= input(17);
output(1, 1) <= input(18);
output(1, 2) <= input(19);
output(1, 3) <= input(20);
output(1, 4) <= input(21);
output(1, 5) <= input(22);
output(1, 6) <= input(23);
output(1, 7) <= input(24);
output(1, 8) <= input(25);
output(1, 9) <= input(26);
output(1, 10) <= input(27);
output(1, 11) <= input(28);
output(1, 12) <= input(29);
output(1, 13) <= input(30);
output(1, 14) <= input(31);
output(1, 15) <= input(33);
output(1, 16) <= input(17);
output(1, 17) <= input(18);
output(1, 18) <= input(19);
output(1, 19) <= input(20);
output(1, 20) <= input(21);
output(1, 21) <= input(22);
output(1, 22) <= input(23);
output(1, 23) <= input(24);
output(1, 24) <= input(25);
output(1, 25) <= input(26);
output(1, 26) <= input(27);
output(1, 27) <= input(28);
output(1, 28) <= input(29);
output(1, 29) <= input(30);
output(1, 30) <= input(31);
output(1, 31) <= input(33);
output(1, 32) <= input(17);
output(1, 33) <= input(18);
output(1, 34) <= input(19);
output(1, 35) <= input(20);
output(1, 36) <= input(21);
output(1, 37) <= input(22);
output(1, 38) <= input(23);
output(1, 39) <= input(24);
output(1, 40) <= input(25);
output(1, 41) <= input(26);
output(1, 42) <= input(27);
output(1, 43) <= input(28);
output(1, 44) <= input(29);
output(1, 45) <= input(30);
output(1, 46) <= input(31);
output(1, 47) <= input(33);
output(1, 48) <= input(17);
output(1, 49) <= input(18);
output(1, 50) <= input(19);
output(1, 51) <= input(20);
output(1, 52) <= input(21);
output(1, 53) <= input(22);
output(1, 54) <= input(23);
output(1, 55) <= input(24);
output(1, 56) <= input(25);
output(1, 57) <= input(26);
output(1, 58) <= input(27);
output(1, 59) <= input(28);
output(1, 60) <= input(29);
output(1, 61) <= input(30);
output(1, 62) <= input(31);
output(1, 63) <= input(33);
output(1, 64) <= input(17);
output(1, 65) <= input(18);
output(1, 66) <= input(19);
output(1, 67) <= input(20);
output(1, 68) <= input(21);
output(1, 69) <= input(22);
output(1, 70) <= input(23);
output(1, 71) <= input(24);
output(1, 72) <= input(25);
output(1, 73) <= input(26);
output(1, 74) <= input(27);
output(1, 75) <= input(28);
output(1, 76) <= input(29);
output(1, 77) <= input(30);
output(1, 78) <= input(31);
output(1, 79) <= input(33);
output(1, 80) <= input(17);
output(1, 81) <= input(18);
output(1, 82) <= input(19);
output(1, 83) <= input(20);
output(1, 84) <= input(21);
output(1, 85) <= input(22);
output(1, 86) <= input(23);
output(1, 87) <= input(24);
output(1, 88) <= input(25);
output(1, 89) <= input(26);
output(1, 90) <= input(27);
output(1, 91) <= input(28);
output(1, 92) <= input(29);
output(1, 93) <= input(30);
output(1, 94) <= input(31);
output(1, 95) <= input(33);
output(1, 96) <= input(17);
output(1, 97) <= input(18);
output(1, 98) <= input(19);
output(1, 99) <= input(20);
output(1, 100) <= input(21);
output(1, 101) <= input(22);
output(1, 102) <= input(23);
output(1, 103) <= input(24);
output(1, 104) <= input(25);
output(1, 105) <= input(26);
output(1, 106) <= input(27);
output(1, 107) <= input(28);
output(1, 108) <= input(29);
output(1, 109) <= input(30);
output(1, 110) <= input(31);
output(1, 111) <= input(33);
output(1, 112) <= input(17);
output(1, 113) <= input(18);
output(1, 114) <= input(19);
output(1, 115) <= input(20);
output(1, 116) <= input(21);
output(1, 117) <= input(22);
output(1, 118) <= input(23);
output(1, 119) <= input(24);
output(1, 120) <= input(25);
output(1, 121) <= input(26);
output(1, 122) <= input(27);
output(1, 123) <= input(28);
output(1, 124) <= input(29);
output(1, 125) <= input(30);
output(1, 126) <= input(31);
output(1, 127) <= input(33);
output(1, 128) <= input(0);
output(1, 129) <= input(1);
output(1, 130) <= input(2);
output(1, 131) <= input(3);
output(1, 132) <= input(4);
output(1, 133) <= input(5);
output(1, 134) <= input(6);
output(1, 135) <= input(7);
output(1, 136) <= input(8);
output(1, 137) <= input(9);
output(1, 138) <= input(10);
output(1, 139) <= input(11);
output(1, 140) <= input(12);
output(1, 141) <= input(13);
output(1, 142) <= input(14);
output(1, 143) <= input(15);
output(1, 144) <= input(0);
output(1, 145) <= input(1);
output(1, 146) <= input(2);
output(1, 147) <= input(3);
output(1, 148) <= input(4);
output(1, 149) <= input(5);
output(1, 150) <= input(6);
output(1, 151) <= input(7);
output(1, 152) <= input(8);
output(1, 153) <= input(9);
output(1, 154) <= input(10);
output(1, 155) <= input(11);
output(1, 156) <= input(12);
output(1, 157) <= input(13);
output(1, 158) <= input(14);
output(1, 159) <= input(15);
output(1, 160) <= input(0);
output(1, 161) <= input(1);
output(1, 162) <= input(2);
output(1, 163) <= input(3);
output(1, 164) <= input(4);
output(1, 165) <= input(5);
output(1, 166) <= input(6);
output(1, 167) <= input(7);
output(1, 168) <= input(8);
output(1, 169) <= input(9);
output(1, 170) <= input(10);
output(1, 171) <= input(11);
output(1, 172) <= input(12);
output(1, 173) <= input(13);
output(1, 174) <= input(14);
output(1, 175) <= input(15);
output(1, 176) <= input(0);
output(1, 177) <= input(1);
output(1, 178) <= input(2);
output(1, 179) <= input(3);
output(1, 180) <= input(4);
output(1, 181) <= input(5);
output(1, 182) <= input(6);
output(1, 183) <= input(7);
output(1, 184) <= input(8);
output(1, 185) <= input(9);
output(1, 186) <= input(10);
output(1, 187) <= input(11);
output(1, 188) <= input(12);
output(1, 189) <= input(13);
output(1, 190) <= input(14);
output(1, 191) <= input(15);
output(1, 192) <= input(0);
output(1, 193) <= input(1);
output(1, 194) <= input(2);
output(1, 195) <= input(3);
output(1, 196) <= input(4);
output(1, 197) <= input(5);
output(1, 198) <= input(6);
output(1, 199) <= input(7);
output(1, 200) <= input(8);
output(1, 201) <= input(9);
output(1, 202) <= input(10);
output(1, 203) <= input(11);
output(1, 204) <= input(12);
output(1, 205) <= input(13);
output(1, 206) <= input(14);
output(1, 207) <= input(15);
output(1, 208) <= input(0);
output(1, 209) <= input(1);
output(1, 210) <= input(2);
output(1, 211) <= input(3);
output(1, 212) <= input(4);
output(1, 213) <= input(5);
output(1, 214) <= input(6);
output(1, 215) <= input(7);
output(1, 216) <= input(8);
output(1, 217) <= input(9);
output(1, 218) <= input(10);
output(1, 219) <= input(11);
output(1, 220) <= input(12);
output(1, 221) <= input(13);
output(1, 222) <= input(14);
output(1, 223) <= input(15);
output(1, 224) <= input(0);
output(1, 225) <= input(1);
output(1, 226) <= input(2);
output(1, 227) <= input(3);
output(1, 228) <= input(4);
output(1, 229) <= input(5);
output(1, 230) <= input(6);
output(1, 231) <= input(7);
output(1, 232) <= input(8);
output(1, 233) <= input(9);
output(1, 234) <= input(10);
output(1, 235) <= input(11);
output(1, 236) <= input(12);
output(1, 237) <= input(13);
output(1, 238) <= input(14);
output(1, 239) <= input(15);
output(1, 240) <= input(0);
output(1, 241) <= input(1);
output(1, 242) <= input(2);
output(1, 243) <= input(3);
output(1, 244) <= input(4);
output(1, 245) <= input(5);
output(1, 246) <= input(6);
output(1, 247) <= input(7);
output(1, 248) <= input(8);
output(1, 249) <= input(9);
output(1, 250) <= input(10);
output(1, 251) <= input(11);
output(1, 252) <= input(12);
output(1, 253) <= input(13);
output(1, 254) <= input(14);
output(1, 255) <= input(15);
output(2, 0) <= input(1);
output(2, 1) <= input(2);
output(2, 2) <= input(3);
output(2, 3) <= input(4);
output(2, 4) <= input(5);
output(2, 5) <= input(6);
output(2, 6) <= input(7);
output(2, 7) <= input(8);
output(2, 8) <= input(9);
output(2, 9) <= input(10);
output(2, 10) <= input(11);
output(2, 11) <= input(12);
output(2, 12) <= input(13);
output(2, 13) <= input(14);
output(2, 14) <= input(15);
output(2, 15) <= input(34);
output(2, 16) <= input(1);
output(2, 17) <= input(2);
output(2, 18) <= input(3);
output(2, 19) <= input(4);
output(2, 20) <= input(5);
output(2, 21) <= input(6);
output(2, 22) <= input(7);
output(2, 23) <= input(8);
output(2, 24) <= input(9);
output(2, 25) <= input(10);
output(2, 26) <= input(11);
output(2, 27) <= input(12);
output(2, 28) <= input(13);
output(2, 29) <= input(14);
output(2, 30) <= input(15);
output(2, 31) <= input(34);
output(2, 32) <= input(1);
output(2, 33) <= input(2);
output(2, 34) <= input(3);
output(2, 35) <= input(4);
output(2, 36) <= input(5);
output(2, 37) <= input(6);
output(2, 38) <= input(7);
output(2, 39) <= input(8);
output(2, 40) <= input(9);
output(2, 41) <= input(10);
output(2, 42) <= input(11);
output(2, 43) <= input(12);
output(2, 44) <= input(13);
output(2, 45) <= input(14);
output(2, 46) <= input(15);
output(2, 47) <= input(34);
output(2, 48) <= input(1);
output(2, 49) <= input(2);
output(2, 50) <= input(3);
output(2, 51) <= input(4);
output(2, 52) <= input(5);
output(2, 53) <= input(6);
output(2, 54) <= input(7);
output(2, 55) <= input(8);
output(2, 56) <= input(9);
output(2, 57) <= input(10);
output(2, 58) <= input(11);
output(2, 59) <= input(12);
output(2, 60) <= input(13);
output(2, 61) <= input(14);
output(2, 62) <= input(15);
output(2, 63) <= input(34);
output(2, 64) <= input(1);
output(2, 65) <= input(2);
output(2, 66) <= input(3);
output(2, 67) <= input(4);
output(2, 68) <= input(5);
output(2, 69) <= input(6);
output(2, 70) <= input(7);
output(2, 71) <= input(8);
output(2, 72) <= input(9);
output(2, 73) <= input(10);
output(2, 74) <= input(11);
output(2, 75) <= input(12);
output(2, 76) <= input(13);
output(2, 77) <= input(14);
output(2, 78) <= input(15);
output(2, 79) <= input(34);
output(2, 80) <= input(1);
output(2, 81) <= input(2);
output(2, 82) <= input(3);
output(2, 83) <= input(4);
output(2, 84) <= input(5);
output(2, 85) <= input(6);
output(2, 86) <= input(7);
output(2, 87) <= input(8);
output(2, 88) <= input(9);
output(2, 89) <= input(10);
output(2, 90) <= input(11);
output(2, 91) <= input(12);
output(2, 92) <= input(13);
output(2, 93) <= input(14);
output(2, 94) <= input(15);
output(2, 95) <= input(34);
output(2, 96) <= input(1);
output(2, 97) <= input(2);
output(2, 98) <= input(3);
output(2, 99) <= input(4);
output(2, 100) <= input(5);
output(2, 101) <= input(6);
output(2, 102) <= input(7);
output(2, 103) <= input(8);
output(2, 104) <= input(9);
output(2, 105) <= input(10);
output(2, 106) <= input(11);
output(2, 107) <= input(12);
output(2, 108) <= input(13);
output(2, 109) <= input(14);
output(2, 110) <= input(15);
output(2, 111) <= input(34);
output(2, 112) <= input(1);
output(2, 113) <= input(2);
output(2, 114) <= input(3);
output(2, 115) <= input(4);
output(2, 116) <= input(5);
output(2, 117) <= input(6);
output(2, 118) <= input(7);
output(2, 119) <= input(8);
output(2, 120) <= input(9);
output(2, 121) <= input(10);
output(2, 122) <= input(11);
output(2, 123) <= input(12);
output(2, 124) <= input(13);
output(2, 125) <= input(14);
output(2, 126) <= input(15);
output(2, 127) <= input(34);
output(2, 128) <= input(1);
output(2, 129) <= input(2);
output(2, 130) <= input(3);
output(2, 131) <= input(4);
output(2, 132) <= input(5);
output(2, 133) <= input(6);
output(2, 134) <= input(7);
output(2, 135) <= input(8);
output(2, 136) <= input(9);
output(2, 137) <= input(10);
output(2, 138) <= input(11);
output(2, 139) <= input(12);
output(2, 140) <= input(13);
output(2, 141) <= input(14);
output(2, 142) <= input(15);
output(2, 143) <= input(34);
output(2, 144) <= input(1);
output(2, 145) <= input(2);
output(2, 146) <= input(3);
output(2, 147) <= input(4);
output(2, 148) <= input(5);
output(2, 149) <= input(6);
output(2, 150) <= input(7);
output(2, 151) <= input(8);
output(2, 152) <= input(9);
output(2, 153) <= input(10);
output(2, 154) <= input(11);
output(2, 155) <= input(12);
output(2, 156) <= input(13);
output(2, 157) <= input(14);
output(2, 158) <= input(15);
output(2, 159) <= input(34);
output(2, 160) <= input(1);
output(2, 161) <= input(2);
output(2, 162) <= input(3);
output(2, 163) <= input(4);
output(2, 164) <= input(5);
output(2, 165) <= input(6);
output(2, 166) <= input(7);
output(2, 167) <= input(8);
output(2, 168) <= input(9);
output(2, 169) <= input(10);
output(2, 170) <= input(11);
output(2, 171) <= input(12);
output(2, 172) <= input(13);
output(2, 173) <= input(14);
output(2, 174) <= input(15);
output(2, 175) <= input(34);
output(2, 176) <= input(1);
output(2, 177) <= input(2);
output(2, 178) <= input(3);
output(2, 179) <= input(4);
output(2, 180) <= input(5);
output(2, 181) <= input(6);
output(2, 182) <= input(7);
output(2, 183) <= input(8);
output(2, 184) <= input(9);
output(2, 185) <= input(10);
output(2, 186) <= input(11);
output(2, 187) <= input(12);
output(2, 188) <= input(13);
output(2, 189) <= input(14);
output(2, 190) <= input(15);
output(2, 191) <= input(34);
output(2, 192) <= input(1);
output(2, 193) <= input(2);
output(2, 194) <= input(3);
output(2, 195) <= input(4);
output(2, 196) <= input(5);
output(2, 197) <= input(6);
output(2, 198) <= input(7);
output(2, 199) <= input(8);
output(2, 200) <= input(9);
output(2, 201) <= input(10);
output(2, 202) <= input(11);
output(2, 203) <= input(12);
output(2, 204) <= input(13);
output(2, 205) <= input(14);
output(2, 206) <= input(15);
output(2, 207) <= input(34);
output(2, 208) <= input(1);
output(2, 209) <= input(2);
output(2, 210) <= input(3);
output(2, 211) <= input(4);
output(2, 212) <= input(5);
output(2, 213) <= input(6);
output(2, 214) <= input(7);
output(2, 215) <= input(8);
output(2, 216) <= input(9);
output(2, 217) <= input(10);
output(2, 218) <= input(11);
output(2, 219) <= input(12);
output(2, 220) <= input(13);
output(2, 221) <= input(14);
output(2, 222) <= input(15);
output(2, 223) <= input(34);
output(2, 224) <= input(1);
output(2, 225) <= input(2);
output(2, 226) <= input(3);
output(2, 227) <= input(4);
output(2, 228) <= input(5);
output(2, 229) <= input(6);
output(2, 230) <= input(7);
output(2, 231) <= input(8);
output(2, 232) <= input(9);
output(2, 233) <= input(10);
output(2, 234) <= input(11);
output(2, 235) <= input(12);
output(2, 236) <= input(13);
output(2, 237) <= input(14);
output(2, 238) <= input(15);
output(2, 239) <= input(34);
output(2, 240) <= input(1);
output(2, 241) <= input(2);
output(2, 242) <= input(3);
output(2, 243) <= input(4);
output(2, 244) <= input(5);
output(2, 245) <= input(6);
output(2, 246) <= input(7);
output(2, 247) <= input(8);
output(2, 248) <= input(9);
output(2, 249) <= input(10);
output(2, 250) <= input(11);
output(2, 251) <= input(12);
output(2, 252) <= input(13);
output(2, 253) <= input(14);
output(2, 254) <= input(15);
output(2, 255) <= input(34);
output(3, 0) <= input(2);
output(3, 1) <= input(3);
output(3, 2) <= input(4);
output(3, 3) <= input(5);
output(3, 4) <= input(6);
output(3, 5) <= input(7);
output(3, 6) <= input(8);
output(3, 7) <= input(9);
output(3, 8) <= input(10);
output(3, 9) <= input(11);
output(3, 10) <= input(12);
output(3, 11) <= input(13);
output(3, 12) <= input(14);
output(3, 13) <= input(15);
output(3, 14) <= input(34);
output(3, 15) <= input(35);
output(3, 16) <= input(2);
output(3, 17) <= input(3);
output(3, 18) <= input(4);
output(3, 19) <= input(5);
output(3, 20) <= input(6);
output(3, 21) <= input(7);
output(3, 22) <= input(8);
output(3, 23) <= input(9);
output(3, 24) <= input(10);
output(3, 25) <= input(11);
output(3, 26) <= input(12);
output(3, 27) <= input(13);
output(3, 28) <= input(14);
output(3, 29) <= input(15);
output(3, 30) <= input(34);
output(3, 31) <= input(35);
output(3, 32) <= input(2);
output(3, 33) <= input(3);
output(3, 34) <= input(4);
output(3, 35) <= input(5);
output(3, 36) <= input(6);
output(3, 37) <= input(7);
output(3, 38) <= input(8);
output(3, 39) <= input(9);
output(3, 40) <= input(10);
output(3, 41) <= input(11);
output(3, 42) <= input(12);
output(3, 43) <= input(13);
output(3, 44) <= input(14);
output(3, 45) <= input(15);
output(3, 46) <= input(34);
output(3, 47) <= input(35);
output(3, 48) <= input(2);
output(3, 49) <= input(3);
output(3, 50) <= input(4);
output(3, 51) <= input(5);
output(3, 52) <= input(6);
output(3, 53) <= input(7);
output(3, 54) <= input(8);
output(3, 55) <= input(9);
output(3, 56) <= input(10);
output(3, 57) <= input(11);
output(3, 58) <= input(12);
output(3, 59) <= input(13);
output(3, 60) <= input(14);
output(3, 61) <= input(15);
output(3, 62) <= input(34);
output(3, 63) <= input(35);
output(3, 64) <= input(2);
output(3, 65) <= input(3);
output(3, 66) <= input(4);
output(3, 67) <= input(5);
output(3, 68) <= input(6);
output(3, 69) <= input(7);
output(3, 70) <= input(8);
output(3, 71) <= input(9);
output(3, 72) <= input(10);
output(3, 73) <= input(11);
output(3, 74) <= input(12);
output(3, 75) <= input(13);
output(3, 76) <= input(14);
output(3, 77) <= input(15);
output(3, 78) <= input(34);
output(3, 79) <= input(35);
output(3, 80) <= input(2);
output(3, 81) <= input(3);
output(3, 82) <= input(4);
output(3, 83) <= input(5);
output(3, 84) <= input(6);
output(3, 85) <= input(7);
output(3, 86) <= input(8);
output(3, 87) <= input(9);
output(3, 88) <= input(10);
output(3, 89) <= input(11);
output(3, 90) <= input(12);
output(3, 91) <= input(13);
output(3, 92) <= input(14);
output(3, 93) <= input(15);
output(3, 94) <= input(34);
output(3, 95) <= input(35);
output(3, 96) <= input(2);
output(3, 97) <= input(3);
output(3, 98) <= input(4);
output(3, 99) <= input(5);
output(3, 100) <= input(6);
output(3, 101) <= input(7);
output(3, 102) <= input(8);
output(3, 103) <= input(9);
output(3, 104) <= input(10);
output(3, 105) <= input(11);
output(3, 106) <= input(12);
output(3, 107) <= input(13);
output(3, 108) <= input(14);
output(3, 109) <= input(15);
output(3, 110) <= input(34);
output(3, 111) <= input(35);
output(3, 112) <= input(2);
output(3, 113) <= input(3);
output(3, 114) <= input(4);
output(3, 115) <= input(5);
output(3, 116) <= input(6);
output(3, 117) <= input(7);
output(3, 118) <= input(8);
output(3, 119) <= input(9);
output(3, 120) <= input(10);
output(3, 121) <= input(11);
output(3, 122) <= input(12);
output(3, 123) <= input(13);
output(3, 124) <= input(14);
output(3, 125) <= input(15);
output(3, 126) <= input(34);
output(3, 127) <= input(35);
output(3, 128) <= input(2);
output(3, 129) <= input(3);
output(3, 130) <= input(4);
output(3, 131) <= input(5);
output(3, 132) <= input(6);
output(3, 133) <= input(7);
output(3, 134) <= input(8);
output(3, 135) <= input(9);
output(3, 136) <= input(10);
output(3, 137) <= input(11);
output(3, 138) <= input(12);
output(3, 139) <= input(13);
output(3, 140) <= input(14);
output(3, 141) <= input(15);
output(3, 142) <= input(34);
output(3, 143) <= input(35);
output(3, 144) <= input(2);
output(3, 145) <= input(3);
output(3, 146) <= input(4);
output(3, 147) <= input(5);
output(3, 148) <= input(6);
output(3, 149) <= input(7);
output(3, 150) <= input(8);
output(3, 151) <= input(9);
output(3, 152) <= input(10);
output(3, 153) <= input(11);
output(3, 154) <= input(12);
output(3, 155) <= input(13);
output(3, 156) <= input(14);
output(3, 157) <= input(15);
output(3, 158) <= input(34);
output(3, 159) <= input(35);
output(3, 160) <= input(2);
output(3, 161) <= input(3);
output(3, 162) <= input(4);
output(3, 163) <= input(5);
output(3, 164) <= input(6);
output(3, 165) <= input(7);
output(3, 166) <= input(8);
output(3, 167) <= input(9);
output(3, 168) <= input(10);
output(3, 169) <= input(11);
output(3, 170) <= input(12);
output(3, 171) <= input(13);
output(3, 172) <= input(14);
output(3, 173) <= input(15);
output(3, 174) <= input(34);
output(3, 175) <= input(35);
output(3, 176) <= input(2);
output(3, 177) <= input(3);
output(3, 178) <= input(4);
output(3, 179) <= input(5);
output(3, 180) <= input(6);
output(3, 181) <= input(7);
output(3, 182) <= input(8);
output(3, 183) <= input(9);
output(3, 184) <= input(10);
output(3, 185) <= input(11);
output(3, 186) <= input(12);
output(3, 187) <= input(13);
output(3, 188) <= input(14);
output(3, 189) <= input(15);
output(3, 190) <= input(34);
output(3, 191) <= input(35);
output(3, 192) <= input(2);
output(3, 193) <= input(3);
output(3, 194) <= input(4);
output(3, 195) <= input(5);
output(3, 196) <= input(6);
output(3, 197) <= input(7);
output(3, 198) <= input(8);
output(3, 199) <= input(9);
output(3, 200) <= input(10);
output(3, 201) <= input(11);
output(3, 202) <= input(12);
output(3, 203) <= input(13);
output(3, 204) <= input(14);
output(3, 205) <= input(15);
output(3, 206) <= input(34);
output(3, 207) <= input(35);
output(3, 208) <= input(2);
output(3, 209) <= input(3);
output(3, 210) <= input(4);
output(3, 211) <= input(5);
output(3, 212) <= input(6);
output(3, 213) <= input(7);
output(3, 214) <= input(8);
output(3, 215) <= input(9);
output(3, 216) <= input(10);
output(3, 217) <= input(11);
output(3, 218) <= input(12);
output(3, 219) <= input(13);
output(3, 220) <= input(14);
output(3, 221) <= input(15);
output(3, 222) <= input(34);
output(3, 223) <= input(35);
output(3, 224) <= input(2);
output(3, 225) <= input(3);
output(3, 226) <= input(4);
output(3, 227) <= input(5);
output(3, 228) <= input(6);
output(3, 229) <= input(7);
output(3, 230) <= input(8);
output(3, 231) <= input(9);
output(3, 232) <= input(10);
output(3, 233) <= input(11);
output(3, 234) <= input(12);
output(3, 235) <= input(13);
output(3, 236) <= input(14);
output(3, 237) <= input(15);
output(3, 238) <= input(34);
output(3, 239) <= input(35);
output(3, 240) <= input(2);
output(3, 241) <= input(3);
output(3, 242) <= input(4);
output(3, 243) <= input(5);
output(3, 244) <= input(6);
output(3, 245) <= input(7);
output(3, 246) <= input(8);
output(3, 247) <= input(9);
output(3, 248) <= input(10);
output(3, 249) <= input(11);
output(3, 250) <= input(12);
output(3, 251) <= input(13);
output(3, 252) <= input(14);
output(3, 253) <= input(15);
output(3, 254) <= input(34);
output(3, 255) <= input(35);
output(4, 0) <= input(19);
output(4, 1) <= input(20);
output(4, 2) <= input(21);
output(4, 3) <= input(22);
output(4, 4) <= input(23);
output(4, 5) <= input(24);
output(4, 6) <= input(25);
output(4, 7) <= input(26);
output(4, 8) <= input(27);
output(4, 9) <= input(28);
output(4, 10) <= input(29);
output(4, 11) <= input(30);
output(4, 12) <= input(31);
output(4, 13) <= input(33);
output(4, 14) <= input(36);
output(4, 15) <= input(37);
output(4, 16) <= input(19);
output(4, 17) <= input(20);
output(4, 18) <= input(21);
output(4, 19) <= input(22);
output(4, 20) <= input(23);
output(4, 21) <= input(24);
output(4, 22) <= input(25);
output(4, 23) <= input(26);
output(4, 24) <= input(27);
output(4, 25) <= input(28);
output(4, 26) <= input(29);
output(4, 27) <= input(30);
output(4, 28) <= input(31);
output(4, 29) <= input(33);
output(4, 30) <= input(36);
output(4, 31) <= input(37);
output(4, 32) <= input(19);
output(4, 33) <= input(20);
output(4, 34) <= input(21);
output(4, 35) <= input(22);
output(4, 36) <= input(23);
output(4, 37) <= input(24);
output(4, 38) <= input(25);
output(4, 39) <= input(26);
output(4, 40) <= input(27);
output(4, 41) <= input(28);
output(4, 42) <= input(29);
output(4, 43) <= input(30);
output(4, 44) <= input(31);
output(4, 45) <= input(33);
output(4, 46) <= input(36);
output(4, 47) <= input(37);
output(4, 48) <= input(19);
output(4, 49) <= input(20);
output(4, 50) <= input(21);
output(4, 51) <= input(22);
output(4, 52) <= input(23);
output(4, 53) <= input(24);
output(4, 54) <= input(25);
output(4, 55) <= input(26);
output(4, 56) <= input(27);
output(4, 57) <= input(28);
output(4, 58) <= input(29);
output(4, 59) <= input(30);
output(4, 60) <= input(31);
output(4, 61) <= input(33);
output(4, 62) <= input(36);
output(4, 63) <= input(37);
output(4, 64) <= input(19);
output(4, 65) <= input(20);
output(4, 66) <= input(21);
output(4, 67) <= input(22);
output(4, 68) <= input(23);
output(4, 69) <= input(24);
output(4, 70) <= input(25);
output(4, 71) <= input(26);
output(4, 72) <= input(27);
output(4, 73) <= input(28);
output(4, 74) <= input(29);
output(4, 75) <= input(30);
output(4, 76) <= input(31);
output(4, 77) <= input(33);
output(4, 78) <= input(36);
output(4, 79) <= input(37);
output(4, 80) <= input(19);
output(4, 81) <= input(20);
output(4, 82) <= input(21);
output(4, 83) <= input(22);
output(4, 84) <= input(23);
output(4, 85) <= input(24);
output(4, 86) <= input(25);
output(4, 87) <= input(26);
output(4, 88) <= input(27);
output(4, 89) <= input(28);
output(4, 90) <= input(29);
output(4, 91) <= input(30);
output(4, 92) <= input(31);
output(4, 93) <= input(33);
output(4, 94) <= input(36);
output(4, 95) <= input(37);
output(4, 96) <= input(19);
output(4, 97) <= input(20);
output(4, 98) <= input(21);
output(4, 99) <= input(22);
output(4, 100) <= input(23);
output(4, 101) <= input(24);
output(4, 102) <= input(25);
output(4, 103) <= input(26);
output(4, 104) <= input(27);
output(4, 105) <= input(28);
output(4, 106) <= input(29);
output(4, 107) <= input(30);
output(4, 108) <= input(31);
output(4, 109) <= input(33);
output(4, 110) <= input(36);
output(4, 111) <= input(37);
output(4, 112) <= input(19);
output(4, 113) <= input(20);
output(4, 114) <= input(21);
output(4, 115) <= input(22);
output(4, 116) <= input(23);
output(4, 117) <= input(24);
output(4, 118) <= input(25);
output(4, 119) <= input(26);
output(4, 120) <= input(27);
output(4, 121) <= input(28);
output(4, 122) <= input(29);
output(4, 123) <= input(30);
output(4, 124) <= input(31);
output(4, 125) <= input(33);
output(4, 126) <= input(36);
output(4, 127) <= input(37);
output(4, 128) <= input(19);
output(4, 129) <= input(20);
output(4, 130) <= input(21);
output(4, 131) <= input(22);
output(4, 132) <= input(23);
output(4, 133) <= input(24);
output(4, 134) <= input(25);
output(4, 135) <= input(26);
output(4, 136) <= input(27);
output(4, 137) <= input(28);
output(4, 138) <= input(29);
output(4, 139) <= input(30);
output(4, 140) <= input(31);
output(4, 141) <= input(33);
output(4, 142) <= input(36);
output(4, 143) <= input(37);
output(4, 144) <= input(19);
output(4, 145) <= input(20);
output(4, 146) <= input(21);
output(4, 147) <= input(22);
output(4, 148) <= input(23);
output(4, 149) <= input(24);
output(4, 150) <= input(25);
output(4, 151) <= input(26);
output(4, 152) <= input(27);
output(4, 153) <= input(28);
output(4, 154) <= input(29);
output(4, 155) <= input(30);
output(4, 156) <= input(31);
output(4, 157) <= input(33);
output(4, 158) <= input(36);
output(4, 159) <= input(37);
output(4, 160) <= input(19);
output(4, 161) <= input(20);
output(4, 162) <= input(21);
output(4, 163) <= input(22);
output(4, 164) <= input(23);
output(4, 165) <= input(24);
output(4, 166) <= input(25);
output(4, 167) <= input(26);
output(4, 168) <= input(27);
output(4, 169) <= input(28);
output(4, 170) <= input(29);
output(4, 171) <= input(30);
output(4, 172) <= input(31);
output(4, 173) <= input(33);
output(4, 174) <= input(36);
output(4, 175) <= input(37);
output(4, 176) <= input(19);
output(4, 177) <= input(20);
output(4, 178) <= input(21);
output(4, 179) <= input(22);
output(4, 180) <= input(23);
output(4, 181) <= input(24);
output(4, 182) <= input(25);
output(4, 183) <= input(26);
output(4, 184) <= input(27);
output(4, 185) <= input(28);
output(4, 186) <= input(29);
output(4, 187) <= input(30);
output(4, 188) <= input(31);
output(4, 189) <= input(33);
output(4, 190) <= input(36);
output(4, 191) <= input(37);
output(4, 192) <= input(19);
output(4, 193) <= input(20);
output(4, 194) <= input(21);
output(4, 195) <= input(22);
output(4, 196) <= input(23);
output(4, 197) <= input(24);
output(4, 198) <= input(25);
output(4, 199) <= input(26);
output(4, 200) <= input(27);
output(4, 201) <= input(28);
output(4, 202) <= input(29);
output(4, 203) <= input(30);
output(4, 204) <= input(31);
output(4, 205) <= input(33);
output(4, 206) <= input(36);
output(4, 207) <= input(37);
output(4, 208) <= input(19);
output(4, 209) <= input(20);
output(4, 210) <= input(21);
output(4, 211) <= input(22);
output(4, 212) <= input(23);
output(4, 213) <= input(24);
output(4, 214) <= input(25);
output(4, 215) <= input(26);
output(4, 216) <= input(27);
output(4, 217) <= input(28);
output(4, 218) <= input(29);
output(4, 219) <= input(30);
output(4, 220) <= input(31);
output(4, 221) <= input(33);
output(4, 222) <= input(36);
output(4, 223) <= input(37);
output(4, 224) <= input(19);
output(4, 225) <= input(20);
output(4, 226) <= input(21);
output(4, 227) <= input(22);
output(4, 228) <= input(23);
output(4, 229) <= input(24);
output(4, 230) <= input(25);
output(4, 231) <= input(26);
output(4, 232) <= input(27);
output(4, 233) <= input(28);
output(4, 234) <= input(29);
output(4, 235) <= input(30);
output(4, 236) <= input(31);
output(4, 237) <= input(33);
output(4, 238) <= input(36);
output(4, 239) <= input(37);
output(4, 240) <= input(3);
output(4, 241) <= input(4);
output(4, 242) <= input(5);
output(4, 243) <= input(6);
output(4, 244) <= input(7);
output(4, 245) <= input(8);
output(4, 246) <= input(9);
output(4, 247) <= input(10);
output(4, 248) <= input(11);
output(4, 249) <= input(12);
output(4, 250) <= input(13);
output(4, 251) <= input(14);
output(4, 252) <= input(15);
output(4, 253) <= input(34);
output(4, 254) <= input(35);
output(4, 255) <= input(38);
output(5, 0) <= input(3);
output(5, 1) <= input(4);
output(5, 2) <= input(5);
output(5, 3) <= input(6);
output(5, 4) <= input(7);
output(5, 5) <= input(8);
output(5, 6) <= input(9);
output(5, 7) <= input(10);
output(5, 8) <= input(11);
output(5, 9) <= input(12);
output(5, 10) <= input(13);
output(5, 11) <= input(14);
output(5, 12) <= input(15);
output(5, 13) <= input(34);
output(5, 14) <= input(35);
output(5, 15) <= input(38);
output(5, 16) <= input(3);
output(5, 17) <= input(4);
output(5, 18) <= input(5);
output(5, 19) <= input(6);
output(5, 20) <= input(7);
output(5, 21) <= input(8);
output(5, 22) <= input(9);
output(5, 23) <= input(10);
output(5, 24) <= input(11);
output(5, 25) <= input(12);
output(5, 26) <= input(13);
output(5, 27) <= input(14);
output(5, 28) <= input(15);
output(5, 29) <= input(34);
output(5, 30) <= input(35);
output(5, 31) <= input(38);
output(5, 32) <= input(3);
output(5, 33) <= input(4);
output(5, 34) <= input(5);
output(5, 35) <= input(6);
output(5, 36) <= input(7);
output(5, 37) <= input(8);
output(5, 38) <= input(9);
output(5, 39) <= input(10);
output(5, 40) <= input(11);
output(5, 41) <= input(12);
output(5, 42) <= input(13);
output(5, 43) <= input(14);
output(5, 44) <= input(15);
output(5, 45) <= input(34);
output(5, 46) <= input(35);
output(5, 47) <= input(38);
output(5, 48) <= input(3);
output(5, 49) <= input(4);
output(5, 50) <= input(5);
output(5, 51) <= input(6);
output(5, 52) <= input(7);
output(5, 53) <= input(8);
output(5, 54) <= input(9);
output(5, 55) <= input(10);
output(5, 56) <= input(11);
output(5, 57) <= input(12);
output(5, 58) <= input(13);
output(5, 59) <= input(14);
output(5, 60) <= input(15);
output(5, 61) <= input(34);
output(5, 62) <= input(35);
output(5, 63) <= input(38);
output(5, 64) <= input(3);
output(5, 65) <= input(4);
output(5, 66) <= input(5);
output(5, 67) <= input(6);
output(5, 68) <= input(7);
output(5, 69) <= input(8);
output(5, 70) <= input(9);
output(5, 71) <= input(10);
output(5, 72) <= input(11);
output(5, 73) <= input(12);
output(5, 74) <= input(13);
output(5, 75) <= input(14);
output(5, 76) <= input(15);
output(5, 77) <= input(34);
output(5, 78) <= input(35);
output(5, 79) <= input(38);
output(5, 80) <= input(3);
output(5, 81) <= input(4);
output(5, 82) <= input(5);
output(5, 83) <= input(6);
output(5, 84) <= input(7);
output(5, 85) <= input(8);
output(5, 86) <= input(9);
output(5, 87) <= input(10);
output(5, 88) <= input(11);
output(5, 89) <= input(12);
output(5, 90) <= input(13);
output(5, 91) <= input(14);
output(5, 92) <= input(15);
output(5, 93) <= input(34);
output(5, 94) <= input(35);
output(5, 95) <= input(38);
output(5, 96) <= input(3);
output(5, 97) <= input(4);
output(5, 98) <= input(5);
output(5, 99) <= input(6);
output(5, 100) <= input(7);
output(5, 101) <= input(8);
output(5, 102) <= input(9);
output(5, 103) <= input(10);
output(5, 104) <= input(11);
output(5, 105) <= input(12);
output(5, 106) <= input(13);
output(5, 107) <= input(14);
output(5, 108) <= input(15);
output(5, 109) <= input(34);
output(5, 110) <= input(35);
output(5, 111) <= input(38);
output(5, 112) <= input(20);
output(5, 113) <= input(21);
output(5, 114) <= input(22);
output(5, 115) <= input(23);
output(5, 116) <= input(24);
output(5, 117) <= input(25);
output(5, 118) <= input(26);
output(5, 119) <= input(27);
output(5, 120) <= input(28);
output(5, 121) <= input(29);
output(5, 122) <= input(30);
output(5, 123) <= input(31);
output(5, 124) <= input(33);
output(5, 125) <= input(36);
output(5, 126) <= input(37);
output(5, 127) <= input(39);
output(5, 128) <= input(20);
output(5, 129) <= input(21);
output(5, 130) <= input(22);
output(5, 131) <= input(23);
output(5, 132) <= input(24);
output(5, 133) <= input(25);
output(5, 134) <= input(26);
output(5, 135) <= input(27);
output(5, 136) <= input(28);
output(5, 137) <= input(29);
output(5, 138) <= input(30);
output(5, 139) <= input(31);
output(5, 140) <= input(33);
output(5, 141) <= input(36);
output(5, 142) <= input(37);
output(5, 143) <= input(39);
output(5, 144) <= input(20);
output(5, 145) <= input(21);
output(5, 146) <= input(22);
output(5, 147) <= input(23);
output(5, 148) <= input(24);
output(5, 149) <= input(25);
output(5, 150) <= input(26);
output(5, 151) <= input(27);
output(5, 152) <= input(28);
output(5, 153) <= input(29);
output(5, 154) <= input(30);
output(5, 155) <= input(31);
output(5, 156) <= input(33);
output(5, 157) <= input(36);
output(5, 158) <= input(37);
output(5, 159) <= input(39);
output(5, 160) <= input(20);
output(5, 161) <= input(21);
output(5, 162) <= input(22);
output(5, 163) <= input(23);
output(5, 164) <= input(24);
output(5, 165) <= input(25);
output(5, 166) <= input(26);
output(5, 167) <= input(27);
output(5, 168) <= input(28);
output(5, 169) <= input(29);
output(5, 170) <= input(30);
output(5, 171) <= input(31);
output(5, 172) <= input(33);
output(5, 173) <= input(36);
output(5, 174) <= input(37);
output(5, 175) <= input(39);
output(5, 176) <= input(20);
output(5, 177) <= input(21);
output(5, 178) <= input(22);
output(5, 179) <= input(23);
output(5, 180) <= input(24);
output(5, 181) <= input(25);
output(5, 182) <= input(26);
output(5, 183) <= input(27);
output(5, 184) <= input(28);
output(5, 185) <= input(29);
output(5, 186) <= input(30);
output(5, 187) <= input(31);
output(5, 188) <= input(33);
output(5, 189) <= input(36);
output(5, 190) <= input(37);
output(5, 191) <= input(39);
output(5, 192) <= input(20);
output(5, 193) <= input(21);
output(5, 194) <= input(22);
output(5, 195) <= input(23);
output(5, 196) <= input(24);
output(5, 197) <= input(25);
output(5, 198) <= input(26);
output(5, 199) <= input(27);
output(5, 200) <= input(28);
output(5, 201) <= input(29);
output(5, 202) <= input(30);
output(5, 203) <= input(31);
output(5, 204) <= input(33);
output(5, 205) <= input(36);
output(5, 206) <= input(37);
output(5, 207) <= input(39);
output(5, 208) <= input(20);
output(5, 209) <= input(21);
output(5, 210) <= input(22);
output(5, 211) <= input(23);
output(5, 212) <= input(24);
output(5, 213) <= input(25);
output(5, 214) <= input(26);
output(5, 215) <= input(27);
output(5, 216) <= input(28);
output(5, 217) <= input(29);
output(5, 218) <= input(30);
output(5, 219) <= input(31);
output(5, 220) <= input(33);
output(5, 221) <= input(36);
output(5, 222) <= input(37);
output(5, 223) <= input(39);
output(5, 224) <= input(20);
output(5, 225) <= input(21);
output(5, 226) <= input(22);
output(5, 227) <= input(23);
output(5, 228) <= input(24);
output(5, 229) <= input(25);
output(5, 230) <= input(26);
output(5, 231) <= input(27);
output(5, 232) <= input(28);
output(5, 233) <= input(29);
output(5, 234) <= input(30);
output(5, 235) <= input(31);
output(5, 236) <= input(33);
output(5, 237) <= input(36);
output(5, 238) <= input(37);
output(5, 239) <= input(39);
output(5, 240) <= input(4);
output(5, 241) <= input(5);
output(5, 242) <= input(6);
output(5, 243) <= input(7);
output(5, 244) <= input(8);
output(5, 245) <= input(9);
output(5, 246) <= input(10);
output(5, 247) <= input(11);
output(5, 248) <= input(12);
output(5, 249) <= input(13);
output(5, 250) <= input(14);
output(5, 251) <= input(15);
output(5, 252) <= input(34);
output(5, 253) <= input(35);
output(5, 254) <= input(38);
output(5, 255) <= input(40);
output(6, 0) <= input(20);
output(6, 1) <= input(21);
output(6, 2) <= input(22);
output(6, 3) <= input(23);
output(6, 4) <= input(24);
output(6, 5) <= input(25);
output(6, 6) <= input(26);
output(6, 7) <= input(27);
output(6, 8) <= input(28);
output(6, 9) <= input(29);
output(6, 10) <= input(30);
output(6, 11) <= input(31);
output(6, 12) <= input(33);
output(6, 13) <= input(36);
output(6, 14) <= input(37);
output(6, 15) <= input(39);
output(6, 16) <= input(20);
output(6, 17) <= input(21);
output(6, 18) <= input(22);
output(6, 19) <= input(23);
output(6, 20) <= input(24);
output(6, 21) <= input(25);
output(6, 22) <= input(26);
output(6, 23) <= input(27);
output(6, 24) <= input(28);
output(6, 25) <= input(29);
output(6, 26) <= input(30);
output(6, 27) <= input(31);
output(6, 28) <= input(33);
output(6, 29) <= input(36);
output(6, 30) <= input(37);
output(6, 31) <= input(39);
output(6, 32) <= input(20);
output(6, 33) <= input(21);
output(6, 34) <= input(22);
output(6, 35) <= input(23);
output(6, 36) <= input(24);
output(6, 37) <= input(25);
output(6, 38) <= input(26);
output(6, 39) <= input(27);
output(6, 40) <= input(28);
output(6, 41) <= input(29);
output(6, 42) <= input(30);
output(6, 43) <= input(31);
output(6, 44) <= input(33);
output(6, 45) <= input(36);
output(6, 46) <= input(37);
output(6, 47) <= input(39);
output(6, 48) <= input(20);
output(6, 49) <= input(21);
output(6, 50) <= input(22);
output(6, 51) <= input(23);
output(6, 52) <= input(24);
output(6, 53) <= input(25);
output(6, 54) <= input(26);
output(6, 55) <= input(27);
output(6, 56) <= input(28);
output(6, 57) <= input(29);
output(6, 58) <= input(30);
output(6, 59) <= input(31);
output(6, 60) <= input(33);
output(6, 61) <= input(36);
output(6, 62) <= input(37);
output(6, 63) <= input(39);
output(6, 64) <= input(20);
output(6, 65) <= input(21);
output(6, 66) <= input(22);
output(6, 67) <= input(23);
output(6, 68) <= input(24);
output(6, 69) <= input(25);
output(6, 70) <= input(26);
output(6, 71) <= input(27);
output(6, 72) <= input(28);
output(6, 73) <= input(29);
output(6, 74) <= input(30);
output(6, 75) <= input(31);
output(6, 76) <= input(33);
output(6, 77) <= input(36);
output(6, 78) <= input(37);
output(6, 79) <= input(39);
output(6, 80) <= input(4);
output(6, 81) <= input(5);
output(6, 82) <= input(6);
output(6, 83) <= input(7);
output(6, 84) <= input(8);
output(6, 85) <= input(9);
output(6, 86) <= input(10);
output(6, 87) <= input(11);
output(6, 88) <= input(12);
output(6, 89) <= input(13);
output(6, 90) <= input(14);
output(6, 91) <= input(15);
output(6, 92) <= input(34);
output(6, 93) <= input(35);
output(6, 94) <= input(38);
output(6, 95) <= input(40);
output(6, 96) <= input(4);
output(6, 97) <= input(5);
output(6, 98) <= input(6);
output(6, 99) <= input(7);
output(6, 100) <= input(8);
output(6, 101) <= input(9);
output(6, 102) <= input(10);
output(6, 103) <= input(11);
output(6, 104) <= input(12);
output(6, 105) <= input(13);
output(6, 106) <= input(14);
output(6, 107) <= input(15);
output(6, 108) <= input(34);
output(6, 109) <= input(35);
output(6, 110) <= input(38);
output(6, 111) <= input(40);
output(6, 112) <= input(4);
output(6, 113) <= input(5);
output(6, 114) <= input(6);
output(6, 115) <= input(7);
output(6, 116) <= input(8);
output(6, 117) <= input(9);
output(6, 118) <= input(10);
output(6, 119) <= input(11);
output(6, 120) <= input(12);
output(6, 121) <= input(13);
output(6, 122) <= input(14);
output(6, 123) <= input(15);
output(6, 124) <= input(34);
output(6, 125) <= input(35);
output(6, 126) <= input(38);
output(6, 127) <= input(40);
output(6, 128) <= input(4);
output(6, 129) <= input(5);
output(6, 130) <= input(6);
output(6, 131) <= input(7);
output(6, 132) <= input(8);
output(6, 133) <= input(9);
output(6, 134) <= input(10);
output(6, 135) <= input(11);
output(6, 136) <= input(12);
output(6, 137) <= input(13);
output(6, 138) <= input(14);
output(6, 139) <= input(15);
output(6, 140) <= input(34);
output(6, 141) <= input(35);
output(6, 142) <= input(38);
output(6, 143) <= input(40);
output(6, 144) <= input(4);
output(6, 145) <= input(5);
output(6, 146) <= input(6);
output(6, 147) <= input(7);
output(6, 148) <= input(8);
output(6, 149) <= input(9);
output(6, 150) <= input(10);
output(6, 151) <= input(11);
output(6, 152) <= input(12);
output(6, 153) <= input(13);
output(6, 154) <= input(14);
output(6, 155) <= input(15);
output(6, 156) <= input(34);
output(6, 157) <= input(35);
output(6, 158) <= input(38);
output(6, 159) <= input(40);
output(6, 160) <= input(21);
output(6, 161) <= input(22);
output(6, 162) <= input(23);
output(6, 163) <= input(24);
output(6, 164) <= input(25);
output(6, 165) <= input(26);
output(6, 166) <= input(27);
output(6, 167) <= input(28);
output(6, 168) <= input(29);
output(6, 169) <= input(30);
output(6, 170) <= input(31);
output(6, 171) <= input(33);
output(6, 172) <= input(36);
output(6, 173) <= input(37);
output(6, 174) <= input(39);
output(6, 175) <= input(41);
output(6, 176) <= input(21);
output(6, 177) <= input(22);
output(6, 178) <= input(23);
output(6, 179) <= input(24);
output(6, 180) <= input(25);
output(6, 181) <= input(26);
output(6, 182) <= input(27);
output(6, 183) <= input(28);
output(6, 184) <= input(29);
output(6, 185) <= input(30);
output(6, 186) <= input(31);
output(6, 187) <= input(33);
output(6, 188) <= input(36);
output(6, 189) <= input(37);
output(6, 190) <= input(39);
output(6, 191) <= input(41);
output(6, 192) <= input(21);
output(6, 193) <= input(22);
output(6, 194) <= input(23);
output(6, 195) <= input(24);
output(6, 196) <= input(25);
output(6, 197) <= input(26);
output(6, 198) <= input(27);
output(6, 199) <= input(28);
output(6, 200) <= input(29);
output(6, 201) <= input(30);
output(6, 202) <= input(31);
output(6, 203) <= input(33);
output(6, 204) <= input(36);
output(6, 205) <= input(37);
output(6, 206) <= input(39);
output(6, 207) <= input(41);
output(6, 208) <= input(21);
output(6, 209) <= input(22);
output(6, 210) <= input(23);
output(6, 211) <= input(24);
output(6, 212) <= input(25);
output(6, 213) <= input(26);
output(6, 214) <= input(27);
output(6, 215) <= input(28);
output(6, 216) <= input(29);
output(6, 217) <= input(30);
output(6, 218) <= input(31);
output(6, 219) <= input(33);
output(6, 220) <= input(36);
output(6, 221) <= input(37);
output(6, 222) <= input(39);
output(6, 223) <= input(41);
output(6, 224) <= input(21);
output(6, 225) <= input(22);
output(6, 226) <= input(23);
output(6, 227) <= input(24);
output(6, 228) <= input(25);
output(6, 229) <= input(26);
output(6, 230) <= input(27);
output(6, 231) <= input(28);
output(6, 232) <= input(29);
output(6, 233) <= input(30);
output(6, 234) <= input(31);
output(6, 235) <= input(33);
output(6, 236) <= input(36);
output(6, 237) <= input(37);
output(6, 238) <= input(39);
output(6, 239) <= input(41);
output(6, 240) <= input(5);
output(6, 241) <= input(6);
output(6, 242) <= input(7);
output(6, 243) <= input(8);
output(6, 244) <= input(9);
output(6, 245) <= input(10);
output(6, 246) <= input(11);
output(6, 247) <= input(12);
output(6, 248) <= input(13);
output(6, 249) <= input(14);
output(6, 250) <= input(15);
output(6, 251) <= input(34);
output(6, 252) <= input(35);
output(6, 253) <= input(38);
output(6, 254) <= input(40);
output(6, 255) <= input(42);
output(7, 0) <= input(4);
output(7, 1) <= input(5);
output(7, 2) <= input(6);
output(7, 3) <= input(7);
output(7, 4) <= input(8);
output(7, 5) <= input(9);
output(7, 6) <= input(10);
output(7, 7) <= input(11);
output(7, 8) <= input(12);
output(7, 9) <= input(13);
output(7, 10) <= input(14);
output(7, 11) <= input(15);
output(7, 12) <= input(34);
output(7, 13) <= input(35);
output(7, 14) <= input(38);
output(7, 15) <= input(40);
output(7, 16) <= input(4);
output(7, 17) <= input(5);
output(7, 18) <= input(6);
output(7, 19) <= input(7);
output(7, 20) <= input(8);
output(7, 21) <= input(9);
output(7, 22) <= input(10);
output(7, 23) <= input(11);
output(7, 24) <= input(12);
output(7, 25) <= input(13);
output(7, 26) <= input(14);
output(7, 27) <= input(15);
output(7, 28) <= input(34);
output(7, 29) <= input(35);
output(7, 30) <= input(38);
output(7, 31) <= input(40);
output(7, 32) <= input(4);
output(7, 33) <= input(5);
output(7, 34) <= input(6);
output(7, 35) <= input(7);
output(7, 36) <= input(8);
output(7, 37) <= input(9);
output(7, 38) <= input(10);
output(7, 39) <= input(11);
output(7, 40) <= input(12);
output(7, 41) <= input(13);
output(7, 42) <= input(14);
output(7, 43) <= input(15);
output(7, 44) <= input(34);
output(7, 45) <= input(35);
output(7, 46) <= input(38);
output(7, 47) <= input(40);
output(7, 48) <= input(21);
output(7, 49) <= input(22);
output(7, 50) <= input(23);
output(7, 51) <= input(24);
output(7, 52) <= input(25);
output(7, 53) <= input(26);
output(7, 54) <= input(27);
output(7, 55) <= input(28);
output(7, 56) <= input(29);
output(7, 57) <= input(30);
output(7, 58) <= input(31);
output(7, 59) <= input(33);
output(7, 60) <= input(36);
output(7, 61) <= input(37);
output(7, 62) <= input(39);
output(7, 63) <= input(41);
output(7, 64) <= input(21);
output(7, 65) <= input(22);
output(7, 66) <= input(23);
output(7, 67) <= input(24);
output(7, 68) <= input(25);
output(7, 69) <= input(26);
output(7, 70) <= input(27);
output(7, 71) <= input(28);
output(7, 72) <= input(29);
output(7, 73) <= input(30);
output(7, 74) <= input(31);
output(7, 75) <= input(33);
output(7, 76) <= input(36);
output(7, 77) <= input(37);
output(7, 78) <= input(39);
output(7, 79) <= input(41);
output(7, 80) <= input(21);
output(7, 81) <= input(22);
output(7, 82) <= input(23);
output(7, 83) <= input(24);
output(7, 84) <= input(25);
output(7, 85) <= input(26);
output(7, 86) <= input(27);
output(7, 87) <= input(28);
output(7, 88) <= input(29);
output(7, 89) <= input(30);
output(7, 90) <= input(31);
output(7, 91) <= input(33);
output(7, 92) <= input(36);
output(7, 93) <= input(37);
output(7, 94) <= input(39);
output(7, 95) <= input(41);
output(7, 96) <= input(21);
output(7, 97) <= input(22);
output(7, 98) <= input(23);
output(7, 99) <= input(24);
output(7, 100) <= input(25);
output(7, 101) <= input(26);
output(7, 102) <= input(27);
output(7, 103) <= input(28);
output(7, 104) <= input(29);
output(7, 105) <= input(30);
output(7, 106) <= input(31);
output(7, 107) <= input(33);
output(7, 108) <= input(36);
output(7, 109) <= input(37);
output(7, 110) <= input(39);
output(7, 111) <= input(41);
output(7, 112) <= input(5);
output(7, 113) <= input(6);
output(7, 114) <= input(7);
output(7, 115) <= input(8);
output(7, 116) <= input(9);
output(7, 117) <= input(10);
output(7, 118) <= input(11);
output(7, 119) <= input(12);
output(7, 120) <= input(13);
output(7, 121) <= input(14);
output(7, 122) <= input(15);
output(7, 123) <= input(34);
output(7, 124) <= input(35);
output(7, 125) <= input(38);
output(7, 126) <= input(40);
output(7, 127) <= input(42);
output(7, 128) <= input(5);
output(7, 129) <= input(6);
output(7, 130) <= input(7);
output(7, 131) <= input(8);
output(7, 132) <= input(9);
output(7, 133) <= input(10);
output(7, 134) <= input(11);
output(7, 135) <= input(12);
output(7, 136) <= input(13);
output(7, 137) <= input(14);
output(7, 138) <= input(15);
output(7, 139) <= input(34);
output(7, 140) <= input(35);
output(7, 141) <= input(38);
output(7, 142) <= input(40);
output(7, 143) <= input(42);
output(7, 144) <= input(5);
output(7, 145) <= input(6);
output(7, 146) <= input(7);
output(7, 147) <= input(8);
output(7, 148) <= input(9);
output(7, 149) <= input(10);
output(7, 150) <= input(11);
output(7, 151) <= input(12);
output(7, 152) <= input(13);
output(7, 153) <= input(14);
output(7, 154) <= input(15);
output(7, 155) <= input(34);
output(7, 156) <= input(35);
output(7, 157) <= input(38);
output(7, 158) <= input(40);
output(7, 159) <= input(42);
output(7, 160) <= input(5);
output(7, 161) <= input(6);
output(7, 162) <= input(7);
output(7, 163) <= input(8);
output(7, 164) <= input(9);
output(7, 165) <= input(10);
output(7, 166) <= input(11);
output(7, 167) <= input(12);
output(7, 168) <= input(13);
output(7, 169) <= input(14);
output(7, 170) <= input(15);
output(7, 171) <= input(34);
output(7, 172) <= input(35);
output(7, 173) <= input(38);
output(7, 174) <= input(40);
output(7, 175) <= input(42);
output(7, 176) <= input(22);
output(7, 177) <= input(23);
output(7, 178) <= input(24);
output(7, 179) <= input(25);
output(7, 180) <= input(26);
output(7, 181) <= input(27);
output(7, 182) <= input(28);
output(7, 183) <= input(29);
output(7, 184) <= input(30);
output(7, 185) <= input(31);
output(7, 186) <= input(33);
output(7, 187) <= input(36);
output(7, 188) <= input(37);
output(7, 189) <= input(39);
output(7, 190) <= input(41);
output(7, 191) <= input(43);
output(7, 192) <= input(22);
output(7, 193) <= input(23);
output(7, 194) <= input(24);
output(7, 195) <= input(25);
output(7, 196) <= input(26);
output(7, 197) <= input(27);
output(7, 198) <= input(28);
output(7, 199) <= input(29);
output(7, 200) <= input(30);
output(7, 201) <= input(31);
output(7, 202) <= input(33);
output(7, 203) <= input(36);
output(7, 204) <= input(37);
output(7, 205) <= input(39);
output(7, 206) <= input(41);
output(7, 207) <= input(43);
output(7, 208) <= input(22);
output(7, 209) <= input(23);
output(7, 210) <= input(24);
output(7, 211) <= input(25);
output(7, 212) <= input(26);
output(7, 213) <= input(27);
output(7, 214) <= input(28);
output(7, 215) <= input(29);
output(7, 216) <= input(30);
output(7, 217) <= input(31);
output(7, 218) <= input(33);
output(7, 219) <= input(36);
output(7, 220) <= input(37);
output(7, 221) <= input(39);
output(7, 222) <= input(41);
output(7, 223) <= input(43);
output(7, 224) <= input(22);
output(7, 225) <= input(23);
output(7, 226) <= input(24);
output(7, 227) <= input(25);
output(7, 228) <= input(26);
output(7, 229) <= input(27);
output(7, 230) <= input(28);
output(7, 231) <= input(29);
output(7, 232) <= input(30);
output(7, 233) <= input(31);
output(7, 234) <= input(33);
output(7, 235) <= input(36);
output(7, 236) <= input(37);
output(7, 237) <= input(39);
output(7, 238) <= input(41);
output(7, 239) <= input(43);
output(7, 240) <= input(6);
output(7, 241) <= input(7);
output(7, 242) <= input(8);
output(7, 243) <= input(9);
output(7, 244) <= input(10);
output(7, 245) <= input(11);
output(7, 246) <= input(12);
output(7, 247) <= input(13);
output(7, 248) <= input(14);
output(7, 249) <= input(15);
output(7, 250) <= input(34);
output(7, 251) <= input(35);
output(7, 252) <= input(38);
output(7, 253) <= input(40);
output(7, 254) <= input(42);
output(7, 255) <= input(44);
when "1110" =>
output(0, 0) <= input(0);
output(0, 1) <= input(1);
output(0, 2) <= input(2);
output(0, 3) <= input(3);
output(0, 4) <= input(4);
output(0, 5) <= input(5);
output(0, 6) <= input(6);
output(0, 7) <= input(7);
output(0, 8) <= input(8);
output(0, 9) <= input(9);
output(0, 10) <= input(10);
output(0, 11) <= input(11);
output(0, 12) <= input(12);
output(0, 13) <= input(13);
output(0, 14) <= input(14);
output(0, 15) <= input(15);
output(0, 16) <= input(0);
output(0, 17) <= input(1);
output(0, 18) <= input(2);
output(0, 19) <= input(3);
output(0, 20) <= input(4);
output(0, 21) <= input(5);
output(0, 22) <= input(6);
output(0, 23) <= input(7);
output(0, 24) <= input(8);
output(0, 25) <= input(9);
output(0, 26) <= input(10);
output(0, 27) <= input(11);
output(0, 28) <= input(12);
output(0, 29) <= input(13);
output(0, 30) <= input(14);
output(0, 31) <= input(15);
output(0, 32) <= input(16);
output(0, 33) <= input(17);
output(0, 34) <= input(18);
output(0, 35) <= input(19);
output(0, 36) <= input(20);
output(0, 37) <= input(21);
output(0, 38) <= input(22);
output(0, 39) <= input(23);
output(0, 40) <= input(24);
output(0, 41) <= input(25);
output(0, 42) <= input(26);
output(0, 43) <= input(27);
output(0, 44) <= input(28);
output(0, 45) <= input(29);
output(0, 46) <= input(30);
output(0, 47) <= input(31);
output(0, 48) <= input(16);
output(0, 49) <= input(17);
output(0, 50) <= input(18);
output(0, 51) <= input(19);
output(0, 52) <= input(20);
output(0, 53) <= input(21);
output(0, 54) <= input(22);
output(0, 55) <= input(23);
output(0, 56) <= input(24);
output(0, 57) <= input(25);
output(0, 58) <= input(26);
output(0, 59) <= input(27);
output(0, 60) <= input(28);
output(0, 61) <= input(29);
output(0, 62) <= input(30);
output(0, 63) <= input(31);
output(0, 64) <= input(16);
output(0, 65) <= input(17);
output(0, 66) <= input(18);
output(0, 67) <= input(19);
output(0, 68) <= input(20);
output(0, 69) <= input(21);
output(0, 70) <= input(22);
output(0, 71) <= input(23);
output(0, 72) <= input(24);
output(0, 73) <= input(25);
output(0, 74) <= input(26);
output(0, 75) <= input(27);
output(0, 76) <= input(28);
output(0, 77) <= input(29);
output(0, 78) <= input(30);
output(0, 79) <= input(31);
output(0, 80) <= input(1);
output(0, 81) <= input(2);
output(0, 82) <= input(3);
output(0, 83) <= input(4);
output(0, 84) <= input(5);
output(0, 85) <= input(6);
output(0, 86) <= input(7);
output(0, 87) <= input(8);
output(0, 88) <= input(9);
output(0, 89) <= input(10);
output(0, 90) <= input(11);
output(0, 91) <= input(12);
output(0, 92) <= input(13);
output(0, 93) <= input(14);
output(0, 94) <= input(15);
output(0, 95) <= input(32);
output(0, 96) <= input(1);
output(0, 97) <= input(2);
output(0, 98) <= input(3);
output(0, 99) <= input(4);
output(0, 100) <= input(5);
output(0, 101) <= input(6);
output(0, 102) <= input(7);
output(0, 103) <= input(8);
output(0, 104) <= input(9);
output(0, 105) <= input(10);
output(0, 106) <= input(11);
output(0, 107) <= input(12);
output(0, 108) <= input(13);
output(0, 109) <= input(14);
output(0, 110) <= input(15);
output(0, 111) <= input(32);
output(0, 112) <= input(17);
output(0, 113) <= input(18);
output(0, 114) <= input(19);
output(0, 115) <= input(20);
output(0, 116) <= input(21);
output(0, 117) <= input(22);
output(0, 118) <= input(23);
output(0, 119) <= input(24);
output(0, 120) <= input(25);
output(0, 121) <= input(26);
output(0, 122) <= input(27);
output(0, 123) <= input(28);
output(0, 124) <= input(29);
output(0, 125) <= input(30);
output(0, 126) <= input(31);
output(0, 127) <= input(33);
output(0, 128) <= input(17);
output(0, 129) <= input(18);
output(0, 130) <= input(19);
output(0, 131) <= input(20);
output(0, 132) <= input(21);
output(0, 133) <= input(22);
output(0, 134) <= input(23);
output(0, 135) <= input(24);
output(0, 136) <= input(25);
output(0, 137) <= input(26);
output(0, 138) <= input(27);
output(0, 139) <= input(28);
output(0, 140) <= input(29);
output(0, 141) <= input(30);
output(0, 142) <= input(31);
output(0, 143) <= input(33);
output(0, 144) <= input(17);
output(0, 145) <= input(18);
output(0, 146) <= input(19);
output(0, 147) <= input(20);
output(0, 148) <= input(21);
output(0, 149) <= input(22);
output(0, 150) <= input(23);
output(0, 151) <= input(24);
output(0, 152) <= input(25);
output(0, 153) <= input(26);
output(0, 154) <= input(27);
output(0, 155) <= input(28);
output(0, 156) <= input(29);
output(0, 157) <= input(30);
output(0, 158) <= input(31);
output(0, 159) <= input(33);
output(0, 160) <= input(2);
output(0, 161) <= input(3);
output(0, 162) <= input(4);
output(0, 163) <= input(5);
output(0, 164) <= input(6);
output(0, 165) <= input(7);
output(0, 166) <= input(8);
output(0, 167) <= input(9);
output(0, 168) <= input(10);
output(0, 169) <= input(11);
output(0, 170) <= input(12);
output(0, 171) <= input(13);
output(0, 172) <= input(14);
output(0, 173) <= input(15);
output(0, 174) <= input(32);
output(0, 175) <= input(34);
output(0, 176) <= input(2);
output(0, 177) <= input(3);
output(0, 178) <= input(4);
output(0, 179) <= input(5);
output(0, 180) <= input(6);
output(0, 181) <= input(7);
output(0, 182) <= input(8);
output(0, 183) <= input(9);
output(0, 184) <= input(10);
output(0, 185) <= input(11);
output(0, 186) <= input(12);
output(0, 187) <= input(13);
output(0, 188) <= input(14);
output(0, 189) <= input(15);
output(0, 190) <= input(32);
output(0, 191) <= input(34);
output(0, 192) <= input(2);
output(0, 193) <= input(3);
output(0, 194) <= input(4);
output(0, 195) <= input(5);
output(0, 196) <= input(6);
output(0, 197) <= input(7);
output(0, 198) <= input(8);
output(0, 199) <= input(9);
output(0, 200) <= input(10);
output(0, 201) <= input(11);
output(0, 202) <= input(12);
output(0, 203) <= input(13);
output(0, 204) <= input(14);
output(0, 205) <= input(15);
output(0, 206) <= input(32);
output(0, 207) <= input(34);
output(0, 208) <= input(18);
output(0, 209) <= input(19);
output(0, 210) <= input(20);
output(0, 211) <= input(21);
output(0, 212) <= input(22);
output(0, 213) <= input(23);
output(0, 214) <= input(24);
output(0, 215) <= input(25);
output(0, 216) <= input(26);
output(0, 217) <= input(27);
output(0, 218) <= input(28);
output(0, 219) <= input(29);
output(0, 220) <= input(30);
output(0, 221) <= input(31);
output(0, 222) <= input(33);
output(0, 223) <= input(35);
output(0, 224) <= input(18);
output(0, 225) <= input(19);
output(0, 226) <= input(20);
output(0, 227) <= input(21);
output(0, 228) <= input(22);
output(0, 229) <= input(23);
output(0, 230) <= input(24);
output(0, 231) <= input(25);
output(0, 232) <= input(26);
output(0, 233) <= input(27);
output(0, 234) <= input(28);
output(0, 235) <= input(29);
output(0, 236) <= input(30);
output(0, 237) <= input(31);
output(0, 238) <= input(33);
output(0, 239) <= input(35);
output(0, 240) <= input(3);
output(0, 241) <= input(4);
output(0, 242) <= input(5);
output(0, 243) <= input(6);
output(0, 244) <= input(7);
output(0, 245) <= input(8);
output(0, 246) <= input(9);
output(0, 247) <= input(10);
output(0, 248) <= input(11);
output(0, 249) <= input(12);
output(0, 250) <= input(13);
output(0, 251) <= input(14);
output(0, 252) <= input(15);
output(0, 253) <= input(32);
output(0, 254) <= input(34);
output(0, 255) <= input(36);
output(1, 0) <= input(1);
output(1, 1) <= input(2);
output(1, 2) <= input(3);
output(1, 3) <= input(4);
output(1, 4) <= input(5);
output(1, 5) <= input(6);
output(1, 6) <= input(7);
output(1, 7) <= input(8);
output(1, 8) <= input(9);
output(1, 9) <= input(10);
output(1, 10) <= input(11);
output(1, 11) <= input(12);
output(1, 12) <= input(13);
output(1, 13) <= input(14);
output(1, 14) <= input(15);
output(1, 15) <= input(32);
output(1, 16) <= input(17);
output(1, 17) <= input(18);
output(1, 18) <= input(19);
output(1, 19) <= input(20);
output(1, 20) <= input(21);
output(1, 21) <= input(22);
output(1, 22) <= input(23);
output(1, 23) <= input(24);
output(1, 24) <= input(25);
output(1, 25) <= input(26);
output(1, 26) <= input(27);
output(1, 27) <= input(28);
output(1, 28) <= input(29);
output(1, 29) <= input(30);
output(1, 30) <= input(31);
output(1, 31) <= input(33);
output(1, 32) <= input(17);
output(1, 33) <= input(18);
output(1, 34) <= input(19);
output(1, 35) <= input(20);
output(1, 36) <= input(21);
output(1, 37) <= input(22);
output(1, 38) <= input(23);
output(1, 39) <= input(24);
output(1, 40) <= input(25);
output(1, 41) <= input(26);
output(1, 42) <= input(27);
output(1, 43) <= input(28);
output(1, 44) <= input(29);
output(1, 45) <= input(30);
output(1, 46) <= input(31);
output(1, 47) <= input(33);
output(1, 48) <= input(2);
output(1, 49) <= input(3);
output(1, 50) <= input(4);
output(1, 51) <= input(5);
output(1, 52) <= input(6);
output(1, 53) <= input(7);
output(1, 54) <= input(8);
output(1, 55) <= input(9);
output(1, 56) <= input(10);
output(1, 57) <= input(11);
output(1, 58) <= input(12);
output(1, 59) <= input(13);
output(1, 60) <= input(14);
output(1, 61) <= input(15);
output(1, 62) <= input(32);
output(1, 63) <= input(34);
output(1, 64) <= input(2);
output(1, 65) <= input(3);
output(1, 66) <= input(4);
output(1, 67) <= input(5);
output(1, 68) <= input(6);
output(1, 69) <= input(7);
output(1, 70) <= input(8);
output(1, 71) <= input(9);
output(1, 72) <= input(10);
output(1, 73) <= input(11);
output(1, 74) <= input(12);
output(1, 75) <= input(13);
output(1, 76) <= input(14);
output(1, 77) <= input(15);
output(1, 78) <= input(32);
output(1, 79) <= input(34);
output(1, 80) <= input(18);
output(1, 81) <= input(19);
output(1, 82) <= input(20);
output(1, 83) <= input(21);
output(1, 84) <= input(22);
output(1, 85) <= input(23);
output(1, 86) <= input(24);
output(1, 87) <= input(25);
output(1, 88) <= input(26);
output(1, 89) <= input(27);
output(1, 90) <= input(28);
output(1, 91) <= input(29);
output(1, 92) <= input(30);
output(1, 93) <= input(31);
output(1, 94) <= input(33);
output(1, 95) <= input(35);
output(1, 96) <= input(18);
output(1, 97) <= input(19);
output(1, 98) <= input(20);
output(1, 99) <= input(21);
output(1, 100) <= input(22);
output(1, 101) <= input(23);
output(1, 102) <= input(24);
output(1, 103) <= input(25);
output(1, 104) <= input(26);
output(1, 105) <= input(27);
output(1, 106) <= input(28);
output(1, 107) <= input(29);
output(1, 108) <= input(30);
output(1, 109) <= input(31);
output(1, 110) <= input(33);
output(1, 111) <= input(35);
output(1, 112) <= input(3);
output(1, 113) <= input(4);
output(1, 114) <= input(5);
output(1, 115) <= input(6);
output(1, 116) <= input(7);
output(1, 117) <= input(8);
output(1, 118) <= input(9);
output(1, 119) <= input(10);
output(1, 120) <= input(11);
output(1, 121) <= input(12);
output(1, 122) <= input(13);
output(1, 123) <= input(14);
output(1, 124) <= input(15);
output(1, 125) <= input(32);
output(1, 126) <= input(34);
output(1, 127) <= input(36);
output(1, 128) <= input(3);
output(1, 129) <= input(4);
output(1, 130) <= input(5);
output(1, 131) <= input(6);
output(1, 132) <= input(7);
output(1, 133) <= input(8);
output(1, 134) <= input(9);
output(1, 135) <= input(10);
output(1, 136) <= input(11);
output(1, 137) <= input(12);
output(1, 138) <= input(13);
output(1, 139) <= input(14);
output(1, 140) <= input(15);
output(1, 141) <= input(32);
output(1, 142) <= input(34);
output(1, 143) <= input(36);
output(1, 144) <= input(19);
output(1, 145) <= input(20);
output(1, 146) <= input(21);
output(1, 147) <= input(22);
output(1, 148) <= input(23);
output(1, 149) <= input(24);
output(1, 150) <= input(25);
output(1, 151) <= input(26);
output(1, 152) <= input(27);
output(1, 153) <= input(28);
output(1, 154) <= input(29);
output(1, 155) <= input(30);
output(1, 156) <= input(31);
output(1, 157) <= input(33);
output(1, 158) <= input(35);
output(1, 159) <= input(37);
output(1, 160) <= input(19);
output(1, 161) <= input(20);
output(1, 162) <= input(21);
output(1, 163) <= input(22);
output(1, 164) <= input(23);
output(1, 165) <= input(24);
output(1, 166) <= input(25);
output(1, 167) <= input(26);
output(1, 168) <= input(27);
output(1, 169) <= input(28);
output(1, 170) <= input(29);
output(1, 171) <= input(30);
output(1, 172) <= input(31);
output(1, 173) <= input(33);
output(1, 174) <= input(35);
output(1, 175) <= input(37);
output(1, 176) <= input(4);
output(1, 177) <= input(5);
output(1, 178) <= input(6);
output(1, 179) <= input(7);
output(1, 180) <= input(8);
output(1, 181) <= input(9);
output(1, 182) <= input(10);
output(1, 183) <= input(11);
output(1, 184) <= input(12);
output(1, 185) <= input(13);
output(1, 186) <= input(14);
output(1, 187) <= input(15);
output(1, 188) <= input(32);
output(1, 189) <= input(34);
output(1, 190) <= input(36);
output(1, 191) <= input(38);
output(1, 192) <= input(4);
output(1, 193) <= input(5);
output(1, 194) <= input(6);
output(1, 195) <= input(7);
output(1, 196) <= input(8);
output(1, 197) <= input(9);
output(1, 198) <= input(10);
output(1, 199) <= input(11);
output(1, 200) <= input(12);
output(1, 201) <= input(13);
output(1, 202) <= input(14);
output(1, 203) <= input(15);
output(1, 204) <= input(32);
output(1, 205) <= input(34);
output(1, 206) <= input(36);
output(1, 207) <= input(38);
output(1, 208) <= input(20);
output(1, 209) <= input(21);
output(1, 210) <= input(22);
output(1, 211) <= input(23);
output(1, 212) <= input(24);
output(1, 213) <= input(25);
output(1, 214) <= input(26);
output(1, 215) <= input(27);
output(1, 216) <= input(28);
output(1, 217) <= input(29);
output(1, 218) <= input(30);
output(1, 219) <= input(31);
output(1, 220) <= input(33);
output(1, 221) <= input(35);
output(1, 222) <= input(37);
output(1, 223) <= input(39);
output(1, 224) <= input(20);
output(1, 225) <= input(21);
output(1, 226) <= input(22);
output(1, 227) <= input(23);
output(1, 228) <= input(24);
output(1, 229) <= input(25);
output(1, 230) <= input(26);
output(1, 231) <= input(27);
output(1, 232) <= input(28);
output(1, 233) <= input(29);
output(1, 234) <= input(30);
output(1, 235) <= input(31);
output(1, 236) <= input(33);
output(1, 237) <= input(35);
output(1, 238) <= input(37);
output(1, 239) <= input(39);
output(1, 240) <= input(5);
output(1, 241) <= input(6);
output(1, 242) <= input(7);
output(1, 243) <= input(8);
output(1, 244) <= input(9);
output(1, 245) <= input(10);
output(1, 246) <= input(11);
output(1, 247) <= input(12);
output(1, 248) <= input(13);
output(1, 249) <= input(14);
output(1, 250) <= input(15);
output(1, 251) <= input(32);
output(1, 252) <= input(34);
output(1, 253) <= input(36);
output(1, 254) <= input(38);
output(1, 255) <= input(40);
output(2, 0) <= input(2);
output(2, 1) <= input(3);
output(2, 2) <= input(4);
output(2, 3) <= input(5);
output(2, 4) <= input(6);
output(2, 5) <= input(7);
output(2, 6) <= input(8);
output(2, 7) <= input(9);
output(2, 8) <= input(10);
output(2, 9) <= input(11);
output(2, 10) <= input(12);
output(2, 11) <= input(13);
output(2, 12) <= input(14);
output(2, 13) <= input(15);
output(2, 14) <= input(32);
output(2, 15) <= input(34);
output(2, 16) <= input(18);
output(2, 17) <= input(19);
output(2, 18) <= input(20);
output(2, 19) <= input(21);
output(2, 20) <= input(22);
output(2, 21) <= input(23);
output(2, 22) <= input(24);
output(2, 23) <= input(25);
output(2, 24) <= input(26);
output(2, 25) <= input(27);
output(2, 26) <= input(28);
output(2, 27) <= input(29);
output(2, 28) <= input(30);
output(2, 29) <= input(31);
output(2, 30) <= input(33);
output(2, 31) <= input(35);
output(2, 32) <= input(18);
output(2, 33) <= input(19);
output(2, 34) <= input(20);
output(2, 35) <= input(21);
output(2, 36) <= input(22);
output(2, 37) <= input(23);
output(2, 38) <= input(24);
output(2, 39) <= input(25);
output(2, 40) <= input(26);
output(2, 41) <= input(27);
output(2, 42) <= input(28);
output(2, 43) <= input(29);
output(2, 44) <= input(30);
output(2, 45) <= input(31);
output(2, 46) <= input(33);
output(2, 47) <= input(35);
output(2, 48) <= input(3);
output(2, 49) <= input(4);
output(2, 50) <= input(5);
output(2, 51) <= input(6);
output(2, 52) <= input(7);
output(2, 53) <= input(8);
output(2, 54) <= input(9);
output(2, 55) <= input(10);
output(2, 56) <= input(11);
output(2, 57) <= input(12);
output(2, 58) <= input(13);
output(2, 59) <= input(14);
output(2, 60) <= input(15);
output(2, 61) <= input(32);
output(2, 62) <= input(34);
output(2, 63) <= input(36);
output(2, 64) <= input(19);
output(2, 65) <= input(20);
output(2, 66) <= input(21);
output(2, 67) <= input(22);
output(2, 68) <= input(23);
output(2, 69) <= input(24);
output(2, 70) <= input(25);
output(2, 71) <= input(26);
output(2, 72) <= input(27);
output(2, 73) <= input(28);
output(2, 74) <= input(29);
output(2, 75) <= input(30);
output(2, 76) <= input(31);
output(2, 77) <= input(33);
output(2, 78) <= input(35);
output(2, 79) <= input(37);
output(2, 80) <= input(19);
output(2, 81) <= input(20);
output(2, 82) <= input(21);
output(2, 83) <= input(22);
output(2, 84) <= input(23);
output(2, 85) <= input(24);
output(2, 86) <= input(25);
output(2, 87) <= input(26);
output(2, 88) <= input(27);
output(2, 89) <= input(28);
output(2, 90) <= input(29);
output(2, 91) <= input(30);
output(2, 92) <= input(31);
output(2, 93) <= input(33);
output(2, 94) <= input(35);
output(2, 95) <= input(37);
output(2, 96) <= input(4);
output(2, 97) <= input(5);
output(2, 98) <= input(6);
output(2, 99) <= input(7);
output(2, 100) <= input(8);
output(2, 101) <= input(9);
output(2, 102) <= input(10);
output(2, 103) <= input(11);
output(2, 104) <= input(12);
output(2, 105) <= input(13);
output(2, 106) <= input(14);
output(2, 107) <= input(15);
output(2, 108) <= input(32);
output(2, 109) <= input(34);
output(2, 110) <= input(36);
output(2, 111) <= input(38);
output(2, 112) <= input(20);
output(2, 113) <= input(21);
output(2, 114) <= input(22);
output(2, 115) <= input(23);
output(2, 116) <= input(24);
output(2, 117) <= input(25);
output(2, 118) <= input(26);
output(2, 119) <= input(27);
output(2, 120) <= input(28);
output(2, 121) <= input(29);
output(2, 122) <= input(30);
output(2, 123) <= input(31);
output(2, 124) <= input(33);
output(2, 125) <= input(35);
output(2, 126) <= input(37);
output(2, 127) <= input(39);
output(2, 128) <= input(20);
output(2, 129) <= input(21);
output(2, 130) <= input(22);
output(2, 131) <= input(23);
output(2, 132) <= input(24);
output(2, 133) <= input(25);
output(2, 134) <= input(26);
output(2, 135) <= input(27);
output(2, 136) <= input(28);
output(2, 137) <= input(29);
output(2, 138) <= input(30);
output(2, 139) <= input(31);
output(2, 140) <= input(33);
output(2, 141) <= input(35);
output(2, 142) <= input(37);
output(2, 143) <= input(39);
output(2, 144) <= input(5);
output(2, 145) <= input(6);
output(2, 146) <= input(7);
output(2, 147) <= input(8);
output(2, 148) <= input(9);
output(2, 149) <= input(10);
output(2, 150) <= input(11);
output(2, 151) <= input(12);
output(2, 152) <= input(13);
output(2, 153) <= input(14);
output(2, 154) <= input(15);
output(2, 155) <= input(32);
output(2, 156) <= input(34);
output(2, 157) <= input(36);
output(2, 158) <= input(38);
output(2, 159) <= input(40);
output(2, 160) <= input(5);
output(2, 161) <= input(6);
output(2, 162) <= input(7);
output(2, 163) <= input(8);
output(2, 164) <= input(9);
output(2, 165) <= input(10);
output(2, 166) <= input(11);
output(2, 167) <= input(12);
output(2, 168) <= input(13);
output(2, 169) <= input(14);
output(2, 170) <= input(15);
output(2, 171) <= input(32);
output(2, 172) <= input(34);
output(2, 173) <= input(36);
output(2, 174) <= input(38);
output(2, 175) <= input(40);
output(2, 176) <= input(21);
output(2, 177) <= input(22);
output(2, 178) <= input(23);
output(2, 179) <= input(24);
output(2, 180) <= input(25);
output(2, 181) <= input(26);
output(2, 182) <= input(27);
output(2, 183) <= input(28);
output(2, 184) <= input(29);
output(2, 185) <= input(30);
output(2, 186) <= input(31);
output(2, 187) <= input(33);
output(2, 188) <= input(35);
output(2, 189) <= input(37);
output(2, 190) <= input(39);
output(2, 191) <= input(41);
output(2, 192) <= input(6);
output(2, 193) <= input(7);
output(2, 194) <= input(8);
output(2, 195) <= input(9);
output(2, 196) <= input(10);
output(2, 197) <= input(11);
output(2, 198) <= input(12);
output(2, 199) <= input(13);
output(2, 200) <= input(14);
output(2, 201) <= input(15);
output(2, 202) <= input(32);
output(2, 203) <= input(34);
output(2, 204) <= input(36);
output(2, 205) <= input(38);
output(2, 206) <= input(40);
output(2, 207) <= input(42);
output(2, 208) <= input(6);
output(2, 209) <= input(7);
output(2, 210) <= input(8);
output(2, 211) <= input(9);
output(2, 212) <= input(10);
output(2, 213) <= input(11);
output(2, 214) <= input(12);
output(2, 215) <= input(13);
output(2, 216) <= input(14);
output(2, 217) <= input(15);
output(2, 218) <= input(32);
output(2, 219) <= input(34);
output(2, 220) <= input(36);
output(2, 221) <= input(38);
output(2, 222) <= input(40);
output(2, 223) <= input(42);
output(2, 224) <= input(22);
output(2, 225) <= input(23);
output(2, 226) <= input(24);
output(2, 227) <= input(25);
output(2, 228) <= input(26);
output(2, 229) <= input(27);
output(2, 230) <= input(28);
output(2, 231) <= input(29);
output(2, 232) <= input(30);
output(2, 233) <= input(31);
output(2, 234) <= input(33);
output(2, 235) <= input(35);
output(2, 236) <= input(37);
output(2, 237) <= input(39);
output(2, 238) <= input(41);
output(2, 239) <= input(43);
output(2, 240) <= input(7);
output(2, 241) <= input(8);
output(2, 242) <= input(9);
output(2, 243) <= input(10);
output(2, 244) <= input(11);
output(2, 245) <= input(12);
output(2, 246) <= input(13);
output(2, 247) <= input(14);
output(2, 248) <= input(15);
output(2, 249) <= input(32);
output(2, 250) <= input(34);
output(2, 251) <= input(36);
output(2, 252) <= input(38);
output(2, 253) <= input(40);
output(2, 254) <= input(42);
output(2, 255) <= input(44);
output(3, 0) <= input(3);
output(3, 1) <= input(4);
output(3, 2) <= input(5);
output(3, 3) <= input(6);
output(3, 4) <= input(7);
output(3, 5) <= input(8);
output(3, 6) <= input(9);
output(3, 7) <= input(10);
output(3, 8) <= input(11);
output(3, 9) <= input(12);
output(3, 10) <= input(13);
output(3, 11) <= input(14);
output(3, 12) <= input(15);
output(3, 13) <= input(32);
output(3, 14) <= input(34);
output(3, 15) <= input(36);
output(3, 16) <= input(19);
output(3, 17) <= input(20);
output(3, 18) <= input(21);
output(3, 19) <= input(22);
output(3, 20) <= input(23);
output(3, 21) <= input(24);
output(3, 22) <= input(25);
output(3, 23) <= input(26);
output(3, 24) <= input(27);
output(3, 25) <= input(28);
output(3, 26) <= input(29);
output(3, 27) <= input(30);
output(3, 28) <= input(31);
output(3, 29) <= input(33);
output(3, 30) <= input(35);
output(3, 31) <= input(37);
output(3, 32) <= input(4);
output(3, 33) <= input(5);
output(3, 34) <= input(6);
output(3, 35) <= input(7);
output(3, 36) <= input(8);
output(3, 37) <= input(9);
output(3, 38) <= input(10);
output(3, 39) <= input(11);
output(3, 40) <= input(12);
output(3, 41) <= input(13);
output(3, 42) <= input(14);
output(3, 43) <= input(15);
output(3, 44) <= input(32);
output(3, 45) <= input(34);
output(3, 46) <= input(36);
output(3, 47) <= input(38);
output(3, 48) <= input(20);
output(3, 49) <= input(21);
output(3, 50) <= input(22);
output(3, 51) <= input(23);
output(3, 52) <= input(24);
output(3, 53) <= input(25);
output(3, 54) <= input(26);
output(3, 55) <= input(27);
output(3, 56) <= input(28);
output(3, 57) <= input(29);
output(3, 58) <= input(30);
output(3, 59) <= input(31);
output(3, 60) <= input(33);
output(3, 61) <= input(35);
output(3, 62) <= input(37);
output(3, 63) <= input(39);
output(3, 64) <= input(20);
output(3, 65) <= input(21);
output(3, 66) <= input(22);
output(3, 67) <= input(23);
output(3, 68) <= input(24);
output(3, 69) <= input(25);
output(3, 70) <= input(26);
output(3, 71) <= input(27);
output(3, 72) <= input(28);
output(3, 73) <= input(29);
output(3, 74) <= input(30);
output(3, 75) <= input(31);
output(3, 76) <= input(33);
output(3, 77) <= input(35);
output(3, 78) <= input(37);
output(3, 79) <= input(39);
output(3, 80) <= input(5);
output(3, 81) <= input(6);
output(3, 82) <= input(7);
output(3, 83) <= input(8);
output(3, 84) <= input(9);
output(3, 85) <= input(10);
output(3, 86) <= input(11);
output(3, 87) <= input(12);
output(3, 88) <= input(13);
output(3, 89) <= input(14);
output(3, 90) <= input(15);
output(3, 91) <= input(32);
output(3, 92) <= input(34);
output(3, 93) <= input(36);
output(3, 94) <= input(38);
output(3, 95) <= input(40);
output(3, 96) <= input(21);
output(3, 97) <= input(22);
output(3, 98) <= input(23);
output(3, 99) <= input(24);
output(3, 100) <= input(25);
output(3, 101) <= input(26);
output(3, 102) <= input(27);
output(3, 103) <= input(28);
output(3, 104) <= input(29);
output(3, 105) <= input(30);
output(3, 106) <= input(31);
output(3, 107) <= input(33);
output(3, 108) <= input(35);
output(3, 109) <= input(37);
output(3, 110) <= input(39);
output(3, 111) <= input(41);
output(3, 112) <= input(6);
output(3, 113) <= input(7);
output(3, 114) <= input(8);
output(3, 115) <= input(9);
output(3, 116) <= input(10);
output(3, 117) <= input(11);
output(3, 118) <= input(12);
output(3, 119) <= input(13);
output(3, 120) <= input(14);
output(3, 121) <= input(15);
output(3, 122) <= input(32);
output(3, 123) <= input(34);
output(3, 124) <= input(36);
output(3, 125) <= input(38);
output(3, 126) <= input(40);
output(3, 127) <= input(42);
output(3, 128) <= input(6);
output(3, 129) <= input(7);
output(3, 130) <= input(8);
output(3, 131) <= input(9);
output(3, 132) <= input(10);
output(3, 133) <= input(11);
output(3, 134) <= input(12);
output(3, 135) <= input(13);
output(3, 136) <= input(14);
output(3, 137) <= input(15);
output(3, 138) <= input(32);
output(3, 139) <= input(34);
output(3, 140) <= input(36);
output(3, 141) <= input(38);
output(3, 142) <= input(40);
output(3, 143) <= input(42);
output(3, 144) <= input(22);
output(3, 145) <= input(23);
output(3, 146) <= input(24);
output(3, 147) <= input(25);
output(3, 148) <= input(26);
output(3, 149) <= input(27);
output(3, 150) <= input(28);
output(3, 151) <= input(29);
output(3, 152) <= input(30);
output(3, 153) <= input(31);
output(3, 154) <= input(33);
output(3, 155) <= input(35);
output(3, 156) <= input(37);
output(3, 157) <= input(39);
output(3, 158) <= input(41);
output(3, 159) <= input(43);
output(3, 160) <= input(7);
output(3, 161) <= input(8);
output(3, 162) <= input(9);
output(3, 163) <= input(10);
output(3, 164) <= input(11);
output(3, 165) <= input(12);
output(3, 166) <= input(13);
output(3, 167) <= input(14);
output(3, 168) <= input(15);
output(3, 169) <= input(32);
output(3, 170) <= input(34);
output(3, 171) <= input(36);
output(3, 172) <= input(38);
output(3, 173) <= input(40);
output(3, 174) <= input(42);
output(3, 175) <= input(44);
output(3, 176) <= input(23);
output(3, 177) <= input(24);
output(3, 178) <= input(25);
output(3, 179) <= input(26);
output(3, 180) <= input(27);
output(3, 181) <= input(28);
output(3, 182) <= input(29);
output(3, 183) <= input(30);
output(3, 184) <= input(31);
output(3, 185) <= input(33);
output(3, 186) <= input(35);
output(3, 187) <= input(37);
output(3, 188) <= input(39);
output(3, 189) <= input(41);
output(3, 190) <= input(43);
output(3, 191) <= input(45);
output(3, 192) <= input(23);
output(3, 193) <= input(24);
output(3, 194) <= input(25);
output(3, 195) <= input(26);
output(3, 196) <= input(27);
output(3, 197) <= input(28);
output(3, 198) <= input(29);
output(3, 199) <= input(30);
output(3, 200) <= input(31);
output(3, 201) <= input(33);
output(3, 202) <= input(35);
output(3, 203) <= input(37);
output(3, 204) <= input(39);
output(3, 205) <= input(41);
output(3, 206) <= input(43);
output(3, 207) <= input(45);
output(3, 208) <= input(8);
output(3, 209) <= input(9);
output(3, 210) <= input(10);
output(3, 211) <= input(11);
output(3, 212) <= input(12);
output(3, 213) <= input(13);
output(3, 214) <= input(14);
output(3, 215) <= input(15);
output(3, 216) <= input(32);
output(3, 217) <= input(34);
output(3, 218) <= input(36);
output(3, 219) <= input(38);
output(3, 220) <= input(40);
output(3, 221) <= input(42);
output(3, 222) <= input(44);
output(3, 223) <= input(46);
output(3, 224) <= input(24);
output(3, 225) <= input(25);
output(3, 226) <= input(26);
output(3, 227) <= input(27);
output(3, 228) <= input(28);
output(3, 229) <= input(29);
output(3, 230) <= input(30);
output(3, 231) <= input(31);
output(3, 232) <= input(33);
output(3, 233) <= input(35);
output(3, 234) <= input(37);
output(3, 235) <= input(39);
output(3, 236) <= input(41);
output(3, 237) <= input(43);
output(3, 238) <= input(45);
output(3, 239) <= input(47);
output(3, 240) <= input(9);
output(3, 241) <= input(10);
output(3, 242) <= input(11);
output(3, 243) <= input(12);
output(3, 244) <= input(13);
output(3, 245) <= input(14);
output(3, 246) <= input(15);
output(3, 247) <= input(32);
output(3, 248) <= input(34);
output(3, 249) <= input(36);
output(3, 250) <= input(38);
output(3, 251) <= input(40);
output(3, 252) <= input(42);
output(3, 253) <= input(44);
output(3, 254) <= input(46);
output(3, 255) <= input(48);
output(4, 0) <= input(4);
output(4, 1) <= input(5);
output(4, 2) <= input(6);
output(4, 3) <= input(7);
output(4, 4) <= input(8);
output(4, 5) <= input(9);
output(4, 6) <= input(10);
output(4, 7) <= input(11);
output(4, 8) <= input(12);
output(4, 9) <= input(13);
output(4, 10) <= input(14);
output(4, 11) <= input(15);
output(4, 12) <= input(32);
output(4, 13) <= input(34);
output(4, 14) <= input(36);
output(4, 15) <= input(38);
output(4, 16) <= input(20);
output(4, 17) <= input(21);
output(4, 18) <= input(22);
output(4, 19) <= input(23);
output(4, 20) <= input(24);
output(4, 21) <= input(25);
output(4, 22) <= input(26);
output(4, 23) <= input(27);
output(4, 24) <= input(28);
output(4, 25) <= input(29);
output(4, 26) <= input(30);
output(4, 27) <= input(31);
output(4, 28) <= input(33);
output(4, 29) <= input(35);
output(4, 30) <= input(37);
output(4, 31) <= input(39);
output(4, 32) <= input(5);
output(4, 33) <= input(6);
output(4, 34) <= input(7);
output(4, 35) <= input(8);
output(4, 36) <= input(9);
output(4, 37) <= input(10);
output(4, 38) <= input(11);
output(4, 39) <= input(12);
output(4, 40) <= input(13);
output(4, 41) <= input(14);
output(4, 42) <= input(15);
output(4, 43) <= input(32);
output(4, 44) <= input(34);
output(4, 45) <= input(36);
output(4, 46) <= input(38);
output(4, 47) <= input(40);
output(4, 48) <= input(21);
output(4, 49) <= input(22);
output(4, 50) <= input(23);
output(4, 51) <= input(24);
output(4, 52) <= input(25);
output(4, 53) <= input(26);
output(4, 54) <= input(27);
output(4, 55) <= input(28);
output(4, 56) <= input(29);
output(4, 57) <= input(30);
output(4, 58) <= input(31);
output(4, 59) <= input(33);
output(4, 60) <= input(35);
output(4, 61) <= input(37);
output(4, 62) <= input(39);
output(4, 63) <= input(41);
output(4, 64) <= input(6);
output(4, 65) <= input(7);
output(4, 66) <= input(8);
output(4, 67) <= input(9);
output(4, 68) <= input(10);
output(4, 69) <= input(11);
output(4, 70) <= input(12);
output(4, 71) <= input(13);
output(4, 72) <= input(14);
output(4, 73) <= input(15);
output(4, 74) <= input(32);
output(4, 75) <= input(34);
output(4, 76) <= input(36);
output(4, 77) <= input(38);
output(4, 78) <= input(40);
output(4, 79) <= input(42);
output(4, 80) <= input(22);
output(4, 81) <= input(23);
output(4, 82) <= input(24);
output(4, 83) <= input(25);
output(4, 84) <= input(26);
output(4, 85) <= input(27);
output(4, 86) <= input(28);
output(4, 87) <= input(29);
output(4, 88) <= input(30);
output(4, 89) <= input(31);
output(4, 90) <= input(33);
output(4, 91) <= input(35);
output(4, 92) <= input(37);
output(4, 93) <= input(39);
output(4, 94) <= input(41);
output(4, 95) <= input(43);
output(4, 96) <= input(7);
output(4, 97) <= input(8);
output(4, 98) <= input(9);
output(4, 99) <= input(10);
output(4, 100) <= input(11);
output(4, 101) <= input(12);
output(4, 102) <= input(13);
output(4, 103) <= input(14);
output(4, 104) <= input(15);
output(4, 105) <= input(32);
output(4, 106) <= input(34);
output(4, 107) <= input(36);
output(4, 108) <= input(38);
output(4, 109) <= input(40);
output(4, 110) <= input(42);
output(4, 111) <= input(44);
output(4, 112) <= input(23);
output(4, 113) <= input(24);
output(4, 114) <= input(25);
output(4, 115) <= input(26);
output(4, 116) <= input(27);
output(4, 117) <= input(28);
output(4, 118) <= input(29);
output(4, 119) <= input(30);
output(4, 120) <= input(31);
output(4, 121) <= input(33);
output(4, 122) <= input(35);
output(4, 123) <= input(37);
output(4, 124) <= input(39);
output(4, 125) <= input(41);
output(4, 126) <= input(43);
output(4, 127) <= input(45);
output(4, 128) <= input(23);
output(4, 129) <= input(24);
output(4, 130) <= input(25);
output(4, 131) <= input(26);
output(4, 132) <= input(27);
output(4, 133) <= input(28);
output(4, 134) <= input(29);
output(4, 135) <= input(30);
output(4, 136) <= input(31);
output(4, 137) <= input(33);
output(4, 138) <= input(35);
output(4, 139) <= input(37);
output(4, 140) <= input(39);
output(4, 141) <= input(41);
output(4, 142) <= input(43);
output(4, 143) <= input(45);
output(4, 144) <= input(8);
output(4, 145) <= input(9);
output(4, 146) <= input(10);
output(4, 147) <= input(11);
output(4, 148) <= input(12);
output(4, 149) <= input(13);
output(4, 150) <= input(14);
output(4, 151) <= input(15);
output(4, 152) <= input(32);
output(4, 153) <= input(34);
output(4, 154) <= input(36);
output(4, 155) <= input(38);
output(4, 156) <= input(40);
output(4, 157) <= input(42);
output(4, 158) <= input(44);
output(4, 159) <= input(46);
output(4, 160) <= input(24);
output(4, 161) <= input(25);
output(4, 162) <= input(26);
output(4, 163) <= input(27);
output(4, 164) <= input(28);
output(4, 165) <= input(29);
output(4, 166) <= input(30);
output(4, 167) <= input(31);
output(4, 168) <= input(33);
output(4, 169) <= input(35);
output(4, 170) <= input(37);
output(4, 171) <= input(39);
output(4, 172) <= input(41);
output(4, 173) <= input(43);
output(4, 174) <= input(45);
output(4, 175) <= input(47);
output(4, 176) <= input(9);
output(4, 177) <= input(10);
output(4, 178) <= input(11);
output(4, 179) <= input(12);
output(4, 180) <= input(13);
output(4, 181) <= input(14);
output(4, 182) <= input(15);
output(4, 183) <= input(32);
output(4, 184) <= input(34);
output(4, 185) <= input(36);
output(4, 186) <= input(38);
output(4, 187) <= input(40);
output(4, 188) <= input(42);
output(4, 189) <= input(44);
output(4, 190) <= input(46);
output(4, 191) <= input(48);
output(4, 192) <= input(25);
output(4, 193) <= input(26);
output(4, 194) <= input(27);
output(4, 195) <= input(28);
output(4, 196) <= input(29);
output(4, 197) <= input(30);
output(4, 198) <= input(31);
output(4, 199) <= input(33);
output(4, 200) <= input(35);
output(4, 201) <= input(37);
output(4, 202) <= input(39);
output(4, 203) <= input(41);
output(4, 204) <= input(43);
output(4, 205) <= input(45);
output(4, 206) <= input(47);
output(4, 207) <= input(49);
output(4, 208) <= input(10);
output(4, 209) <= input(11);
output(4, 210) <= input(12);
output(4, 211) <= input(13);
output(4, 212) <= input(14);
output(4, 213) <= input(15);
output(4, 214) <= input(32);
output(4, 215) <= input(34);
output(4, 216) <= input(36);
output(4, 217) <= input(38);
output(4, 218) <= input(40);
output(4, 219) <= input(42);
output(4, 220) <= input(44);
output(4, 221) <= input(46);
output(4, 222) <= input(48);
output(4, 223) <= input(50);
output(4, 224) <= input(26);
output(4, 225) <= input(27);
output(4, 226) <= input(28);
output(4, 227) <= input(29);
output(4, 228) <= input(30);
output(4, 229) <= input(31);
output(4, 230) <= input(33);
output(4, 231) <= input(35);
output(4, 232) <= input(37);
output(4, 233) <= input(39);
output(4, 234) <= input(41);
output(4, 235) <= input(43);
output(4, 236) <= input(45);
output(4, 237) <= input(47);
output(4, 238) <= input(49);
output(4, 239) <= input(51);
output(4, 240) <= input(11);
output(4, 241) <= input(12);
output(4, 242) <= input(13);
output(4, 243) <= input(14);
output(4, 244) <= input(15);
output(4, 245) <= input(32);
output(4, 246) <= input(34);
output(4, 247) <= input(36);
output(4, 248) <= input(38);
output(4, 249) <= input(40);
output(4, 250) <= input(42);
output(4, 251) <= input(44);
output(4, 252) <= input(46);
output(4, 253) <= input(48);
output(4, 254) <= input(50);
output(4, 255) <= input(52);
output(5, 0) <= input(21);
output(5, 1) <= input(22);
output(5, 2) <= input(23);
output(5, 3) <= input(24);
output(5, 4) <= input(25);
output(5, 5) <= input(26);
output(5, 6) <= input(27);
output(5, 7) <= input(28);
output(5, 8) <= input(29);
output(5, 9) <= input(30);
output(5, 10) <= input(31);
output(5, 11) <= input(33);
output(5, 12) <= input(35);
output(5, 13) <= input(37);
output(5, 14) <= input(39);
output(5, 15) <= input(41);
output(5, 16) <= input(6);
output(5, 17) <= input(7);
output(5, 18) <= input(8);
output(5, 19) <= input(9);
output(5, 20) <= input(10);
output(5, 21) <= input(11);
output(5, 22) <= input(12);
output(5, 23) <= input(13);
output(5, 24) <= input(14);
output(5, 25) <= input(15);
output(5, 26) <= input(32);
output(5, 27) <= input(34);
output(5, 28) <= input(36);
output(5, 29) <= input(38);
output(5, 30) <= input(40);
output(5, 31) <= input(42);
output(5, 32) <= input(22);
output(5, 33) <= input(23);
output(5, 34) <= input(24);
output(5, 35) <= input(25);
output(5, 36) <= input(26);
output(5, 37) <= input(27);
output(5, 38) <= input(28);
output(5, 39) <= input(29);
output(5, 40) <= input(30);
output(5, 41) <= input(31);
output(5, 42) <= input(33);
output(5, 43) <= input(35);
output(5, 44) <= input(37);
output(5, 45) <= input(39);
output(5, 46) <= input(41);
output(5, 47) <= input(43);
output(5, 48) <= input(7);
output(5, 49) <= input(8);
output(5, 50) <= input(9);
output(5, 51) <= input(10);
output(5, 52) <= input(11);
output(5, 53) <= input(12);
output(5, 54) <= input(13);
output(5, 55) <= input(14);
output(5, 56) <= input(15);
output(5, 57) <= input(32);
output(5, 58) <= input(34);
output(5, 59) <= input(36);
output(5, 60) <= input(38);
output(5, 61) <= input(40);
output(5, 62) <= input(42);
output(5, 63) <= input(44);
output(5, 64) <= input(23);
output(5, 65) <= input(24);
output(5, 66) <= input(25);
output(5, 67) <= input(26);
output(5, 68) <= input(27);
output(5, 69) <= input(28);
output(5, 70) <= input(29);
output(5, 71) <= input(30);
output(5, 72) <= input(31);
output(5, 73) <= input(33);
output(5, 74) <= input(35);
output(5, 75) <= input(37);
output(5, 76) <= input(39);
output(5, 77) <= input(41);
output(5, 78) <= input(43);
output(5, 79) <= input(45);
output(5, 80) <= input(8);
output(5, 81) <= input(9);
output(5, 82) <= input(10);
output(5, 83) <= input(11);
output(5, 84) <= input(12);
output(5, 85) <= input(13);
output(5, 86) <= input(14);
output(5, 87) <= input(15);
output(5, 88) <= input(32);
output(5, 89) <= input(34);
output(5, 90) <= input(36);
output(5, 91) <= input(38);
output(5, 92) <= input(40);
output(5, 93) <= input(42);
output(5, 94) <= input(44);
output(5, 95) <= input(46);
output(5, 96) <= input(24);
output(5, 97) <= input(25);
output(5, 98) <= input(26);
output(5, 99) <= input(27);
output(5, 100) <= input(28);
output(5, 101) <= input(29);
output(5, 102) <= input(30);
output(5, 103) <= input(31);
output(5, 104) <= input(33);
output(5, 105) <= input(35);
output(5, 106) <= input(37);
output(5, 107) <= input(39);
output(5, 108) <= input(41);
output(5, 109) <= input(43);
output(5, 110) <= input(45);
output(5, 111) <= input(47);
output(5, 112) <= input(9);
output(5, 113) <= input(10);
output(5, 114) <= input(11);
output(5, 115) <= input(12);
output(5, 116) <= input(13);
output(5, 117) <= input(14);
output(5, 118) <= input(15);
output(5, 119) <= input(32);
output(5, 120) <= input(34);
output(5, 121) <= input(36);
output(5, 122) <= input(38);
output(5, 123) <= input(40);
output(5, 124) <= input(42);
output(5, 125) <= input(44);
output(5, 126) <= input(46);
output(5, 127) <= input(48);
output(5, 128) <= input(25);
output(5, 129) <= input(26);
output(5, 130) <= input(27);
output(5, 131) <= input(28);
output(5, 132) <= input(29);
output(5, 133) <= input(30);
output(5, 134) <= input(31);
output(5, 135) <= input(33);
output(5, 136) <= input(35);
output(5, 137) <= input(37);
output(5, 138) <= input(39);
output(5, 139) <= input(41);
output(5, 140) <= input(43);
output(5, 141) <= input(45);
output(5, 142) <= input(47);
output(5, 143) <= input(49);
output(5, 144) <= input(10);
output(5, 145) <= input(11);
output(5, 146) <= input(12);
output(5, 147) <= input(13);
output(5, 148) <= input(14);
output(5, 149) <= input(15);
output(5, 150) <= input(32);
output(5, 151) <= input(34);
output(5, 152) <= input(36);
output(5, 153) <= input(38);
output(5, 154) <= input(40);
output(5, 155) <= input(42);
output(5, 156) <= input(44);
output(5, 157) <= input(46);
output(5, 158) <= input(48);
output(5, 159) <= input(50);
output(5, 160) <= input(26);
output(5, 161) <= input(27);
output(5, 162) <= input(28);
output(5, 163) <= input(29);
output(5, 164) <= input(30);
output(5, 165) <= input(31);
output(5, 166) <= input(33);
output(5, 167) <= input(35);
output(5, 168) <= input(37);
output(5, 169) <= input(39);
output(5, 170) <= input(41);
output(5, 171) <= input(43);
output(5, 172) <= input(45);
output(5, 173) <= input(47);
output(5, 174) <= input(49);
output(5, 175) <= input(51);
output(5, 176) <= input(11);
output(5, 177) <= input(12);
output(5, 178) <= input(13);
output(5, 179) <= input(14);
output(5, 180) <= input(15);
output(5, 181) <= input(32);
output(5, 182) <= input(34);
output(5, 183) <= input(36);
output(5, 184) <= input(38);
output(5, 185) <= input(40);
output(5, 186) <= input(42);
output(5, 187) <= input(44);
output(5, 188) <= input(46);
output(5, 189) <= input(48);
output(5, 190) <= input(50);
output(5, 191) <= input(52);
output(5, 192) <= input(27);
output(5, 193) <= input(28);
output(5, 194) <= input(29);
output(5, 195) <= input(30);
output(5, 196) <= input(31);
output(5, 197) <= input(33);
output(5, 198) <= input(35);
output(5, 199) <= input(37);
output(5, 200) <= input(39);
output(5, 201) <= input(41);
output(5, 202) <= input(43);
output(5, 203) <= input(45);
output(5, 204) <= input(47);
output(5, 205) <= input(49);
output(5, 206) <= input(51);
output(5, 207) <= input(53);
output(5, 208) <= input(12);
output(5, 209) <= input(13);
output(5, 210) <= input(14);
output(5, 211) <= input(15);
output(5, 212) <= input(32);
output(5, 213) <= input(34);
output(5, 214) <= input(36);
output(5, 215) <= input(38);
output(5, 216) <= input(40);
output(5, 217) <= input(42);
output(5, 218) <= input(44);
output(5, 219) <= input(46);
output(5, 220) <= input(48);
output(5, 221) <= input(50);
output(5, 222) <= input(52);
output(5, 223) <= input(54);
output(5, 224) <= input(28);
output(5, 225) <= input(29);
output(5, 226) <= input(30);
output(5, 227) <= input(31);
output(5, 228) <= input(33);
output(5, 229) <= input(35);
output(5, 230) <= input(37);
output(5, 231) <= input(39);
output(5, 232) <= input(41);
output(5, 233) <= input(43);
output(5, 234) <= input(45);
output(5, 235) <= input(47);
output(5, 236) <= input(49);
output(5, 237) <= input(51);
output(5, 238) <= input(53);
output(5, 239) <= input(55);
output(5, 240) <= input(13);
output(5, 241) <= input(14);
output(5, 242) <= input(15);
output(5, 243) <= input(32);
output(5, 244) <= input(34);
output(5, 245) <= input(36);
output(5, 246) <= input(38);
output(5, 247) <= input(40);
output(5, 248) <= input(42);
output(5, 249) <= input(44);
output(5, 250) <= input(46);
output(5, 251) <= input(48);
output(5, 252) <= input(50);
output(5, 253) <= input(52);
output(5, 254) <= input(54);
output(5, 255) <= input(56);
when "1111" =>
output(0, 0) <= input(0);
output(0, 1) <= input(1);
output(0, 2) <= input(2);
output(0, 3) <= input(3);
output(0, 4) <= input(4);
output(0, 5) <= input(5);
output(0, 6) <= input(6);
output(0, 7) <= input(7);
output(0, 8) <= input(8);
output(0, 9) <= input(9);
output(0, 10) <= input(10);
output(0, 11) <= input(11);
output(0, 12) <= input(12);
output(0, 13) <= input(13);
output(0, 14) <= input(14);
output(0, 15) <= input(15);
output(0, 16) <= input(16);
output(0, 17) <= input(17);
output(0, 18) <= input(18);
output(0, 19) <= input(19);
output(0, 20) <= input(20);
output(0, 21) <= input(21);
output(0, 22) <= input(22);
output(0, 23) <= input(23);
output(0, 24) <= input(24);
output(0, 25) <= input(25);
output(0, 26) <= input(26);
output(0, 27) <= input(27);
output(0, 28) <= input(28);
output(0, 29) <= input(29);
output(0, 30) <= input(30);
output(0, 31) <= input(31);
output(0, 32) <= input(1);
output(0, 33) <= input(2);
output(0, 34) <= input(3);
output(0, 35) <= input(4);
output(0, 36) <= input(5);
output(0, 37) <= input(6);
output(0, 38) <= input(7);
output(0, 39) <= input(8);
output(0, 40) <= input(9);
output(0, 41) <= input(10);
output(0, 42) <= input(11);
output(0, 43) <= input(12);
output(0, 44) <= input(13);
output(0, 45) <= input(14);
output(0, 46) <= input(15);
output(0, 47) <= input(32);
output(0, 48) <= input(17);
output(0, 49) <= input(18);
output(0, 50) <= input(19);
output(0, 51) <= input(20);
output(0, 52) <= input(21);
output(0, 53) <= input(22);
output(0, 54) <= input(23);
output(0, 55) <= input(24);
output(0, 56) <= input(25);
output(0, 57) <= input(26);
output(0, 58) <= input(27);
output(0, 59) <= input(28);
output(0, 60) <= input(29);
output(0, 61) <= input(30);
output(0, 62) <= input(31);
output(0, 63) <= input(33);
output(0, 64) <= input(2);
output(0, 65) <= input(3);
output(0, 66) <= input(4);
output(0, 67) <= input(5);
output(0, 68) <= input(6);
output(0, 69) <= input(7);
output(0, 70) <= input(8);
output(0, 71) <= input(9);
output(0, 72) <= input(10);
output(0, 73) <= input(11);
output(0, 74) <= input(12);
output(0, 75) <= input(13);
output(0, 76) <= input(14);
output(0, 77) <= input(15);
output(0, 78) <= input(32);
output(0, 79) <= input(34);
output(0, 80) <= input(18);
output(0, 81) <= input(19);
output(0, 82) <= input(20);
output(0, 83) <= input(21);
output(0, 84) <= input(22);
output(0, 85) <= input(23);
output(0, 86) <= input(24);
output(0, 87) <= input(25);
output(0, 88) <= input(26);
output(0, 89) <= input(27);
output(0, 90) <= input(28);
output(0, 91) <= input(29);
output(0, 92) <= input(30);
output(0, 93) <= input(31);
output(0, 94) <= input(33);
output(0, 95) <= input(35);
output(0, 96) <= input(3);
output(0, 97) <= input(4);
output(0, 98) <= input(5);
output(0, 99) <= input(6);
output(0, 100) <= input(7);
output(0, 101) <= input(8);
output(0, 102) <= input(9);
output(0, 103) <= input(10);
output(0, 104) <= input(11);
output(0, 105) <= input(12);
output(0, 106) <= input(13);
output(0, 107) <= input(14);
output(0, 108) <= input(15);
output(0, 109) <= input(32);
output(0, 110) <= input(34);
output(0, 111) <= input(36);
output(0, 112) <= input(4);
output(0, 113) <= input(5);
output(0, 114) <= input(6);
output(0, 115) <= input(7);
output(0, 116) <= input(8);
output(0, 117) <= input(9);
output(0, 118) <= input(10);
output(0, 119) <= input(11);
output(0, 120) <= input(12);
output(0, 121) <= input(13);
output(0, 122) <= input(14);
output(0, 123) <= input(15);
output(0, 124) <= input(32);
output(0, 125) <= input(34);
output(0, 126) <= input(36);
output(0, 127) <= input(37);
output(0, 128) <= input(20);
output(0, 129) <= input(21);
output(0, 130) <= input(22);
output(0, 131) <= input(23);
output(0, 132) <= input(24);
output(0, 133) <= input(25);
output(0, 134) <= input(26);
output(0, 135) <= input(27);
output(0, 136) <= input(28);
output(0, 137) <= input(29);
output(0, 138) <= input(30);
output(0, 139) <= input(31);
output(0, 140) <= input(33);
output(0, 141) <= input(35);
output(0, 142) <= input(38);
output(0, 143) <= input(39);
output(0, 144) <= input(5);
output(0, 145) <= input(6);
output(0, 146) <= input(7);
output(0, 147) <= input(8);
output(0, 148) <= input(9);
output(0, 149) <= input(10);
output(0, 150) <= input(11);
output(0, 151) <= input(12);
output(0, 152) <= input(13);
output(0, 153) <= input(14);
output(0, 154) <= input(15);
output(0, 155) <= input(32);
output(0, 156) <= input(34);
output(0, 157) <= input(36);
output(0, 158) <= input(37);
output(0, 159) <= input(40);
output(0, 160) <= input(21);
output(0, 161) <= input(22);
output(0, 162) <= input(23);
output(0, 163) <= input(24);
output(0, 164) <= input(25);
output(0, 165) <= input(26);
output(0, 166) <= input(27);
output(0, 167) <= input(28);
output(0, 168) <= input(29);
output(0, 169) <= input(30);
output(0, 170) <= input(31);
output(0, 171) <= input(33);
output(0, 172) <= input(35);
output(0, 173) <= input(38);
output(0, 174) <= input(39);
output(0, 175) <= input(41);
output(0, 176) <= input(6);
output(0, 177) <= input(7);
output(0, 178) <= input(8);
output(0, 179) <= input(9);
output(0, 180) <= input(10);
output(0, 181) <= input(11);
output(0, 182) <= input(12);
output(0, 183) <= input(13);
output(0, 184) <= input(14);
output(0, 185) <= input(15);
output(0, 186) <= input(32);
output(0, 187) <= input(34);
output(0, 188) <= input(36);
output(0, 189) <= input(37);
output(0, 190) <= input(40);
output(0, 191) <= input(42);
output(0, 192) <= input(22);
output(0, 193) <= input(23);
output(0, 194) <= input(24);
output(0, 195) <= input(25);
output(0, 196) <= input(26);
output(0, 197) <= input(27);
output(0, 198) <= input(28);
output(0, 199) <= input(29);
output(0, 200) <= input(30);
output(0, 201) <= input(31);
output(0, 202) <= input(33);
output(0, 203) <= input(35);
output(0, 204) <= input(38);
output(0, 205) <= input(39);
output(0, 206) <= input(41);
output(0, 207) <= input(43);
output(0, 208) <= input(7);
output(0, 209) <= input(8);
output(0, 210) <= input(9);
output(0, 211) <= input(10);
output(0, 212) <= input(11);
output(0, 213) <= input(12);
output(0, 214) <= input(13);
output(0, 215) <= input(14);
output(0, 216) <= input(15);
output(0, 217) <= input(32);
output(0, 218) <= input(34);
output(0, 219) <= input(36);
output(0, 220) <= input(37);
output(0, 221) <= input(40);
output(0, 222) <= input(42);
output(0, 223) <= input(44);
output(0, 224) <= input(23);
output(0, 225) <= input(24);
output(0, 226) <= input(25);
output(0, 227) <= input(26);
output(0, 228) <= input(27);
output(0, 229) <= input(28);
output(0, 230) <= input(29);
output(0, 231) <= input(30);
output(0, 232) <= input(31);
output(0, 233) <= input(33);
output(0, 234) <= input(35);
output(0, 235) <= input(38);
output(0, 236) <= input(39);
output(0, 237) <= input(41);
output(0, 238) <= input(43);
output(0, 239) <= input(45);
output(0, 240) <= input(24);
output(0, 241) <= input(25);
output(0, 242) <= input(26);
output(0, 243) <= input(27);
output(0, 244) <= input(28);
output(0, 245) <= input(29);
output(0, 246) <= input(30);
output(0, 247) <= input(31);
output(0, 248) <= input(33);
output(0, 249) <= input(35);
output(0, 250) <= input(38);
output(0, 251) <= input(39);
output(0, 252) <= input(41);
output(0, 253) <= input(43);
output(0, 254) <= input(45);
output(0, 255) <= input(46);
output(1, 0) <= input(1);
output(1, 1) <= input(2);
output(1, 2) <= input(3);
output(1, 3) <= input(4);
output(1, 4) <= input(5);
output(1, 5) <= input(6);
output(1, 6) <= input(7);
output(1, 7) <= input(8);
output(1, 8) <= input(9);
output(1, 9) <= input(10);
output(1, 10) <= input(11);
output(1, 11) <= input(12);
output(1, 12) <= input(13);
output(1, 13) <= input(14);
output(1, 14) <= input(15);
output(1, 15) <= input(32);
output(1, 16) <= input(17);
output(1, 17) <= input(18);
output(1, 18) <= input(19);
output(1, 19) <= input(20);
output(1, 20) <= input(21);
output(1, 21) <= input(22);
output(1, 22) <= input(23);
output(1, 23) <= input(24);
output(1, 24) <= input(25);
output(1, 25) <= input(26);
output(1, 26) <= input(27);
output(1, 27) <= input(28);
output(1, 28) <= input(29);
output(1, 29) <= input(30);
output(1, 30) <= input(31);
output(1, 31) <= input(33);
output(1, 32) <= input(2);
output(1, 33) <= input(3);
output(1, 34) <= input(4);
output(1, 35) <= input(5);
output(1, 36) <= input(6);
output(1, 37) <= input(7);
output(1, 38) <= input(8);
output(1, 39) <= input(9);
output(1, 40) <= input(10);
output(1, 41) <= input(11);
output(1, 42) <= input(12);
output(1, 43) <= input(13);
output(1, 44) <= input(14);
output(1, 45) <= input(15);
output(1, 46) <= input(32);
output(1, 47) <= input(34);
output(1, 48) <= input(3);
output(1, 49) <= input(4);
output(1, 50) <= input(5);
output(1, 51) <= input(6);
output(1, 52) <= input(7);
output(1, 53) <= input(8);
output(1, 54) <= input(9);
output(1, 55) <= input(10);
output(1, 56) <= input(11);
output(1, 57) <= input(12);
output(1, 58) <= input(13);
output(1, 59) <= input(14);
output(1, 60) <= input(15);
output(1, 61) <= input(32);
output(1, 62) <= input(34);
output(1, 63) <= input(36);
output(1, 64) <= input(19);
output(1, 65) <= input(20);
output(1, 66) <= input(21);
output(1, 67) <= input(22);
output(1, 68) <= input(23);
output(1, 69) <= input(24);
output(1, 70) <= input(25);
output(1, 71) <= input(26);
output(1, 72) <= input(27);
output(1, 73) <= input(28);
output(1, 74) <= input(29);
output(1, 75) <= input(30);
output(1, 76) <= input(31);
output(1, 77) <= input(33);
output(1, 78) <= input(35);
output(1, 79) <= input(38);
output(1, 80) <= input(4);
output(1, 81) <= input(5);
output(1, 82) <= input(6);
output(1, 83) <= input(7);
output(1, 84) <= input(8);
output(1, 85) <= input(9);
output(1, 86) <= input(10);
output(1, 87) <= input(11);
output(1, 88) <= input(12);
output(1, 89) <= input(13);
output(1, 90) <= input(14);
output(1, 91) <= input(15);
output(1, 92) <= input(32);
output(1, 93) <= input(34);
output(1, 94) <= input(36);
output(1, 95) <= input(37);
output(1, 96) <= input(20);
output(1, 97) <= input(21);
output(1, 98) <= input(22);
output(1, 99) <= input(23);
output(1, 100) <= input(24);
output(1, 101) <= input(25);
output(1, 102) <= input(26);
output(1, 103) <= input(27);
output(1, 104) <= input(28);
output(1, 105) <= input(29);
output(1, 106) <= input(30);
output(1, 107) <= input(31);
output(1, 108) <= input(33);
output(1, 109) <= input(35);
output(1, 110) <= input(38);
output(1, 111) <= input(39);
output(1, 112) <= input(21);
output(1, 113) <= input(22);
output(1, 114) <= input(23);
output(1, 115) <= input(24);
output(1, 116) <= input(25);
output(1, 117) <= input(26);
output(1, 118) <= input(27);
output(1, 119) <= input(28);
output(1, 120) <= input(29);
output(1, 121) <= input(30);
output(1, 122) <= input(31);
output(1, 123) <= input(33);
output(1, 124) <= input(35);
output(1, 125) <= input(38);
output(1, 126) <= input(39);
output(1, 127) <= input(41);
output(1, 128) <= input(6);
output(1, 129) <= input(7);
output(1, 130) <= input(8);
output(1, 131) <= input(9);
output(1, 132) <= input(10);
output(1, 133) <= input(11);
output(1, 134) <= input(12);
output(1, 135) <= input(13);
output(1, 136) <= input(14);
output(1, 137) <= input(15);
output(1, 138) <= input(32);
output(1, 139) <= input(34);
output(1, 140) <= input(36);
output(1, 141) <= input(37);
output(1, 142) <= input(40);
output(1, 143) <= input(42);
output(1, 144) <= input(22);
output(1, 145) <= input(23);
output(1, 146) <= input(24);
output(1, 147) <= input(25);
output(1, 148) <= input(26);
output(1, 149) <= input(27);
output(1, 150) <= input(28);
output(1, 151) <= input(29);
output(1, 152) <= input(30);
output(1, 153) <= input(31);
output(1, 154) <= input(33);
output(1, 155) <= input(35);
output(1, 156) <= input(38);
output(1, 157) <= input(39);
output(1, 158) <= input(41);
output(1, 159) <= input(43);
output(1, 160) <= input(7);
output(1, 161) <= input(8);
output(1, 162) <= input(9);
output(1, 163) <= input(10);
output(1, 164) <= input(11);
output(1, 165) <= input(12);
output(1, 166) <= input(13);
output(1, 167) <= input(14);
output(1, 168) <= input(15);
output(1, 169) <= input(32);
output(1, 170) <= input(34);
output(1, 171) <= input(36);
output(1, 172) <= input(37);
output(1, 173) <= input(40);
output(1, 174) <= input(42);
output(1, 175) <= input(44);
output(1, 176) <= input(8);
output(1, 177) <= input(9);
output(1, 178) <= input(10);
output(1, 179) <= input(11);
output(1, 180) <= input(12);
output(1, 181) <= input(13);
output(1, 182) <= input(14);
output(1, 183) <= input(15);
output(1, 184) <= input(32);
output(1, 185) <= input(34);
output(1, 186) <= input(36);
output(1, 187) <= input(37);
output(1, 188) <= input(40);
output(1, 189) <= input(42);
output(1, 190) <= input(44);
output(1, 191) <= input(47);
output(1, 192) <= input(24);
output(1, 193) <= input(25);
output(1, 194) <= input(26);
output(1, 195) <= input(27);
output(1, 196) <= input(28);
output(1, 197) <= input(29);
output(1, 198) <= input(30);
output(1, 199) <= input(31);
output(1, 200) <= input(33);
output(1, 201) <= input(35);
output(1, 202) <= input(38);
output(1, 203) <= input(39);
output(1, 204) <= input(41);
output(1, 205) <= input(43);
output(1, 206) <= input(45);
output(1, 207) <= input(46);
output(1, 208) <= input(9);
output(1, 209) <= input(10);
output(1, 210) <= input(11);
output(1, 211) <= input(12);
output(1, 212) <= input(13);
output(1, 213) <= input(14);
output(1, 214) <= input(15);
output(1, 215) <= input(32);
output(1, 216) <= input(34);
output(1, 217) <= input(36);
output(1, 218) <= input(37);
output(1, 219) <= input(40);
output(1, 220) <= input(42);
output(1, 221) <= input(44);
output(1, 222) <= input(47);
output(1, 223) <= input(48);
output(1, 224) <= input(25);
output(1, 225) <= input(26);
output(1, 226) <= input(27);
output(1, 227) <= input(28);
output(1, 228) <= input(29);
output(1, 229) <= input(30);
output(1, 230) <= input(31);
output(1, 231) <= input(33);
output(1, 232) <= input(35);
output(1, 233) <= input(38);
output(1, 234) <= input(39);
output(1, 235) <= input(41);
output(1, 236) <= input(43);
output(1, 237) <= input(45);
output(1, 238) <= input(46);
output(1, 239) <= input(49);
output(1, 240) <= input(26);
output(1, 241) <= input(27);
output(1, 242) <= input(28);
output(1, 243) <= input(29);
output(1, 244) <= input(30);
output(1, 245) <= input(31);
output(1, 246) <= input(33);
output(1, 247) <= input(35);
output(1, 248) <= input(38);
output(1, 249) <= input(39);
output(1, 250) <= input(41);
output(1, 251) <= input(43);
output(1, 252) <= input(45);
output(1, 253) <= input(46);
output(1, 254) <= input(49);
output(1, 255) <= input(50);
output(2, 0) <= input(18);
output(2, 1) <= input(19);
output(2, 2) <= input(20);
output(2, 3) <= input(21);
output(2, 4) <= input(22);
output(2, 5) <= input(23);
output(2, 6) <= input(24);
output(2, 7) <= input(25);
output(2, 8) <= input(26);
output(2, 9) <= input(27);
output(2, 10) <= input(28);
output(2, 11) <= input(29);
output(2, 12) <= input(30);
output(2, 13) <= input(31);
output(2, 14) <= input(33);
output(2, 15) <= input(35);
output(2, 16) <= input(3);
output(2, 17) <= input(4);
output(2, 18) <= input(5);
output(2, 19) <= input(6);
output(2, 20) <= input(7);
output(2, 21) <= input(8);
output(2, 22) <= input(9);
output(2, 23) <= input(10);
output(2, 24) <= input(11);
output(2, 25) <= input(12);
output(2, 26) <= input(13);
output(2, 27) <= input(14);
output(2, 28) <= input(15);
output(2, 29) <= input(32);
output(2, 30) <= input(34);
output(2, 31) <= input(36);
output(2, 32) <= input(4);
output(2, 33) <= input(5);
output(2, 34) <= input(6);
output(2, 35) <= input(7);
output(2, 36) <= input(8);
output(2, 37) <= input(9);
output(2, 38) <= input(10);
output(2, 39) <= input(11);
output(2, 40) <= input(12);
output(2, 41) <= input(13);
output(2, 42) <= input(14);
output(2, 43) <= input(15);
output(2, 44) <= input(32);
output(2, 45) <= input(34);
output(2, 46) <= input(36);
output(2, 47) <= input(37);
output(2, 48) <= input(20);
output(2, 49) <= input(21);
output(2, 50) <= input(22);
output(2, 51) <= input(23);
output(2, 52) <= input(24);
output(2, 53) <= input(25);
output(2, 54) <= input(26);
output(2, 55) <= input(27);
output(2, 56) <= input(28);
output(2, 57) <= input(29);
output(2, 58) <= input(30);
output(2, 59) <= input(31);
output(2, 60) <= input(33);
output(2, 61) <= input(35);
output(2, 62) <= input(38);
output(2, 63) <= input(39);
output(2, 64) <= input(21);
output(2, 65) <= input(22);
output(2, 66) <= input(23);
output(2, 67) <= input(24);
output(2, 68) <= input(25);
output(2, 69) <= input(26);
output(2, 70) <= input(27);
output(2, 71) <= input(28);
output(2, 72) <= input(29);
output(2, 73) <= input(30);
output(2, 74) <= input(31);
output(2, 75) <= input(33);
output(2, 76) <= input(35);
output(2, 77) <= input(38);
output(2, 78) <= input(39);
output(2, 79) <= input(41);
output(2, 80) <= input(6);
output(2, 81) <= input(7);
output(2, 82) <= input(8);
output(2, 83) <= input(9);
output(2, 84) <= input(10);
output(2, 85) <= input(11);
output(2, 86) <= input(12);
output(2, 87) <= input(13);
output(2, 88) <= input(14);
output(2, 89) <= input(15);
output(2, 90) <= input(32);
output(2, 91) <= input(34);
output(2, 92) <= input(36);
output(2, 93) <= input(37);
output(2, 94) <= input(40);
output(2, 95) <= input(42);
output(2, 96) <= input(7);
output(2, 97) <= input(8);
output(2, 98) <= input(9);
output(2, 99) <= input(10);
output(2, 100) <= input(11);
output(2, 101) <= input(12);
output(2, 102) <= input(13);
output(2, 103) <= input(14);
output(2, 104) <= input(15);
output(2, 105) <= input(32);
output(2, 106) <= input(34);
output(2, 107) <= input(36);
output(2, 108) <= input(37);
output(2, 109) <= input(40);
output(2, 110) <= input(42);
output(2, 111) <= input(44);
output(2, 112) <= input(23);
output(2, 113) <= input(24);
output(2, 114) <= input(25);
output(2, 115) <= input(26);
output(2, 116) <= input(27);
output(2, 117) <= input(28);
output(2, 118) <= input(29);
output(2, 119) <= input(30);
output(2, 120) <= input(31);
output(2, 121) <= input(33);
output(2, 122) <= input(35);
output(2, 123) <= input(38);
output(2, 124) <= input(39);
output(2, 125) <= input(41);
output(2, 126) <= input(43);
output(2, 127) <= input(45);
output(2, 128) <= input(8);
output(2, 129) <= input(9);
output(2, 130) <= input(10);
output(2, 131) <= input(11);
output(2, 132) <= input(12);
output(2, 133) <= input(13);
output(2, 134) <= input(14);
output(2, 135) <= input(15);
output(2, 136) <= input(32);
output(2, 137) <= input(34);
output(2, 138) <= input(36);
output(2, 139) <= input(37);
output(2, 140) <= input(40);
output(2, 141) <= input(42);
output(2, 142) <= input(44);
output(2, 143) <= input(47);
output(2, 144) <= input(9);
output(2, 145) <= input(10);
output(2, 146) <= input(11);
output(2, 147) <= input(12);
output(2, 148) <= input(13);
output(2, 149) <= input(14);
output(2, 150) <= input(15);
output(2, 151) <= input(32);
output(2, 152) <= input(34);
output(2, 153) <= input(36);
output(2, 154) <= input(37);
output(2, 155) <= input(40);
output(2, 156) <= input(42);
output(2, 157) <= input(44);
output(2, 158) <= input(47);
output(2, 159) <= input(48);
output(2, 160) <= input(25);
output(2, 161) <= input(26);
output(2, 162) <= input(27);
output(2, 163) <= input(28);
output(2, 164) <= input(29);
output(2, 165) <= input(30);
output(2, 166) <= input(31);
output(2, 167) <= input(33);
output(2, 168) <= input(35);
output(2, 169) <= input(38);
output(2, 170) <= input(39);
output(2, 171) <= input(41);
output(2, 172) <= input(43);
output(2, 173) <= input(45);
output(2, 174) <= input(46);
output(2, 175) <= input(49);
output(2, 176) <= input(26);
output(2, 177) <= input(27);
output(2, 178) <= input(28);
output(2, 179) <= input(29);
output(2, 180) <= input(30);
output(2, 181) <= input(31);
output(2, 182) <= input(33);
output(2, 183) <= input(35);
output(2, 184) <= input(38);
output(2, 185) <= input(39);
output(2, 186) <= input(41);
output(2, 187) <= input(43);
output(2, 188) <= input(45);
output(2, 189) <= input(46);
output(2, 190) <= input(49);
output(2, 191) <= input(50);
output(2, 192) <= input(11);
output(2, 193) <= input(12);
output(2, 194) <= input(13);
output(2, 195) <= input(14);
output(2, 196) <= input(15);
output(2, 197) <= input(32);
output(2, 198) <= input(34);
output(2, 199) <= input(36);
output(2, 200) <= input(37);
output(2, 201) <= input(40);
output(2, 202) <= input(42);
output(2, 203) <= input(44);
output(2, 204) <= input(47);
output(2, 205) <= input(48);
output(2, 206) <= input(51);
output(2, 207) <= input(52);
output(2, 208) <= input(12);
output(2, 209) <= input(13);
output(2, 210) <= input(14);
output(2, 211) <= input(15);
output(2, 212) <= input(32);
output(2, 213) <= input(34);
output(2, 214) <= input(36);
output(2, 215) <= input(37);
output(2, 216) <= input(40);
output(2, 217) <= input(42);
output(2, 218) <= input(44);
output(2, 219) <= input(47);
output(2, 220) <= input(48);
output(2, 221) <= input(51);
output(2, 222) <= input(52);
output(2, 223) <= input(53);
output(2, 224) <= input(28);
output(2, 225) <= input(29);
output(2, 226) <= input(30);
output(2, 227) <= input(31);
output(2, 228) <= input(33);
output(2, 229) <= input(35);
output(2, 230) <= input(38);
output(2, 231) <= input(39);
output(2, 232) <= input(41);
output(2, 233) <= input(43);
output(2, 234) <= input(45);
output(2, 235) <= input(46);
output(2, 236) <= input(49);
output(2, 237) <= input(50);
output(2, 238) <= input(54);
output(2, 239) <= input(55);
output(2, 240) <= input(29);
output(2, 241) <= input(30);
output(2, 242) <= input(31);
output(2, 243) <= input(33);
output(2, 244) <= input(35);
output(2, 245) <= input(38);
output(2, 246) <= input(39);
output(2, 247) <= input(41);
output(2, 248) <= input(43);
output(2, 249) <= input(45);
output(2, 250) <= input(46);
output(2, 251) <= input(49);
output(2, 252) <= input(50);
output(2, 253) <= input(54);
output(2, 254) <= input(55);
output(2, 255) <= input(56);
output(3, 0) <= input(4);
output(3, 1) <= input(5);
output(3, 2) <= input(6);
output(3, 3) <= input(7);
output(3, 4) <= input(8);
output(3, 5) <= input(9);
output(3, 6) <= input(10);
output(3, 7) <= input(11);
output(3, 8) <= input(12);
output(3, 9) <= input(13);
output(3, 10) <= input(14);
output(3, 11) <= input(15);
output(3, 12) <= input(32);
output(3, 13) <= input(34);
output(3, 14) <= input(36);
output(3, 15) <= input(37);
output(3, 16) <= input(5);
output(3, 17) <= input(6);
output(3, 18) <= input(7);
output(3, 19) <= input(8);
output(3, 20) <= input(9);
output(3, 21) <= input(10);
output(3, 22) <= input(11);
output(3, 23) <= input(12);
output(3, 24) <= input(13);
output(3, 25) <= input(14);
output(3, 26) <= input(15);
output(3, 27) <= input(32);
output(3, 28) <= input(34);
output(3, 29) <= input(36);
output(3, 30) <= input(37);
output(3, 31) <= input(40);
output(3, 32) <= input(21);
output(3, 33) <= input(22);
output(3, 34) <= input(23);
output(3, 35) <= input(24);
output(3, 36) <= input(25);
output(3, 37) <= input(26);
output(3, 38) <= input(27);
output(3, 39) <= input(28);
output(3, 40) <= input(29);
output(3, 41) <= input(30);
output(3, 42) <= input(31);
output(3, 43) <= input(33);
output(3, 44) <= input(35);
output(3, 45) <= input(38);
output(3, 46) <= input(39);
output(3, 47) <= input(41);
output(3, 48) <= input(22);
output(3, 49) <= input(23);
output(3, 50) <= input(24);
output(3, 51) <= input(25);
output(3, 52) <= input(26);
output(3, 53) <= input(27);
output(3, 54) <= input(28);
output(3, 55) <= input(29);
output(3, 56) <= input(30);
output(3, 57) <= input(31);
output(3, 58) <= input(33);
output(3, 59) <= input(35);
output(3, 60) <= input(38);
output(3, 61) <= input(39);
output(3, 62) <= input(41);
output(3, 63) <= input(43);
output(3, 64) <= input(23);
output(3, 65) <= input(24);
output(3, 66) <= input(25);
output(3, 67) <= input(26);
output(3, 68) <= input(27);
output(3, 69) <= input(28);
output(3, 70) <= input(29);
output(3, 71) <= input(30);
output(3, 72) <= input(31);
output(3, 73) <= input(33);
output(3, 74) <= input(35);
output(3, 75) <= input(38);
output(3, 76) <= input(39);
output(3, 77) <= input(41);
output(3, 78) <= input(43);
output(3, 79) <= input(45);
output(3, 80) <= input(8);
output(3, 81) <= input(9);
output(3, 82) <= input(10);
output(3, 83) <= input(11);
output(3, 84) <= input(12);
output(3, 85) <= input(13);
output(3, 86) <= input(14);
output(3, 87) <= input(15);
output(3, 88) <= input(32);
output(3, 89) <= input(34);
output(3, 90) <= input(36);
output(3, 91) <= input(37);
output(3, 92) <= input(40);
output(3, 93) <= input(42);
output(3, 94) <= input(44);
output(3, 95) <= input(47);
output(3, 96) <= input(9);
output(3, 97) <= input(10);
output(3, 98) <= input(11);
output(3, 99) <= input(12);
output(3, 100) <= input(13);
output(3, 101) <= input(14);
output(3, 102) <= input(15);
output(3, 103) <= input(32);
output(3, 104) <= input(34);
output(3, 105) <= input(36);
output(3, 106) <= input(37);
output(3, 107) <= input(40);
output(3, 108) <= input(42);
output(3, 109) <= input(44);
output(3, 110) <= input(47);
output(3, 111) <= input(48);
output(3, 112) <= input(10);
output(3, 113) <= input(11);
output(3, 114) <= input(12);
output(3, 115) <= input(13);
output(3, 116) <= input(14);
output(3, 117) <= input(15);
output(3, 118) <= input(32);
output(3, 119) <= input(34);
output(3, 120) <= input(36);
output(3, 121) <= input(37);
output(3, 122) <= input(40);
output(3, 123) <= input(42);
output(3, 124) <= input(44);
output(3, 125) <= input(47);
output(3, 126) <= input(48);
output(3, 127) <= input(51);
output(3, 128) <= input(26);
output(3, 129) <= input(27);
output(3, 130) <= input(28);
output(3, 131) <= input(29);
output(3, 132) <= input(30);
output(3, 133) <= input(31);
output(3, 134) <= input(33);
output(3, 135) <= input(35);
output(3, 136) <= input(38);
output(3, 137) <= input(39);
output(3, 138) <= input(41);
output(3, 139) <= input(43);
output(3, 140) <= input(45);
output(3, 141) <= input(46);
output(3, 142) <= input(49);
output(3, 143) <= input(50);
output(3, 144) <= input(27);
output(3, 145) <= input(28);
output(3, 146) <= input(29);
output(3, 147) <= input(30);
output(3, 148) <= input(31);
output(3, 149) <= input(33);
output(3, 150) <= input(35);
output(3, 151) <= input(38);
output(3, 152) <= input(39);
output(3, 153) <= input(41);
output(3, 154) <= input(43);
output(3, 155) <= input(45);
output(3, 156) <= input(46);
output(3, 157) <= input(49);
output(3, 158) <= input(50);
output(3, 159) <= input(54);
output(3, 160) <= input(12);
output(3, 161) <= input(13);
output(3, 162) <= input(14);
output(3, 163) <= input(15);
output(3, 164) <= input(32);
output(3, 165) <= input(34);
output(3, 166) <= input(36);
output(3, 167) <= input(37);
output(3, 168) <= input(40);
output(3, 169) <= input(42);
output(3, 170) <= input(44);
output(3, 171) <= input(47);
output(3, 172) <= input(48);
output(3, 173) <= input(51);
output(3, 174) <= input(52);
output(3, 175) <= input(53);
output(3, 176) <= input(13);
output(3, 177) <= input(14);
output(3, 178) <= input(15);
output(3, 179) <= input(32);
output(3, 180) <= input(34);
output(3, 181) <= input(36);
output(3, 182) <= input(37);
output(3, 183) <= input(40);
output(3, 184) <= input(42);
output(3, 185) <= input(44);
output(3, 186) <= input(47);
output(3, 187) <= input(48);
output(3, 188) <= input(51);
output(3, 189) <= input(52);
output(3, 190) <= input(53);
output(3, 191) <= input(57);
output(3, 192) <= input(14);
output(3, 193) <= input(15);
output(3, 194) <= input(32);
output(3, 195) <= input(34);
output(3, 196) <= input(36);
output(3, 197) <= input(37);
output(3, 198) <= input(40);
output(3, 199) <= input(42);
output(3, 200) <= input(44);
output(3, 201) <= input(47);
output(3, 202) <= input(48);
output(3, 203) <= input(51);
output(3, 204) <= input(52);
output(3, 205) <= input(53);
output(3, 206) <= input(57);
output(3, 207) <= input(58);
output(3, 208) <= input(30);
output(3, 209) <= input(31);
output(3, 210) <= input(33);
output(3, 211) <= input(35);
output(3, 212) <= input(38);
output(3, 213) <= input(39);
output(3, 214) <= input(41);
output(3, 215) <= input(43);
output(3, 216) <= input(45);
output(3, 217) <= input(46);
output(3, 218) <= input(49);
output(3, 219) <= input(50);
output(3, 220) <= input(54);
output(3, 221) <= input(55);
output(3, 222) <= input(56);
output(3, 223) <= input(59);
output(3, 224) <= input(31);
output(3, 225) <= input(33);
output(3, 226) <= input(35);
output(3, 227) <= input(38);
output(3, 228) <= input(39);
output(3, 229) <= input(41);
output(3, 230) <= input(43);
output(3, 231) <= input(45);
output(3, 232) <= input(46);
output(3, 233) <= input(49);
output(3, 234) <= input(50);
output(3, 235) <= input(54);
output(3, 236) <= input(55);
output(3, 237) <= input(56);
output(3, 238) <= input(59);
output(3, 239) <= input(60);
output(3, 240) <= input(33);
output(3, 241) <= input(35);
output(3, 242) <= input(38);
output(3, 243) <= input(39);
output(3, 244) <= input(41);
output(3, 245) <= input(43);
output(3, 246) <= input(45);
output(3, 247) <= input(46);
output(3, 248) <= input(49);
output(3, 249) <= input(50);
output(3, 250) <= input(54);
output(3, 251) <= input(55);
output(3, 252) <= input(56);
output(3, 253) <= input(59);
output(3, 254) <= input(60);
output(3, 255) <= input(61);
output(4, 0) <= input(21);
output(4, 1) <= input(22);
output(4, 2) <= input(23);
output(4, 3) <= input(24);
output(4, 4) <= input(25);
output(4, 5) <= input(26);
output(4, 6) <= input(27);
output(4, 7) <= input(28);
output(4, 8) <= input(29);
output(4, 9) <= input(30);
output(4, 10) <= input(31);
output(4, 11) <= input(33);
output(4, 12) <= input(35);
output(4, 13) <= input(38);
output(4, 14) <= input(39);
output(4, 15) <= input(41);
output(4, 16) <= input(22);
output(4, 17) <= input(23);
output(4, 18) <= input(24);
output(4, 19) <= input(25);
output(4, 20) <= input(26);
output(4, 21) <= input(27);
output(4, 22) <= input(28);
output(4, 23) <= input(29);
output(4, 24) <= input(30);
output(4, 25) <= input(31);
output(4, 26) <= input(33);
output(4, 27) <= input(35);
output(4, 28) <= input(38);
output(4, 29) <= input(39);
output(4, 30) <= input(41);
output(4, 31) <= input(43);
output(4, 32) <= input(23);
output(4, 33) <= input(24);
output(4, 34) <= input(25);
output(4, 35) <= input(26);
output(4, 36) <= input(27);
output(4, 37) <= input(28);
output(4, 38) <= input(29);
output(4, 39) <= input(30);
output(4, 40) <= input(31);
output(4, 41) <= input(33);
output(4, 42) <= input(35);
output(4, 43) <= input(38);
output(4, 44) <= input(39);
output(4, 45) <= input(41);
output(4, 46) <= input(43);
output(4, 47) <= input(45);
output(4, 48) <= input(24);
output(4, 49) <= input(25);
output(4, 50) <= input(26);
output(4, 51) <= input(27);
output(4, 52) <= input(28);
output(4, 53) <= input(29);
output(4, 54) <= input(30);
output(4, 55) <= input(31);
output(4, 56) <= input(33);
output(4, 57) <= input(35);
output(4, 58) <= input(38);
output(4, 59) <= input(39);
output(4, 60) <= input(41);
output(4, 61) <= input(43);
output(4, 62) <= input(45);
output(4, 63) <= input(46);
output(4, 64) <= input(25);
output(4, 65) <= input(26);
output(4, 66) <= input(27);
output(4, 67) <= input(28);
output(4, 68) <= input(29);
output(4, 69) <= input(30);
output(4, 70) <= input(31);
output(4, 71) <= input(33);
output(4, 72) <= input(35);
output(4, 73) <= input(38);
output(4, 74) <= input(39);
output(4, 75) <= input(41);
output(4, 76) <= input(43);
output(4, 77) <= input(45);
output(4, 78) <= input(46);
output(4, 79) <= input(49);
output(4, 80) <= input(10);
output(4, 81) <= input(11);
output(4, 82) <= input(12);
output(4, 83) <= input(13);
output(4, 84) <= input(14);
output(4, 85) <= input(15);
output(4, 86) <= input(32);
output(4, 87) <= input(34);
output(4, 88) <= input(36);
output(4, 89) <= input(37);
output(4, 90) <= input(40);
output(4, 91) <= input(42);
output(4, 92) <= input(44);
output(4, 93) <= input(47);
output(4, 94) <= input(48);
output(4, 95) <= input(51);
output(4, 96) <= input(11);
output(4, 97) <= input(12);
output(4, 98) <= input(13);
output(4, 99) <= input(14);
output(4, 100) <= input(15);
output(4, 101) <= input(32);
output(4, 102) <= input(34);
output(4, 103) <= input(36);
output(4, 104) <= input(37);
output(4, 105) <= input(40);
output(4, 106) <= input(42);
output(4, 107) <= input(44);
output(4, 108) <= input(47);
output(4, 109) <= input(48);
output(4, 110) <= input(51);
output(4, 111) <= input(52);
output(4, 112) <= input(12);
output(4, 113) <= input(13);
output(4, 114) <= input(14);
output(4, 115) <= input(15);
output(4, 116) <= input(32);
output(4, 117) <= input(34);
output(4, 118) <= input(36);
output(4, 119) <= input(37);
output(4, 120) <= input(40);
output(4, 121) <= input(42);
output(4, 122) <= input(44);
output(4, 123) <= input(47);
output(4, 124) <= input(48);
output(4, 125) <= input(51);
output(4, 126) <= input(52);
output(4, 127) <= input(53);
output(4, 128) <= input(13);
output(4, 129) <= input(14);
output(4, 130) <= input(15);
output(4, 131) <= input(32);
output(4, 132) <= input(34);
output(4, 133) <= input(36);
output(4, 134) <= input(37);
output(4, 135) <= input(40);
output(4, 136) <= input(42);
output(4, 137) <= input(44);
output(4, 138) <= input(47);
output(4, 139) <= input(48);
output(4, 140) <= input(51);
output(4, 141) <= input(52);
output(4, 142) <= input(53);
output(4, 143) <= input(57);
output(4, 144) <= input(14);
output(4, 145) <= input(15);
output(4, 146) <= input(32);
output(4, 147) <= input(34);
output(4, 148) <= input(36);
output(4, 149) <= input(37);
output(4, 150) <= input(40);
output(4, 151) <= input(42);
output(4, 152) <= input(44);
output(4, 153) <= input(47);
output(4, 154) <= input(48);
output(4, 155) <= input(51);
output(4, 156) <= input(52);
output(4, 157) <= input(53);
output(4, 158) <= input(57);
output(4, 159) <= input(58);
output(4, 160) <= input(30);
output(4, 161) <= input(31);
output(4, 162) <= input(33);
output(4, 163) <= input(35);
output(4, 164) <= input(38);
output(4, 165) <= input(39);
output(4, 166) <= input(41);
output(4, 167) <= input(43);
output(4, 168) <= input(45);
output(4, 169) <= input(46);
output(4, 170) <= input(49);
output(4, 171) <= input(50);
output(4, 172) <= input(54);
output(4, 173) <= input(55);
output(4, 174) <= input(56);
output(4, 175) <= input(59);
output(4, 176) <= input(31);
output(4, 177) <= input(33);
output(4, 178) <= input(35);
output(4, 179) <= input(38);
output(4, 180) <= input(39);
output(4, 181) <= input(41);
output(4, 182) <= input(43);
output(4, 183) <= input(45);
output(4, 184) <= input(46);
output(4, 185) <= input(49);
output(4, 186) <= input(50);
output(4, 187) <= input(54);
output(4, 188) <= input(55);
output(4, 189) <= input(56);
output(4, 190) <= input(59);
output(4, 191) <= input(60);
output(4, 192) <= input(33);
output(4, 193) <= input(35);
output(4, 194) <= input(38);
output(4, 195) <= input(39);
output(4, 196) <= input(41);
output(4, 197) <= input(43);
output(4, 198) <= input(45);
output(4, 199) <= input(46);
output(4, 200) <= input(49);
output(4, 201) <= input(50);
output(4, 202) <= input(54);
output(4, 203) <= input(55);
output(4, 204) <= input(56);
output(4, 205) <= input(59);
output(4, 206) <= input(60);
output(4, 207) <= input(61);
output(4, 208) <= input(35);
output(4, 209) <= input(38);
output(4, 210) <= input(39);
output(4, 211) <= input(41);
output(4, 212) <= input(43);
output(4, 213) <= input(45);
output(4, 214) <= input(46);
output(4, 215) <= input(49);
output(4, 216) <= input(50);
output(4, 217) <= input(54);
output(4, 218) <= input(55);
output(4, 219) <= input(56);
output(4, 220) <= input(59);
output(4, 221) <= input(60);
output(4, 222) <= input(61);
output(4, 223) <= input(62);
output(4, 224) <= input(38);
output(4, 225) <= input(39);
output(4, 226) <= input(41);
output(4, 227) <= input(43);
output(4, 228) <= input(45);
output(4, 229) <= input(46);
output(4, 230) <= input(49);
output(4, 231) <= input(50);
output(4, 232) <= input(54);
output(4, 233) <= input(55);
output(4, 234) <= input(56);
output(4, 235) <= input(59);
output(4, 236) <= input(60);
output(4, 237) <= input(61);
output(4, 238) <= input(62);
output(4, 239) <= input(63);
output(4, 240) <= input(39);
output(4, 241) <= input(41);
output(4, 242) <= input(43);
output(4, 243) <= input(45);
output(4, 244) <= input(46);
output(4, 245) <= input(49);
output(4, 246) <= input(50);
output(4, 247) <= input(54);
output(4, 248) <= input(55);
output(4, 249) <= input(56);
output(4, 250) <= input(59);
output(4, 251) <= input(60);
output(4, 252) <= input(61);
output(4, 253) <= input(62);
output(4, 254) <= input(63);
output(4, 255) <= input(64);
output(5, 0) <= input(23);
output(5, 1) <= input(24);
output(5, 2) <= input(25);
output(5, 3) <= input(26);
output(5, 4) <= input(27);
output(5, 5) <= input(28);
output(5, 6) <= input(29);
output(5, 7) <= input(30);
output(5, 8) <= input(31);
output(5, 9) <= input(33);
output(5, 10) <= input(35);
output(5, 11) <= input(38);
output(5, 12) <= input(39);
output(5, 13) <= input(41);
output(5, 14) <= input(43);
output(5, 15) <= input(45);
output(5, 16) <= input(24);
output(5, 17) <= input(25);
output(5, 18) <= input(26);
output(5, 19) <= input(27);
output(5, 20) <= input(28);
output(5, 21) <= input(29);
output(5, 22) <= input(30);
output(5, 23) <= input(31);
output(5, 24) <= input(33);
output(5, 25) <= input(35);
output(5, 26) <= input(38);
output(5, 27) <= input(39);
output(5, 28) <= input(41);
output(5, 29) <= input(43);
output(5, 30) <= input(45);
output(5, 31) <= input(46);
output(5, 32) <= input(25);
output(5, 33) <= input(26);
output(5, 34) <= input(27);
output(5, 35) <= input(28);
output(5, 36) <= input(29);
output(5, 37) <= input(30);
output(5, 38) <= input(31);
output(5, 39) <= input(33);
output(5, 40) <= input(35);
output(5, 41) <= input(38);
output(5, 42) <= input(39);
output(5, 43) <= input(41);
output(5, 44) <= input(43);
output(5, 45) <= input(45);
output(5, 46) <= input(46);
output(5, 47) <= input(49);
output(5, 48) <= input(26);
output(5, 49) <= input(27);
output(5, 50) <= input(28);
output(5, 51) <= input(29);
output(5, 52) <= input(30);
output(5, 53) <= input(31);
output(5, 54) <= input(33);
output(5, 55) <= input(35);
output(5, 56) <= input(38);
output(5, 57) <= input(39);
output(5, 58) <= input(41);
output(5, 59) <= input(43);
output(5, 60) <= input(45);
output(5, 61) <= input(46);
output(5, 62) <= input(49);
output(5, 63) <= input(50);
output(5, 64) <= input(27);
output(5, 65) <= input(28);
output(5, 66) <= input(29);
output(5, 67) <= input(30);
output(5, 68) <= input(31);
output(5, 69) <= input(33);
output(5, 70) <= input(35);
output(5, 71) <= input(38);
output(5, 72) <= input(39);
output(5, 73) <= input(41);
output(5, 74) <= input(43);
output(5, 75) <= input(45);
output(5, 76) <= input(46);
output(5, 77) <= input(49);
output(5, 78) <= input(50);
output(5, 79) <= input(54);
output(5, 80) <= input(28);
output(5, 81) <= input(29);
output(5, 82) <= input(30);
output(5, 83) <= input(31);
output(5, 84) <= input(33);
output(5, 85) <= input(35);
output(5, 86) <= input(38);
output(5, 87) <= input(39);
output(5, 88) <= input(41);
output(5, 89) <= input(43);
output(5, 90) <= input(45);
output(5, 91) <= input(46);
output(5, 92) <= input(49);
output(5, 93) <= input(50);
output(5, 94) <= input(54);
output(5, 95) <= input(55);
output(5, 96) <= input(29);
output(5, 97) <= input(30);
output(5, 98) <= input(31);
output(5, 99) <= input(33);
output(5, 100) <= input(35);
output(5, 101) <= input(38);
output(5, 102) <= input(39);
output(5, 103) <= input(41);
output(5, 104) <= input(43);
output(5, 105) <= input(45);
output(5, 106) <= input(46);
output(5, 107) <= input(49);
output(5, 108) <= input(50);
output(5, 109) <= input(54);
output(5, 110) <= input(55);
output(5, 111) <= input(56);
output(5, 112) <= input(30);
output(5, 113) <= input(31);
output(5, 114) <= input(33);
output(5, 115) <= input(35);
output(5, 116) <= input(38);
output(5, 117) <= input(39);
output(5, 118) <= input(41);
output(5, 119) <= input(43);
output(5, 120) <= input(45);
output(5, 121) <= input(46);
output(5, 122) <= input(49);
output(5, 123) <= input(50);
output(5, 124) <= input(54);
output(5, 125) <= input(55);
output(5, 126) <= input(56);
output(5, 127) <= input(59);
output(5, 128) <= input(31);
output(5, 129) <= input(33);
output(5, 130) <= input(35);
output(5, 131) <= input(38);
output(5, 132) <= input(39);
output(5, 133) <= input(41);
output(5, 134) <= input(43);
output(5, 135) <= input(45);
output(5, 136) <= input(46);
output(5, 137) <= input(49);
output(5, 138) <= input(50);
output(5, 139) <= input(54);
output(5, 140) <= input(55);
output(5, 141) <= input(56);
output(5, 142) <= input(59);
output(5, 143) <= input(60);
output(5, 144) <= input(33);
output(5, 145) <= input(35);
output(5, 146) <= input(38);
output(5, 147) <= input(39);
output(5, 148) <= input(41);
output(5, 149) <= input(43);
output(5, 150) <= input(45);
output(5, 151) <= input(46);
output(5, 152) <= input(49);
output(5, 153) <= input(50);
output(5, 154) <= input(54);
output(5, 155) <= input(55);
output(5, 156) <= input(56);
output(5, 157) <= input(59);
output(5, 158) <= input(60);
output(5, 159) <= input(61);
output(5, 160) <= input(35);
output(5, 161) <= input(38);
output(5, 162) <= input(39);
output(5, 163) <= input(41);
output(5, 164) <= input(43);
output(5, 165) <= input(45);
output(5, 166) <= input(46);
output(5, 167) <= input(49);
output(5, 168) <= input(50);
output(5, 169) <= input(54);
output(5, 170) <= input(55);
output(5, 171) <= input(56);
output(5, 172) <= input(59);
output(5, 173) <= input(60);
output(5, 174) <= input(61);
output(5, 175) <= input(62);
output(5, 176) <= input(38);
output(5, 177) <= input(39);
output(5, 178) <= input(41);
output(5, 179) <= input(43);
output(5, 180) <= input(45);
output(5, 181) <= input(46);
output(5, 182) <= input(49);
output(5, 183) <= input(50);
output(5, 184) <= input(54);
output(5, 185) <= input(55);
output(5, 186) <= input(56);
output(5, 187) <= input(59);
output(5, 188) <= input(60);
output(5, 189) <= input(61);
output(5, 190) <= input(62);
output(5, 191) <= input(63);
output(5, 192) <= input(39);
output(5, 193) <= input(41);
output(5, 194) <= input(43);
output(5, 195) <= input(45);
output(5, 196) <= input(46);
output(5, 197) <= input(49);
output(5, 198) <= input(50);
output(5, 199) <= input(54);
output(5, 200) <= input(55);
output(5, 201) <= input(56);
output(5, 202) <= input(59);
output(5, 203) <= input(60);
output(5, 204) <= input(61);
output(5, 205) <= input(62);
output(5, 206) <= input(63);
output(5, 207) <= input(64);
output(5, 208) <= input(41);
output(5, 209) <= input(43);
output(5, 210) <= input(45);
output(5, 211) <= input(46);
output(5, 212) <= input(49);
output(5, 213) <= input(50);
output(5, 214) <= input(54);
output(5, 215) <= input(55);
output(5, 216) <= input(56);
output(5, 217) <= input(59);
output(5, 218) <= input(60);
output(5, 219) <= input(61);
output(5, 220) <= input(62);
output(5, 221) <= input(63);
output(5, 222) <= input(64);
output(5, 223) <= input(65);
output(5, 224) <= input(43);
output(5, 225) <= input(45);
output(5, 226) <= input(46);
output(5, 227) <= input(49);
output(5, 228) <= input(50);
output(5, 229) <= input(54);
output(5, 230) <= input(55);
output(5, 231) <= input(56);
output(5, 232) <= input(59);
output(5, 233) <= input(60);
output(5, 234) <= input(61);
output(5, 235) <= input(62);
output(5, 236) <= input(63);
output(5, 237) <= input(64);
output(5, 238) <= input(65);
output(5, 239) <= input(66);
output(5, 240) <= input(45);
output(5, 241) <= input(46);
output(5, 242) <= input(49);
output(5, 243) <= input(50);
output(5, 244) <= input(54);
output(5, 245) <= input(55);
output(5, 246) <= input(56);
output(5, 247) <= input(59);
output(5, 248) <= input(60);
output(5, 249) <= input(61);
output(5, 250) <= input(62);
output(5, 251) <= input(63);
output(5, 252) <= input(64);
output(5, 253) <= input(65);
output(5, 254) <= input(66);
output(5, 255) <= input(67);
when others => for i in 0 to 7 loop for j in 0 to 255 loop output(i,j) <= "00000000"; end loop; end loop;
end case;
		end if;
	end process;
END comportamental;
